//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283, new_n1284, new_n1285;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  INV_X1    g0004(.A(G68), .ZN(new_n205));
  INV_X1    g0005(.A(G238), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  INV_X1    g0007(.A(G264), .ZN(new_n208));
  OAI22_X1  g0008(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g0009(.A(new_n209), .B1(G50), .B2(G226), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G232), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR3_X1   g0021(.A1(new_n215), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G77), .A2(G244), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n204), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT1), .Z(new_n225));
  NOR2_X1   g0025(.A1(G58), .A2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(G13), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n204), .A2(new_n232), .ZN(new_n233));
  AOI211_X1 g0033(.A(new_n220), .B(new_n233), .C1(new_n214), .C2(new_n208), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT0), .ZN(new_n235));
  NOR3_X1   g0035(.A1(new_n225), .A2(new_n231), .A3(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n217), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  OAI21_X1  g0051(.A(G20), .B1(new_n227), .B2(G50), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT65), .B1(G20), .B2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR3_X1   g0058(.A1(KEYINPUT65), .A2(G20), .A3(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G150), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n252), .B1(new_n255), .B2(new_n256), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n230), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n263), .A2(new_n230), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G1), .B2(new_n229), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G50), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT66), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(G50), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n268), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n269), .B1(new_n268), .B2(new_n273), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n265), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  OR2_X1    g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G222), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G223), .A2(G1698), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G1), .A3(G13), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n285), .B(new_n288), .C1(G77), .C2(new_n281), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G226), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n287), .A2(new_n290), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n289), .B(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(KEYINPUT9), .B(new_n265), .C1(new_n274), .C2(new_n275), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n278), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n296), .A2(G200), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT68), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n278), .A2(new_n298), .A3(KEYINPUT68), .A4(new_n299), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(new_n303), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT69), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT10), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n309), .B1(new_n308), .B2(KEYINPUT10), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n304), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n296), .A2(G179), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n313), .A2(KEYINPUT67), .ZN(new_n314));
  INV_X1    g0114(.A(G169), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n296), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n313), .A2(KEYINPUT67), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n314), .A2(new_n316), .A3(new_n276), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G238), .A2(G1698), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n281), .B(new_n319), .C1(new_n212), .C2(G1698), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n320), .B(new_n288), .C1(G107), .C2(new_n281), .ZN(new_n321));
  INV_X1    g0121(.A(G244), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n321), .B(new_n293), .C1(new_n322), .C2(new_n295), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n315), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n260), .A2(new_n256), .ZN(new_n325));
  OR2_X1    g0125(.A1(KEYINPUT15), .A2(G87), .ZN(new_n326));
  NAND2_X1  g0126(.A1(KEYINPUT15), .A2(G87), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G77), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n328), .A2(new_n255), .B1(new_n229), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n264), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n267), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G77), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n331), .B(new_n333), .C1(G77), .C2(new_n271), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n324), .B(new_n334), .C1(G179), .C2(new_n323), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n312), .A2(new_n318), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT71), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT65), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(new_n229), .A3(new_n253), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n257), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n337), .B1(new_n340), .B2(G159), .ZN(new_n341));
  INV_X1    g0141(.A(G159), .ZN(new_n342));
  AOI211_X1 g0142(.A(KEYINPUT71), .B(new_n342), .C1(new_n339), .C2(new_n257), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g0144(.A1(KEYINPUT3), .A2(G33), .ZN(new_n345));
  NOR2_X1   g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT7), .B1(new_n347), .B2(new_n229), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  NOR4_X1   g0149(.A1(new_n345), .A2(new_n346), .A3(new_n349), .A4(G20), .ZN(new_n350));
  OAI21_X1  g0150(.A(G68), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n211), .A2(new_n205), .ZN(new_n352));
  OAI21_X1  g0152(.A(G20), .B1(new_n352), .B2(new_n226), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n344), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT16), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n344), .A2(new_n351), .A3(KEYINPUT16), .A4(new_n353), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n264), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n294), .A2(G1698), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n281), .B(new_n359), .C1(G223), .C2(G1698), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n288), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n295), .A2(new_n212), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n363), .A2(new_n297), .A3(new_n293), .A4(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n287), .B1(new_n360), .B2(new_n361), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n367), .A2(new_n292), .A3(new_n364), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n366), .B1(new_n368), .B2(G200), .ZN(new_n369));
  INV_X1    g0169(.A(new_n271), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n256), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n256), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n332), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n358), .A2(new_n369), .A3(new_n371), .A4(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT17), .ZN(new_n375));
  OR2_X1    g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n375), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n358), .A2(new_n371), .A3(new_n373), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n368), .A2(G169), .ZN(new_n380));
  NOR4_X1   g0180(.A1(new_n367), .A2(G179), .A3(new_n292), .A4(new_n364), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(KEYINPUT18), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT72), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT18), .B1(new_n379), .B2(new_n382), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  AOI211_X1 g0188(.A(KEYINPUT72), .B(KEYINPUT18), .C1(new_n379), .C2(new_n382), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n378), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT13), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n294), .A2(new_n282), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n212), .A2(G1698), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n393), .B(new_n394), .C1(new_n345), .C2(new_n346), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n292), .B1(new_n397), .B2(new_n288), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n287), .A2(G238), .A3(new_n290), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n392), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n287), .B1(new_n395), .B2(new_n396), .ZN(new_n402));
  NOR4_X1   g0202(.A1(new_n402), .A2(KEYINPUT13), .A3(new_n399), .A4(new_n292), .ZN(new_n403));
  OAI21_X1  g0203(.A(G169), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT14), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n401), .A2(new_n403), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G179), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT14), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n408), .B(G169), .C1(new_n401), .C2(new_n403), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n405), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n370), .A2(new_n205), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT12), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n205), .B2(new_n267), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n254), .A2(G77), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n414), .B1(new_n229), .B2(G68), .C1(new_n260), .C2(new_n272), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n264), .ZN(new_n416));
  OR2_X1    g0216(.A1(new_n416), .A2(KEYINPUT11), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(KEYINPUT11), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n410), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(G200), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT70), .B1(new_n406), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n406), .A2(G190), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT70), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n425), .B(G200), .C1(new_n401), .C2(new_n403), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n419), .A2(new_n423), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n323), .A2(new_n297), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n334), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n323), .A2(G200), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n391), .A2(new_n421), .A3(new_n427), .A4(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n336), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT4), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(G1698), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(G244), .C1(new_n346), .C2(new_n345), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G283), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n322), .B1(new_n279), .B2(new_n280), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n436), .B(new_n437), .C1(new_n438), .C2(KEYINPUT4), .ZN(new_n439));
  OAI21_X1  g0239(.A(G250), .B1(new_n345), .B2(new_n346), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n282), .B1(new_n440), .B2(KEYINPUT4), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n288), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G41), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n270), .B(G45), .C1(new_n443), .C2(KEYINPUT5), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT74), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(KEYINPUT5), .ZN(new_n447));
  INV_X1    g0247(.A(G45), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n448), .A2(G1), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G41), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(KEYINPUT74), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n446), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n453), .A2(G257), .A3(new_n287), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n444), .A2(new_n445), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT74), .B1(new_n449), .B2(new_n451), .ZN(new_n456));
  OAI21_X1  g0256(.A(KEYINPUT75), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT75), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n446), .A2(new_n458), .A3(new_n452), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n287), .A2(G274), .A3(new_n447), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n442), .A2(new_n454), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT76), .B1(new_n463), .B2(new_n422), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n271), .A2(G97), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n253), .A2(G1), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n370), .A2(new_n264), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(new_n213), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n279), .A2(new_n229), .A3(new_n280), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n349), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n347), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n207), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n213), .A2(G107), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n207), .A2(G97), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT73), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(KEYINPUT6), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT6), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(KEYINPUT73), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n476), .B(new_n477), .C1(new_n479), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(KEYINPUT73), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n478), .A2(KEYINPUT6), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(G97), .A4(new_n207), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n229), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n260), .A2(new_n329), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n475), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n466), .B(new_n471), .C1(new_n488), .C2(new_n266), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n463), .A2(G190), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT76), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n462), .A2(new_n492), .A3(G200), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n464), .A2(new_n490), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n462), .A2(new_n315), .ZN(new_n495));
  INV_X1    g0295(.A(G179), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n442), .A2(new_n496), .A3(new_n461), .A4(new_n454), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n489), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n370), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT25), .B1(new_n370), .B2(new_n207), .ZN(new_n500));
  OAI22_X1  g0300(.A1(new_n469), .A2(new_n207), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n229), .A2(G33), .A3(G116), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n229), .A2(G107), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n503), .B(KEYINPUT23), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n229), .B(G87), .C1(new_n345), .C2(new_n346), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n505), .A2(KEYINPUT22), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(KEYINPUT22), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n502), .B(new_n504), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT24), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n505), .B(KEYINPUT22), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT24), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(new_n502), .A4(new_n504), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n501), .B1(new_n513), .B2(new_n264), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n220), .A2(new_n282), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n214), .A2(G1698), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n515), .B(new_n516), .C1(new_n345), .C2(new_n346), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G294), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT81), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n517), .A2(KEYINPUT81), .A3(new_n518), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n288), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n453), .A2(G264), .A3(new_n287), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n461), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n422), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n523), .A2(new_n297), .A3(new_n461), .A4(new_n524), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n514), .A2(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n494), .A2(new_n498), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n514), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n525), .A2(G169), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n523), .A2(G179), .A3(new_n461), .A4(new_n524), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n532), .A2(KEYINPUT82), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT82), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT21), .ZN(new_n537));
  OR3_X1    g0337(.A1(new_n271), .A2(KEYINPUT79), .A3(G116), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT79), .B1(new_n271), .B2(G116), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n468), .A2(G116), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n437), .B(new_n229), .C1(G33), .C2(new_n213), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n216), .A2(G20), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n264), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT20), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n541), .A2(KEYINPUT20), .A3(new_n264), .A4(new_n542), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n540), .A2(new_n547), .A3(KEYINPUT80), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT80), .B1(new_n540), .B2(new_n547), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n282), .A2(G257), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n281), .B(new_n552), .C1(new_n208), .C2(new_n282), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n553), .B(new_n288), .C1(G303), .C2(new_n281), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n453), .A2(G270), .A3(new_n287), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n461), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G169), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n537), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n550), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n548), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(KEYINPUT21), .A3(G169), .A4(new_n556), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n461), .A2(new_n554), .A3(G179), .A4(new_n555), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n556), .A2(G200), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n461), .A2(new_n554), .A3(G190), .A4(new_n555), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n551), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n558), .A2(new_n561), .A3(new_n564), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n206), .A2(new_n282), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n322), .A2(G1698), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n569), .B(new_n570), .C1(new_n345), .C2(new_n346), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G116), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n287), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n220), .B1(new_n448), .B2(G1), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n270), .A2(new_n291), .A3(G45), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n287), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT77), .B1(new_n577), .B2(new_n496), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT77), .ZN(new_n579));
  NOR4_X1   g0379(.A1(new_n573), .A2(new_n579), .A3(new_n576), .A4(G179), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n573), .A2(new_n576), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT78), .ZN(new_n583));
  XNOR2_X1  g0383(.A(new_n328), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n468), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n219), .A2(new_n213), .A3(new_n207), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n396), .A2(new_n229), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT19), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n229), .B(G68), .C1(new_n345), .C2(new_n346), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT19), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n396), .B2(G20), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n264), .B1(new_n370), .B2(new_n328), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n315), .A2(new_n582), .B1(new_n585), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(G200), .B1(new_n573), .B2(new_n576), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n468), .A2(G87), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n595), .A2(new_n593), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n577), .A2(G190), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n581), .A2(new_n594), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n568), .A2(new_n600), .ZN(new_n601));
  AND4_X1   g0401(.A1(new_n433), .A2(new_n530), .A3(new_n536), .A4(new_n601), .ZN(G372));
  INV_X1    g0402(.A(new_n318), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n387), .A2(new_n383), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n427), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n421), .B2(new_n335), .ZN(new_n607));
  INV_X1    g0407(.A(new_n377), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n374), .A2(new_n375), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n605), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n603), .B1(new_n612), .B2(new_n312), .ZN(new_n613));
  INV_X1    g0413(.A(new_n433), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n498), .A2(KEYINPUT83), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n582), .A2(new_n315), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n585), .A2(new_n593), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n577), .A2(new_n496), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n598), .A2(new_n595), .A3(new_n596), .A4(new_n593), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT83), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n489), .A2(new_n495), .A3(new_n623), .A4(new_n497), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n615), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n498), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(KEYINPUT26), .A3(new_n599), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT84), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n628), .A2(KEYINPUT84), .A3(KEYINPUT26), .A4(new_n599), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n627), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n558), .A2(new_n561), .A3(new_n564), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n514), .B1(new_n532), .B2(new_n533), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n621), .B1(new_n514), .B2(new_n528), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n494), .A2(new_n637), .A3(new_n498), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n619), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n633), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n613), .B1(new_n614), .B2(new_n640), .ZN(G369));
  INV_X1    g0441(.A(new_n536), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n232), .A2(G20), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n270), .ZN(new_n644));
  XNOR2_X1  g0444(.A(KEYINPUT85), .B(KEYINPUT27), .ZN(new_n645));
  OR2_X1    g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(G213), .A3(new_n647), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT86), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT86), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n642), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n531), .A2(new_n653), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n656), .A2(new_n529), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n655), .B1(new_n642), .B2(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT88), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT88), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n654), .A2(new_n551), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n568), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n634), .A2(new_n663), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT87), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n662), .A2(G330), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n634), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n653), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n659), .A2(new_n660), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n532), .A2(new_n533), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n531), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(new_n653), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n669), .A2(new_n672), .A3(new_n676), .ZN(G399));
  NOR2_X1   g0477(.A1(new_n233), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n586), .A2(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n228), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT89), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  INV_X1    g0484(.A(new_n619), .ZN(new_n685));
  NOR3_X1   g0485(.A1(new_n600), .A2(KEYINPUT26), .A3(new_n498), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n615), .A2(new_n620), .A3(new_n624), .ZN(new_n687));
  AOI211_X1 g0487(.A(new_n685), .B(new_n686), .C1(KEYINPUT26), .C2(new_n687), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n530), .B(new_n620), .C1(new_n642), .C2(new_n634), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n653), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n690), .A2(KEYINPUT91), .A3(KEYINPUT29), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n690), .A2(KEYINPUT29), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT91), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n654), .B1(new_n633), .B2(new_n639), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT29), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n691), .B1(new_n692), .B2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n601), .A2(new_n530), .A3(new_n536), .A4(new_n654), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n442), .A2(new_n454), .A3(new_n461), .A4(new_n577), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n523), .A2(new_n524), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  NOR4_X1   g0501(.A1(new_n699), .A2(new_n562), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n562), .A2(new_n700), .ZN(new_n703));
  INV_X1    g0503(.A(new_n699), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT30), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n556), .A2(new_n496), .A3(new_n582), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(KEYINPUT90), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT90), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n556), .A2(new_n709), .A3(new_n496), .A4(new_n582), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n462), .A2(new_n525), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n706), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n653), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(KEYINPUT31), .A3(new_n653), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n698), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(G330), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n697), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n684), .B1(new_n722), .B2(G1), .ZN(G364));
  NOR2_X1   g0523(.A1(G13), .A2(G33), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n664), .A2(new_n665), .A3(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n270), .B1(new_n643), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n678), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(KEYINPUT92), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n230), .B1(G20), .B2(new_n315), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n726), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n233), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(G355), .A3(new_n281), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n233), .A2(new_n281), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G45), .B2(new_n228), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n247), .A2(new_n448), .ZN(new_n739));
  OAI221_X1 g0539(.A(new_n736), .B1(G116), .B2(new_n735), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n732), .B1(new_n734), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT93), .Z(new_n742));
  NOR2_X1   g0542(.A1(new_n229), .A2(G179), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G190), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G159), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT32), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n219), .ZN(new_n750));
  NAND2_X1  g0550(.A1(G20), .A2(G179), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT94), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n297), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n743), .A2(new_n297), .A3(G200), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n754), .A2(new_n211), .B1(new_n207), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n496), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n750), .B(new_n756), .C1(G97), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n752), .A2(G200), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G190), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n759), .B(new_n281), .C1(new_n205), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n760), .A2(new_n297), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n748), .B(new_n763), .C1(G50), .C2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT95), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n752), .A2(new_n766), .A3(new_n744), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n766), .B1(new_n752), .B2(new_n744), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n765), .B1(new_n329), .B2(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT96), .Z(new_n771));
  INV_X1    g0571(.A(G311), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  INV_X1    g0574(.A(G329), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n755), .A2(new_n774), .B1(new_n745), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n749), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n776), .A2(KEYINPUT97), .B1(G303), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n764), .ZN(new_n779));
  INV_X1    g0579(.A(G326), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT33), .B(G317), .Z(new_n781));
  OAI221_X1 g0581(.A(new_n778), .B1(new_n779), .B2(new_n780), .C1(new_n762), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n776), .A2(KEYINPUT97), .ZN(new_n783));
  NOR3_X1   g0583(.A1(new_n782), .A2(new_n281), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n754), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G322), .ZN(new_n786));
  INV_X1    g0586(.A(G294), .ZN(new_n787));
  INV_X1    g0587(.A(new_n758), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n784), .B(new_n786), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n771), .B1(new_n773), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT98), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n728), .B(new_n742), .C1(new_n791), .C2(new_n733), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n668), .A2(G330), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n668), .A2(G330), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n794), .A2(new_n731), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(G396));
  INV_X1    g0598(.A(new_n769), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G116), .B1(G303), .B2(new_n764), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n774), .B2(new_n762), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  NOR2_X1   g0602(.A1(new_n749), .A2(new_n207), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n755), .A2(new_n219), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n785), .A2(G294), .B1(G97), .B2(new_n758), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT100), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n803), .B(new_n804), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n802), .A2(new_n347), .A3(new_n807), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n808), .B1(new_n806), .B2(new_n805), .C1(new_n772), .C2(new_n745), .ZN(new_n809));
  XNOR2_X1  g0609(.A(KEYINPUT102), .B(G143), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n799), .A2(G159), .B1(new_n785), .B2(new_n810), .ZN(new_n811));
  AOI22_X1  g0611(.A1(G137), .A2(new_n764), .B1(new_n761), .B2(G150), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n812), .A2(KEYINPUT101), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n812), .A2(KEYINPUT101), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT34), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n755), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n815), .A2(new_n816), .B1(G68), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n777), .A2(G50), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n746), .A2(G132), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n347), .B1(new_n758), .B2(G58), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n809), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n732), .B1(new_n824), .B2(new_n733), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n733), .A2(new_n724), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n335), .A2(new_n653), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n653), .A2(new_n334), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n431), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n830), .B2(new_n335), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n825), .B1(G77), .B2(new_n827), .C1(new_n725), .C2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n831), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n694), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n654), .B(new_n831), .C1(new_n633), .C2(new_n639), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(new_n720), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n832), .B1(new_n731), .B2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT103), .Z(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G384));
  NAND2_X1  g0640(.A1(new_n482), .A2(new_n485), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT104), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT35), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n229), .B(new_n230), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n844), .B(G116), .C1(new_n843), .C2(new_n842), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT36), .ZN(new_n846));
  OAI21_X1  g0646(.A(G77), .B1(new_n211), .B2(new_n205), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n228), .A2(new_n847), .B1(G50), .B2(new_n205), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(G1), .A3(new_n232), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n420), .A2(new_n653), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n421), .A2(new_n850), .A3(new_n427), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n410), .A2(new_n420), .A3(new_n653), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT105), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n494), .A2(new_n637), .A3(new_n498), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n674), .A2(new_n558), .A3(new_n561), .A4(new_n564), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n685), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n627), .A2(new_n631), .A3(new_n632), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n653), .B(new_n833), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n855), .B1(new_n860), .B2(new_n828), .ZN(new_n861));
  INV_X1    g0661(.A(new_n828), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n835), .A2(KEYINPUT105), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n854), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT106), .ZN(new_n865));
  INV_X1    g0665(.A(new_n651), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n379), .B1(new_n382), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g0667(.A(new_n865), .B(KEYINPUT37), .C1(new_n867), .C2(new_n374), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n865), .A2(KEYINPUT37), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n867), .A2(new_n374), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n379), .A2(new_n866), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n391), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n874), .B(KEYINPUT38), .C1(new_n391), .C2(new_n875), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n864), .A2(new_n880), .B1(new_n605), .B2(new_n651), .ZN(new_n881));
  INV_X1    g0681(.A(new_n879), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n386), .B1(new_n384), .B2(new_n383), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n610), .B1(new_n883), .B2(new_n389), .ZN(new_n884));
  INV_X1    g0684(.A(new_n875), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n886), .B2(new_n874), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT39), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(KEYINPUT108), .B(KEYINPUT39), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n867), .A2(new_n374), .A3(new_n871), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n869), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n872), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT107), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n608), .B2(new_n609), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n376), .A2(KEYINPUT107), .A3(new_n377), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n604), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n892), .B1(new_n896), .B2(new_n885), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n879), .B(new_n889), .C1(new_n897), .C2(KEYINPUT38), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n888), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n421), .A2(new_n653), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT109), .B1(new_n881), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n653), .B1(new_n858), .B2(new_n859), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n855), .B(new_n828), .C1(new_n903), .C2(new_n831), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT105), .B1(new_n835), .B2(new_n862), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n880), .B(new_n853), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n605), .A2(new_n651), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT109), .ZN(new_n909));
  INV_X1    g0709(.A(new_n900), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n888), .B2(new_n898), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n433), .B(new_n691), .C1(new_n692), .C2(new_n696), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n613), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n913), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n853), .A2(new_n831), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT31), .B1(new_n714), .B2(new_n653), .ZN(new_n918));
  AOI211_X1 g0718(.A(new_n716), .B(new_n654), .C1(new_n706), .C2(new_n713), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n917), .B1(new_n920), .B2(new_n698), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n880), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT40), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n923), .B1(new_n921), .B2(KEYINPUT110), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n879), .B1(new_n897), .B2(KEYINPUT38), .ZN(new_n926));
  INV_X1    g0726(.A(new_n917), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n719), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT110), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n925), .A2(new_n926), .A3(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n924), .A2(new_n433), .A3(new_n719), .A4(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n928), .B1(new_n878), .B2(new_n879), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n931), .B(G330), .C1(KEYINPUT40), .C2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n614), .A2(new_n720), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI22_X1  g0737(.A1(new_n916), .A2(new_n937), .B1(new_n270), .B2(new_n643), .ZN(new_n938));
  XOR2_X1   g0738(.A(new_n938), .B(KEYINPUT111), .Z(new_n939));
  AND2_X1   g0739(.A1(new_n916), .A2(new_n937), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n846), .B(new_n849), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT112), .Z(G367));
  INV_X1    g0742(.A(G317), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n347), .B1(new_n745), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n761), .A2(G294), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n755), .A2(new_n213), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n758), .A2(G107), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n785), .A2(G303), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n945), .A2(new_n947), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n944), .B(new_n950), .C1(G311), .C2(new_n764), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n777), .A2(G116), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT46), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n951), .B(new_n953), .C1(new_n774), .C2(new_n769), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT113), .Z(new_n955));
  NAND2_X1  g0755(.A1(new_n758), .A2(G68), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n211), .B2(new_n749), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n347), .B(new_n957), .C1(new_n761), .C2(G159), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n746), .A2(G137), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n754), .A2(new_n261), .B1(new_n329), .B2(new_n755), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(new_n764), .C2(new_n810), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n958), .B(new_n961), .C1(new_n272), .C2(new_n769), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n955), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT47), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n964), .A2(new_n733), .ZN(new_n965));
  INV_X1    g0765(.A(new_n732), .ZN(new_n966));
  INV_X1    g0766(.A(new_n737), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n734), .B1(new_n735), .B2(new_n328), .C1(new_n243), .C2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n593), .A2(new_n596), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n653), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n622), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n653), .A2(new_n685), .A3(new_n969), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n726), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n966), .B(new_n968), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n965), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n678), .B(KEYINPUT41), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n494), .A2(new_n498), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n490), .B2(new_n654), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n628), .A2(new_n653), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(new_n672), .B2(new_n676), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT44), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n672), .A2(new_n676), .A3(new_n981), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n983), .A2(new_n669), .A3(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n793), .A2(new_n661), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n669), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n671), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n669), .B(new_n989), .C1(new_n670), .C2(new_n653), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n722), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n669), .B1(new_n983), .B2(new_n986), .ZN(new_n995));
  NOR3_X1   g0795(.A1(new_n988), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n977), .B1(new_n996), .B2(new_n721), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n729), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n662), .A2(new_n978), .A3(new_n671), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n498), .B1(new_n979), .B2(new_n536), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n654), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(KEYINPUT42), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1006), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n981), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n1009), .A2(new_n1010), .B1(new_n669), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1010), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n669), .A2(new_n1011), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(new_n1014), .A3(new_n1008), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n976), .B1(new_n998), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(G387));
  NAND2_X1  g0819(.A1(new_n993), .A2(new_n730), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT114), .ZN(new_n1021));
  XOR2_X1   g0821(.A(KEYINPUT117), .B(G322), .Z(new_n1022));
  AOI22_X1  g0822(.A1(new_n764), .A2(new_n1022), .B1(new_n785), .B2(G317), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n772), .B2(new_n762), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G303), .B2(new_n799), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT48), .Z(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n774), .B2(new_n788), .C1(new_n787), .C2(new_n749), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT49), .Z(new_n1028));
  OAI221_X1 g0828(.A(new_n347), .B1(new_n745), .B2(new_n780), .C1(new_n216), .C2(new_n755), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT118), .Z(new_n1030));
  OAI221_X1 g0830(.A(new_n947), .B1(new_n779), .B2(new_n342), .C1(new_n256), .C2(new_n762), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n584), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(new_n788), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n754), .A2(new_n272), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n745), .A2(new_n261), .ZN(new_n1035));
  NOR4_X1   g0835(.A1(new_n1033), .A2(new_n1034), .A3(new_n347), .A4(new_n1035), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n1036), .B1(new_n205), .B2(new_n769), .C1(new_n329), .C2(new_n749), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1028), .A2(new_n1030), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n732), .B1(new_n1038), .B2(new_n733), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n734), .ZN(new_n1040));
  OR3_X1    g0840(.A1(new_n256), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1041));
  OAI21_X1  g0841(.A(KEYINPUT50), .B1(new_n256), .B2(G50), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1041), .A2(new_n1042), .A3(new_n448), .A4(new_n680), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n205), .A2(new_n329), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n737), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT115), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n448), .B2(new_n240), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n735), .A2(new_n281), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1047), .B1(G107), .B2(new_n735), .C1(new_n680), .C2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT116), .Z(new_n1050));
  OAI221_X1 g0850(.A(new_n1039), .B1(new_n662), .B2(new_n974), .C1(new_n1040), .C2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1021), .A2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n993), .B(new_n721), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n678), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(G393));
  INV_X1    g0857(.A(new_n995), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1058), .A2(new_n730), .A3(new_n987), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n734), .B1(new_n967), .B2(new_n250), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(G97), .B2(new_n233), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n769), .A2(new_n787), .B1(new_n207), .B2(new_n755), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n764), .A2(G317), .B1(new_n785), .B2(G311), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT52), .Z(new_n1064));
  NAND2_X1  g0864(.A1(new_n746), .A2(new_n1022), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n347), .A3(new_n1065), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1062), .B(new_n1066), .C1(G303), .C2(new_n761), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n216), .B2(new_n788), .C1(new_n774), .C2(new_n749), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n764), .A2(G150), .B1(new_n785), .B2(G159), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT51), .Z(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n329), .B2(new_n788), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n347), .B(new_n1071), .C1(G50), .C2(new_n761), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n749), .A2(new_n205), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n804), .B(new_n1073), .C1(new_n746), .C2(new_n810), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1072), .B(new_n1074), .C1(new_n256), .C2(new_n769), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1068), .A2(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n732), .B(new_n1061), .C1(new_n1076), .C2(new_n733), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n974), .B2(new_n981), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1059), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1058), .A2(new_n987), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n679), .B1(new_n1080), .B2(new_n994), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n996), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(G390));
  OAI211_X1 g0884(.A(new_n914), .B(new_n613), .C1(new_n614), .C2(new_n720), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n720), .A2(new_n917), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n719), .A2(G330), .A3(new_n831), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(KEYINPUT120), .A3(new_n854), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(KEYINPUT120), .B1(new_n1088), .B2(new_n854), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n1090), .A2(new_n1091), .B1(new_n905), .B2(new_n904), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n830), .A2(new_n335), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n653), .B(new_n1094), .C1(new_n688), .C2(new_n689), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1095), .A2(new_n828), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n853), .B(KEYINPUT119), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1088), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1087), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1085), .B1(new_n1092), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n853), .B1(new_n904), .B2(new_n905), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n899), .B1(new_n910), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1097), .B1(new_n1095), .B2(new_n828), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1104), .A2(new_n910), .A3(new_n926), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1086), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n888), .B(new_n898), .C1(new_n864), .C2(new_n900), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1108), .A2(new_n1105), .A3(new_n1087), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1101), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n678), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1101), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n777), .A2(G150), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT53), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n785), .A2(G132), .ZN(new_n1117));
  INV_X1    g0917(.A(G128), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1117), .B1(new_n272), .B2(new_n755), .C1(new_n779), .C2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT54), .B(G143), .Z(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n799), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n347), .B1(new_n761), .B2(G137), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1121), .B(new_n1122), .C1(new_n342), .C2(new_n788), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1116), .B(new_n1123), .C1(G125), .C2(new_n746), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n754), .A2(new_n216), .B1(new_n205), .B2(new_n755), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n799), .B2(G97), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n329), .B2(new_n788), .C1(new_n774), .C2(new_n779), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n347), .B1(new_n787), .B2(new_n745), .C1(new_n762), .C2(new_n207), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n1127), .A2(new_n750), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n733), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1130), .A2(new_n966), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n372), .B2(new_n827), .C1(new_n899), .C2(new_n725), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1112), .B2(new_n729), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1114), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(G378));
  INV_X1    g0935(.A(KEYINPUT57), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1103), .A2(new_n1106), .A3(new_n1086), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1087), .B1(new_n1108), .B2(new_n1105), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1085), .B1(new_n1139), .B2(new_n1101), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n866), .A2(new_n276), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT121), .Z(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  XOR2_X1   g0943(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n312), .A2(new_n318), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n312), .B2(new_n318), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1143), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n312), .A2(new_n318), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1144), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1151), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1152));
  AND2_X1   g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n934), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n924), .A2(new_n1155), .A3(G330), .A4(new_n931), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n902), .B2(new_n912), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n909), .B1(new_n908), .B2(new_n911), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n901), .A2(KEYINPUT109), .A3(new_n907), .A4(new_n906), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n1156), .A4(new_n1154), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1136), .B1(new_n1140), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1085), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1110), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1165), .A2(KEYINPUT57), .A3(new_n1161), .A4(new_n1158), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1163), .A2(new_n678), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1158), .A2(new_n730), .A3(new_n1161), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n731), .B1(G50), .B2(new_n827), .ZN(new_n1169));
  INV_X1    g0969(.A(G124), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n253), .B1(new_n745), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n799), .A2(G137), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n761), .A2(G132), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n777), .A2(new_n1120), .B1(new_n758), .B2(G150), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n764), .A2(G125), .B1(new_n785), .B2(G128), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  AOI211_X1 g0976(.A(G41), .B(new_n1171), .C1(new_n1176), .C2(KEYINPUT59), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(KEYINPUT59), .B2(new_n1176), .C1(new_n342), .C2(new_n755), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n347), .B1(new_n207), .B2(new_n754), .C1(new_n769), .C2(new_n1032), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n761), .A2(G97), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n764), .A2(G116), .ZN(new_n1181));
  AOI21_X1  g0981(.A(G41), .B1(new_n746), .B2(G283), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n956), .A4(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n749), .A2(new_n329), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n755), .A2(new_n211), .ZN(new_n1185));
  NOR4_X1   g0985(.A1(new_n1179), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT58), .Z(new_n1187));
  OAI21_X1  g0987(.A(new_n272), .B1(new_n345), .B2(G41), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1178), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1169), .B1(new_n1189), .B2(new_n733), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n1155), .B2(new_n725), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n1168), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1167), .A2(new_n1192), .ZN(G375));
  NOR2_X1   g0993(.A1(new_n779), .A2(new_n787), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1033), .B1(G97), .B2(new_n777), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n799), .A2(G107), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n761), .A2(G116), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n755), .A2(new_n329), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n281), .B(new_n1198), .C1(G303), .C2(new_n746), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1194), .B(new_n1200), .C1(G283), .C2(new_n785), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n749), .A2(new_n342), .B1(new_n745), .B2(new_n1118), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT122), .Z(new_n1203));
  NAND2_X1  g1003(.A1(new_n799), .A2(G150), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n761), .A2(new_n1120), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1185), .B1(new_n764), .B2(G132), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n347), .B1(new_n785), .B2(G137), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1203), .B(new_n1208), .C1(G50), .C2(new_n758), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n733), .B1(new_n1201), .B2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n1210), .B(new_n966), .C1(G68), .C2(new_n827), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1098), .B2(new_n724), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1092), .A2(new_n1100), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(new_n1213), .B2(new_n730), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1085), .A2(new_n1092), .A3(new_n1100), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n977), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1214), .B1(new_n1216), .B2(new_n1101), .ZN(G381));
  NAND3_X1  g1017(.A1(new_n1167), .A2(new_n1134), .A3(new_n1192), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1054), .A2(new_n1021), .A3(new_n797), .A4(new_n1051), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(G384), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1218), .B1(KEYINPUT123), .B2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(G390), .A2(G381), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1220), .A2(KEYINPUT123), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1221), .A2(new_n1018), .A3(new_n1222), .A4(new_n1223), .ZN(G407));
  OAI211_X1 g1024(.A(G407), .B(G213), .C1(G343), .C2(new_n1218), .ZN(G409));
  NAND2_X1  g1025(.A1(G375), .A2(G378), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT124), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1158), .A2(new_n1227), .A3(new_n1161), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n730), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1227), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1191), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT125), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1165), .A2(new_n977), .A3(new_n1161), .A4(new_n1158), .ZN(new_n1234));
  OAI211_X1 g1034(.A(KEYINPUT125), .B(new_n1191), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1233), .A2(new_n1134), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n652), .A2(G213), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT60), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n679), .B1(new_n1215), .B2(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1239), .B(new_n1113), .C1(new_n1238), .C2(new_n1215), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n1214), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(G384), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n839), .A2(new_n1214), .A3(new_n1240), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1226), .A2(new_n1236), .A3(new_n1237), .A4(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(KEYINPUT126), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT63), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1226), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n652), .A2(G213), .A3(G2897), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1244), .B(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT61), .B1(new_n1248), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT63), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1245), .A2(KEYINPUT126), .A3(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT127), .B1(new_n1018), .B2(G390), .ZN(new_n1255));
  OAI21_X1  g1055(.A(G396), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1219), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1016), .B1(new_n997), .B2(new_n729), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1083), .B1(new_n1259), .B2(new_n976), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n998), .A2(new_n1017), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n976), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1261), .A2(G390), .A3(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1258), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT127), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1260), .A2(new_n1263), .A3(new_n1266), .A4(new_n1257), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1247), .A2(new_n1252), .A3(new_n1254), .A4(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1245), .A2(KEYINPUT62), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G375), .A2(G378), .B1(G213), .B2(new_n652), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1236), .A4(new_n1244), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1267), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1255), .A2(new_n1257), .B1(new_n1263), .B2(new_n1260), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1276), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1269), .A2(new_n1280), .ZN(G405));
  NAND2_X1  g1081(.A1(new_n1226), .A2(new_n1218), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n1243), .A3(new_n1242), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1226), .A2(new_n1218), .A3(new_n1244), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1279), .ZN(G402));
endmodule


