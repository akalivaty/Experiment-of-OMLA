//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  NOR2_X1   g001(.A1(G472), .A2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT30), .ZN(new_n190));
  INV_X1    g004(.A(G131), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G134), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(G137), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G137), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n196), .B1(new_n193), .B2(G137), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n191), .B(new_n194), .C1(new_n197), .C2(new_n192), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n193), .A2(G137), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G134), .ZN(new_n201));
  OAI21_X1  g015(.A(G131), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(KEYINPUT1), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n207), .A2(KEYINPUT64), .A3(G146), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT64), .B1(new_n207), .B2(G146), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n204), .B(new_n206), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(G143), .B2(new_n203), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n207), .A2(G146), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n203), .A2(G143), .ZN(new_n214));
  OAI22_X1  g028(.A1(new_n212), .A2(new_n205), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n198), .A2(new_n202), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n203), .B2(G143), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n207), .A2(KEYINPUT64), .A3(G146), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n213), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT0), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(new_n205), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n207), .A2(G146), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n204), .A2(new_n225), .B1(KEYINPUT0), .B2(G128), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n205), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g043(.A1(KEYINPUT65), .A2(G134), .ZN(new_n230));
  NOR2_X1   g044(.A1(KEYINPUT65), .A2(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(G137), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n196), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n192), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n230), .A2(new_n231), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT11), .B1(new_n235), .B2(new_n200), .ZN(new_n236));
  OAI21_X1  g050(.A(G131), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n229), .B1(new_n237), .B2(new_n198), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n190), .B1(new_n217), .B2(new_n238), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n223), .A2(new_n221), .B1(new_n226), .B2(new_n227), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n234), .A2(new_n236), .A3(G131), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n195), .ZN(new_n243));
  NAND2_X1  g057(.A1(KEYINPUT65), .A2(G134), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n200), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT11), .B1(new_n245), .B2(new_n196), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n191), .B1(new_n246), .B2(new_n194), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n240), .B1(new_n241), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n210), .A2(new_n249), .A3(new_n215), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n210), .B2(new_n215), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n198), .B(new_n202), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n248), .A2(new_n252), .A3(KEYINPUT30), .ZN(new_n253));
  INV_X1    g067(.A(G119), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G116), .ZN(new_n255));
  INV_X1    g069(.A(G116), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G119), .ZN(new_n257));
  INV_X1    g071(.A(G113), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n258), .A2(KEYINPUT2), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(KEYINPUT2), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n255), .B(new_n257), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n255), .A2(new_n257), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT2), .B(G113), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n264), .A3(KEYINPUT66), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n262), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n239), .A2(new_n253), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n265), .A2(KEYINPUT68), .A3(new_n267), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(new_n248), .A3(new_n252), .ZN(new_n275));
  INV_X1    g089(.A(G237), .ZN(new_n276));
  INV_X1    g090(.A(G953), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(G210), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n278), .B(G101), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n270), .A2(new_n275), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n270), .A2(KEYINPUT31), .A3(new_n275), .A4(new_n281), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n269), .B1(new_n217), .B2(new_n238), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n275), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT28), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT28), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n275), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n281), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n189), .B1(new_n286), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n187), .B1(new_n295), .B2(KEYINPUT32), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n284), .A2(new_n285), .B1(new_n292), .B2(new_n293), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT32), .ZN(new_n298));
  NOR4_X1   g112(.A1(new_n297), .A2(KEYINPUT72), .A3(new_n298), .A4(new_n189), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n270), .A2(new_n275), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n293), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT70), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(KEYINPUT70), .A3(new_n293), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n289), .A2(KEYINPUT69), .A3(new_n281), .A4(new_n291), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n289), .A2(new_n281), .A3(new_n291), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT69), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT29), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n301), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n198), .A2(new_n202), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n216), .A2(KEYINPUT67), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n210), .A2(new_n215), .A3(new_n249), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n237), .A2(new_n198), .ZN(new_n319));
  AOI22_X1  g133(.A1(new_n315), .A2(new_n318), .B1(new_n319), .B2(new_n240), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(new_n274), .ZN(new_n321));
  INV_X1    g135(.A(new_n275), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT28), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n323), .A2(KEYINPUT29), .A3(new_n281), .A4(new_n291), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT71), .ZN(new_n325));
  OAI21_X1  g139(.A(G472), .B1(new_n314), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n298), .B1(new_n297), .B2(new_n189), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n300), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n254), .A2(G128), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT23), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n205), .A2(G119), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n330), .B1(new_n333), .B2(new_n329), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G110), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n331), .A2(new_n329), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT24), .B(G110), .Z(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G140), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G125), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT16), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G140), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(KEYINPUT73), .A3(G140), .ZN(new_n348));
  AOI22_X1  g162(.A1(new_n347), .A2(new_n348), .B1(G125), .B2(new_n340), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n343), .B1(new_n349), .B2(new_n342), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G146), .ZN(new_n351));
  INV_X1    g165(.A(new_n343), .ZN(new_n352));
  INV_X1    g166(.A(new_n348), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT73), .B1(new_n344), .B2(G140), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n341), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n352), .B1(new_n355), .B2(KEYINPUT16), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n203), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n339), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n341), .A2(new_n345), .A3(new_n203), .ZN(new_n360));
  OAI22_X1  g174(.A1(new_n334), .A2(G110), .B1(new_n336), .B2(new_n337), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n351), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n277), .A2(G221), .A3(G234), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT74), .ZN(new_n364));
  XOR2_X1   g178(.A(KEYINPUT22), .B(G137), .Z(new_n365));
  XNOR2_X1  g179(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n359), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n366), .ZN(new_n368));
  INV_X1    g182(.A(new_n362), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(new_n358), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n371), .A2(KEYINPUT75), .ZN(new_n372));
  INV_X1    g186(.A(G217), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(G234), .B2(new_n301), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(G902), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(KEYINPUT75), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n372), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT76), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n371), .A2(KEYINPUT25), .A3(new_n301), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT25), .B1(new_n371), .B2(new_n301), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n374), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n372), .A2(new_n382), .A3(new_n375), .A4(new_n376), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n378), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n328), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G469), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n388));
  INV_X1    g202(.A(G104), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT3), .B1(new_n389), .B2(G107), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G104), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n389), .A2(G107), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n390), .A2(new_n393), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n389), .A2(G107), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n392), .A2(G104), .ZN(new_n398));
  OAI21_X1  g212(.A(G101), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n396), .A2(new_n399), .A3(KEYINPUT10), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n250), .B2(new_n251), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT80), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n318), .A2(KEYINPUT80), .A3(new_n400), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n319), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT79), .B(KEYINPUT10), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n212), .A2(new_n205), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n210), .B1(new_n221), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n396), .A2(new_n399), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n390), .A2(new_n393), .A3(new_n395), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G101), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT4), .A3(new_n396), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n415), .A3(G101), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n411), .B1(new_n417), .B2(new_n240), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n405), .A2(KEYINPUT81), .A3(new_n406), .A4(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n418), .A2(new_n403), .A3(new_n404), .A4(new_n406), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT81), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(G110), .B(G140), .ZN(new_n424));
  INV_X1    g238(.A(G227), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(G953), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n424), .B(new_n426), .Z(new_n427));
  AOI21_X1  g241(.A(new_n388), .B1(new_n423), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n427), .ZN(new_n429));
  AOI211_X1 g243(.A(KEYINPUT83), .B(new_n429), .C1(new_n419), .C2(new_n422), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n409), .A2(new_n410), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n216), .B2(new_n410), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n432), .A2(new_n319), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n433), .A2(KEYINPUT12), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(KEYINPUT82), .A3(KEYINPUT12), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(KEYINPUT12), .A3(new_n319), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n434), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n428), .A2(new_n430), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n405), .A2(new_n418), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n319), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n427), .B1(new_n423), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n387), .B(new_n301), .C1(new_n441), .C2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n387), .A2(new_n301), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n427), .B1(new_n423), .B2(new_n439), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n423), .A2(new_n427), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n447), .B1(new_n449), .B2(new_n443), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n446), .B1(new_n450), .B2(G469), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n276), .A2(new_n277), .A3(G214), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n207), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n276), .A2(new_n277), .A3(G143), .A4(G214), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(KEYINPUT18), .A2(G131), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n360), .B1(new_n349), .B2(new_n203), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT17), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n454), .A2(new_n191), .A3(new_n455), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT87), .B1(new_n456), .B2(G131), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT87), .ZN(new_n464));
  AOI211_X1 g278(.A(new_n464), .B(new_n191), .C1(new_n454), .C2(new_n455), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n461), .B(new_n462), .C1(new_n463), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n456), .A2(G131), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n464), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n456), .A2(KEYINPUT87), .A3(G131), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(KEYINPUT17), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n351), .A2(new_n357), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n460), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(G113), .B(G122), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(new_n389), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT19), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n341), .A2(new_n345), .A3(new_n477), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n203), .B(new_n478), .C1(new_n349), .C2(new_n477), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n356), .B2(new_n203), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n462), .B1(new_n463), .B2(new_n465), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n351), .A2(KEYINPUT88), .A3(new_n479), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n475), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(new_n460), .ZN(new_n487));
  NOR2_X1   g301(.A1(G475), .A2(G902), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n476), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT20), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT89), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(KEYINPUT89), .A3(KEYINPUT20), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n476), .A2(new_n487), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT20), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT90), .B1(G475), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT90), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n488), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n492), .A2(new_n493), .A3(new_n499), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n475), .A2(KEYINPUT91), .ZN(new_n501));
  AOI21_X1  g315(.A(G902), .B1(new_n473), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n473), .B2(new_n501), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G475), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(G128), .B(G143), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n193), .B(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G122), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G116), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n256), .A2(G122), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n392), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT14), .B1(new_n508), .B2(G116), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT92), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OR3_X1    g329(.A1(new_n508), .A2(KEYINPUT14), .A3(G116), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(KEYINPUT92), .A3(KEYINPUT14), .ZN(new_n517));
  AND4_X1   g331(.A1(new_n509), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n507), .B(new_n512), .C1(new_n518), .C2(new_n392), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n511), .B(new_n392), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n506), .A2(KEYINPUT13), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n207), .A2(G128), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n521), .B(G134), .C1(KEYINPUT13), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n193), .A2(new_n506), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT9), .B(G234), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n527), .B(KEYINPUT77), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(G217), .A3(new_n277), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n526), .B(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G478), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n530), .B(new_n301), .C1(KEYINPUT15), .C2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n526), .A2(G217), .A3(new_n277), .A4(new_n528), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n519), .A2(new_n525), .A3(new_n529), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n301), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT15), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(G478), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT93), .ZN(new_n539));
  OR2_X1    g353(.A1(KEYINPUT94), .A2(G952), .ZN(new_n540));
  NAND2_X1  g354(.A1(KEYINPUT94), .A2(G952), .ZN(new_n541));
  AOI21_X1  g355(.A(G953), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G234), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n276), .ZN(new_n544));
  OAI211_X1 g358(.A(G902), .B(G953), .C1(new_n543), .C2(new_n276), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n545), .B(KEYINPUT95), .Z(new_n546));
  XOR2_X1   g360(.A(KEYINPUT21), .B(G898), .Z(new_n547));
  OAI21_X1  g361(.A(new_n544), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n505), .A2(new_n539), .A3(new_n549), .ZN(new_n550));
  MUX2_X1   g364(.A(new_n216), .B(new_n240), .S(G125), .Z(new_n551));
  NAND2_X1  g365(.A1(new_n277), .A2(G224), .ZN(new_n552));
  XOR2_X1   g366(.A(new_n552), .B(KEYINPUT85), .Z(new_n553));
  XNOR2_X1  g367(.A(new_n551), .B(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n414), .A2(new_n267), .A3(new_n265), .A4(new_n416), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n255), .A2(new_n257), .A3(KEYINPUT5), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n556), .B(G113), .C1(KEYINPUT5), .C2(new_n255), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n410), .A2(new_n261), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(G110), .B(G122), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n555), .A2(new_n558), .A3(new_n560), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(KEYINPUT6), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT84), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT6), .ZN(new_n566));
  AND4_X1   g380(.A1(new_n565), .A2(new_n559), .A3(new_n566), .A4(new_n561), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n560), .B1(new_n555), .B2(new_n558), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n565), .B1(new_n568), .B2(new_n566), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n554), .B(new_n564), .C1(new_n567), .C2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT86), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n410), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n557), .A2(new_n261), .ZN(new_n573));
  OR2_X1    g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n560), .B(KEYINPUT8), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n552), .A2(KEYINPUT7), .ZN(new_n578));
  OR2_X1    g392(.A1(new_n551), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n551), .A2(new_n578), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n577), .A2(new_n563), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n570), .A2(new_n301), .A3(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(G210), .B1(G237), .B2(G902), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n570), .A2(new_n301), .A3(new_n583), .A4(new_n581), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G214), .B1(G237), .B2(G902), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n528), .A2(new_n301), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G221), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(KEYINPUT78), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n452), .A2(new_n550), .A3(new_n590), .A4(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n386), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(new_n394), .ZN(G3));
  INV_X1    g410(.A(new_n593), .ZN(new_n597));
  INV_X1    g411(.A(new_n295), .ZN(new_n598));
  OAI21_X1  g412(.A(G472), .B1(new_n297), .B2(G902), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI211_X1 g414(.A(new_n597), .B(new_n600), .C1(new_n445), .C2(new_n451), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n585), .A2(new_n586), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n602), .B1(new_n603), .B2(new_n588), .ZN(new_n604));
  AOI211_X1 g418(.A(KEYINPUT96), .B(new_n589), .C1(new_n585), .C2(new_n586), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n529), .A2(KEYINPUT98), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n526), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT33), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n530), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n531), .A2(G902), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n612), .A2(new_n613), .B1(new_n531), .B2(new_n535), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n500), .B2(new_n504), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n615), .A2(new_n548), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n601), .A2(new_n385), .A3(new_n606), .A4(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT34), .B(G104), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  NAND3_X1  g433(.A1(new_n494), .A2(new_n495), .A3(new_n488), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n492), .A2(new_n493), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n539), .A2(new_n621), .A3(new_n504), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(new_n385), .A3(new_n548), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n601), .A2(new_n606), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT35), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(new_n392), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n626), .B(new_n628), .ZN(G9));
  NAND2_X1  g443(.A1(new_n359), .A2(new_n362), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n366), .A2(KEYINPUT36), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n375), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n381), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n600), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n594), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT37), .B(G110), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  OAI21_X1  g454(.A(new_n544), .B1(new_n546), .B2(G900), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n539), .A2(new_n621), .A3(new_n504), .A4(new_n641), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n642), .A2(new_n604), .A3(new_n605), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n597), .B1(new_n445), .B2(new_n451), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n328), .A2(new_n643), .A3(new_n644), .A4(new_n634), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  NOR2_X1   g460(.A1(new_n295), .A2(KEYINPUT32), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n296), .A2(new_n299), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(G472), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n293), .B1(new_n321), .B2(new_n322), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n650), .A2(new_n282), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n651), .A2(KEYINPUT101), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(KEYINPUT101), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n652), .A2(new_n653), .A3(G902), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n648), .B1(new_n649), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT102), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n505), .A2(new_n539), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n588), .A3(new_n635), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n658), .B(KEYINPUT103), .Z(new_n659));
  NOR2_X1   g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n641), .B(KEYINPUT39), .Z(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n644), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT40), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n603), .B(KEYINPUT38), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n660), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  AND3_X1   g481(.A1(new_n328), .A2(new_n644), .A3(new_n634), .ZN(new_n668));
  INV_X1    g482(.A(new_n641), .ZN(new_n669));
  AOI211_X1 g483(.A(new_n669), .B(new_n614), .C1(new_n500), .C2(new_n504), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT104), .B1(new_n606), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n614), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n505), .A2(new_n672), .A3(new_n641), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n674));
  NOR4_X1   g488(.A1(new_n673), .A2(new_n604), .A3(new_n605), .A4(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n668), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  NOR2_X1   g491(.A1(new_n428), .A2(new_n430), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n444), .B1(new_n678), .B2(new_n439), .ZN(new_n679));
  OAI21_X1  g493(.A(G469), .B1(new_n679), .B2(G902), .ZN(new_n680));
  AND4_X1   g494(.A1(new_n592), .A2(new_n680), .A3(new_n606), .A4(new_n445), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n384), .B1(new_n648), .B2(new_n326), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n616), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  NAND2_X1  g499(.A1(new_n448), .A2(KEYINPUT83), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n423), .A2(new_n388), .A3(new_n427), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n439), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n444), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n387), .B1(new_n690), .B2(new_n301), .ZN(new_n691));
  AOI211_X1 g505(.A(G469), .B(G902), .C1(new_n688), .C2(new_n689), .ZN(new_n692));
  INV_X1    g506(.A(new_n592), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n694), .A2(new_n328), .A3(new_n624), .A4(new_n606), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT105), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n680), .A2(new_n606), .A3(new_n592), .A4(new_n445), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n286), .A2(new_n294), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(KEYINPUT32), .A3(new_n188), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT72), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n295), .A2(new_n187), .A3(KEYINPUT32), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n327), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n290), .B1(new_n275), .B2(new_n287), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT28), .B1(new_n320), .B2(new_n274), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n703), .A2(new_n704), .A3(new_n310), .A4(new_n293), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT70), .B1(new_n302), .B2(new_n293), .ZN(new_n706));
  AOI211_X1 g520(.A(new_n304), .B(new_n281), .C1(new_n270), .C2(new_n275), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(KEYINPUT29), .B1(new_n309), .B2(new_n310), .ZN(new_n709));
  AOI21_X1  g523(.A(G902), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n324), .B(KEYINPUT71), .Z(new_n711));
  AOI21_X1  g525(.A(new_n649), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n702), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n697), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n715), .A3(new_n624), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n696), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  NAND4_X1  g532(.A1(new_n681), .A2(new_n328), .A3(new_n550), .A4(new_n634), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  AND2_X1   g534(.A1(new_n323), .A2(new_n291), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n286), .B1(new_n721), .B2(new_n281), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n188), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n723), .A2(new_n599), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n657), .A2(new_n724), .A3(new_n385), .A4(new_n548), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n697), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  NOR2_X1   g541(.A1(new_n691), .A2(new_n692), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n723), .A2(new_n599), .A3(new_n634), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n673), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n728), .A2(new_n592), .A3(new_n606), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  NAND2_X1  g546(.A1(new_n699), .A2(new_n327), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT106), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n699), .A2(new_n327), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n326), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n587), .A2(new_n588), .A3(new_n592), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n445), .B2(new_n451), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(new_n739), .A3(new_n385), .A4(new_n670), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT42), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n673), .A2(KEYINPUT42), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n682), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT107), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n741), .A2(new_n743), .A3(KEYINPUT107), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G131), .ZN(G33));
  INV_X1    g563(.A(new_n642), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n328), .A2(new_n739), .A3(new_n385), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  NAND3_X1  g566(.A1(new_n500), .A2(new_n504), .A3(new_n672), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n753), .A2(new_n754), .A3(KEYINPUT43), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n600), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n635), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(KEYINPUT44), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n587), .A2(new_n588), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n757), .A2(new_n761), .A3(new_n758), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n762), .A2(new_n764), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n423), .A2(new_n443), .A3(new_n427), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n423), .A2(new_n439), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n771), .B1(new_n772), .B2(new_n427), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(KEYINPUT45), .B(new_n771), .C1(new_n772), .C2(new_n427), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(G469), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n446), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(KEYINPUT46), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n445), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT46), .B1(new_n777), .B2(new_n778), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n592), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n762), .A2(KEYINPUT109), .A3(new_n764), .A4(new_n767), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n770), .A2(new_n662), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G137), .ZN(G39));
  NAND2_X1  g600(.A1(new_n782), .A2(KEYINPUT47), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n788), .B(new_n592), .C1(new_n780), .C2(new_n781), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n328), .A2(new_n385), .A3(new_n763), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n787), .A2(new_n670), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT110), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  INV_X1    g607(.A(new_n665), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n680), .A2(new_n445), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n385), .B(new_n794), .C1(new_n795), .C2(KEYINPUT49), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n753), .B(new_n796), .C1(KEYINPUT49), .C2(new_n795), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(new_n588), .A3(new_n593), .A4(new_n656), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n694), .A2(new_n589), .A3(new_n794), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT116), .Z(new_n800));
  NAND2_X1  g614(.A1(new_n724), .A2(new_n385), .ZN(new_n801));
  INV_X1    g615(.A(new_n544), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n759), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT115), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n759), .A2(new_n805), .A3(new_n802), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n801), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n800), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n800), .A2(KEYINPUT50), .A3(new_n807), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n787), .A2(new_n789), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n795), .A2(new_n593), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n807), .B(new_n764), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n795), .B(new_n738), .C1(new_n804), .C2(new_n806), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n634), .A3(new_n724), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n795), .A2(new_n738), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n656), .A2(new_n385), .A3(new_n802), .A4(new_n818), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n819), .A2(new_n505), .A3(new_n672), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n812), .A2(new_n815), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT51), .B1(new_n815), .B2(KEYINPUT117), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n542), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n822), .B2(new_n821), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n807), .A2(new_n681), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n675), .A2(new_n671), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n328), .A2(new_n644), .A3(new_n634), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n645), .B(new_n731), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n381), .A2(new_n633), .A3(new_n641), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT113), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n445), .B2(new_n451), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n606), .A2(new_n657), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n655), .A3(new_n592), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n826), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n731), .A2(new_n645), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n676), .A3(KEYINPUT52), .A4(new_n834), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT114), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n676), .A3(new_n834), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n840), .B1(new_n841), .B2(new_n826), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n719), .A2(new_n683), .A3(new_n726), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n716), .B2(new_n696), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n621), .A2(new_n504), .A3(new_n537), .A4(new_n532), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n763), .A3(new_n669), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n328), .A2(new_n644), .A3(new_n849), .A4(new_n634), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n739), .A2(new_n730), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n751), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n594), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n682), .B2(new_n636), .ZN(new_n854));
  INV_X1    g668(.A(new_n590), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n500), .A2(new_n504), .A3(new_n538), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT111), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n856), .B1(new_n615), .B2(new_n857), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(new_n601), .A3(new_n385), .A4(new_n548), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n852), .A2(new_n854), .A3(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n846), .A2(new_n748), .A3(new_n847), .A4(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n616), .B(new_n385), .C1(new_n702), .C2(new_n712), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n697), .B1(new_n864), .B2(new_n725), .ZN(new_n865));
  INV_X1    g679(.A(new_n550), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n697), .A2(new_n713), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n865), .B1(new_n634), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n858), .A2(new_n859), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n590), .A3(new_n548), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n644), .A2(new_n385), .A3(new_n760), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n594), .B1(new_n386), .B2(new_n637), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n717), .A2(new_n868), .A3(new_n874), .A4(new_n852), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n741), .A2(new_n743), .A3(KEYINPUT107), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT107), .B1(new_n741), .B2(new_n743), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT112), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n843), .A2(new_n844), .A3(new_n863), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n836), .A2(new_n838), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n863), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n880), .B(KEYINPUT54), .C1(new_n844), .C2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n865), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n715), .B1(new_n714), .B2(new_n624), .ZN(new_n886));
  NOR4_X1   g700(.A1(new_n697), .A2(new_n713), .A3(KEYINPUT105), .A4(new_n623), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n719), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n751), .A2(new_n850), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(new_n854), .A3(new_n861), .A4(new_n851), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n888), .A2(new_n890), .A3(new_n744), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n891), .B(KEYINPUT53), .C1(new_n839), .C2(new_n842), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n844), .B2(new_n882), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n824), .A2(new_n825), .A3(new_n884), .A4(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n615), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n819), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n816), .A2(new_n385), .A3(new_n737), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(KEYINPUT48), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n900), .B(new_n902), .Z(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n901), .B2(KEYINPUT48), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n897), .A2(new_n899), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n798), .B1(new_n905), .B2(new_n906), .ZN(G75));
  NOR2_X1   g721(.A1(new_n277), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(new_n894), .B2(new_n301), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n882), .A2(new_n844), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n301), .B1(new_n912), .B2(new_n892), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT120), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n583), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n564), .B1(new_n567), .B2(new_n569), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(new_n554), .Z(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT55), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(KEYINPUT56), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n909), .B1(new_n915), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT56), .B1(new_n913), .B2(G210), .ZN(new_n923));
  INV_X1    g737(.A(new_n918), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(G210), .ZN(new_n926));
  AOI211_X1 g740(.A(new_n926), .B(new_n301), .C1(new_n912), .C2(new_n892), .ZN(new_n927));
  OAI211_X1 g741(.A(KEYINPUT119), .B(new_n918), .C1(new_n927), .C2(KEYINPUT56), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(KEYINPUT121), .B1(new_n921), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n912), .A2(new_n892), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT120), .B1(new_n931), .B2(G902), .ZN(new_n932));
  AOI211_X1 g746(.A(new_n910), .B(new_n301), .C1(new_n912), .C2(new_n892), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n584), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n908), .B1(new_n934), .B2(new_n919), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n935), .A2(new_n936), .A3(new_n925), .A4(new_n928), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n930), .A2(new_n937), .ZN(G51));
  NAND2_X1  g752(.A1(new_n931), .A2(KEYINPUT54), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n896), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n778), .A2(KEYINPUT57), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n778), .A2(KEYINPUT57), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n690), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n911), .A2(new_n914), .ZN(new_n945));
  INV_X1    g759(.A(new_n777), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n908), .B1(new_n944), .B2(new_n947), .ZN(G54));
  NAND3_X1  g762(.A1(new_n945), .A2(KEYINPUT58), .A3(G475), .ZN(new_n949));
  INV_X1    g763(.A(new_n494), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n945), .A2(KEYINPUT58), .A3(G475), .A4(new_n494), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n951), .A2(new_n909), .A3(new_n952), .ZN(G60));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT59), .Z(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n896), .B2(new_n939), .ZN(new_n956));
  INV_X1    g770(.A(new_n612), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n896), .A2(new_n884), .ZN(new_n958));
  OAI211_X1 g772(.A(KEYINPUT122), .B(new_n957), .C1(new_n958), .C2(new_n955), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n955), .B1(new_n896), .B2(new_n884), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n961), .B2(new_n612), .ZN(new_n962));
  AOI221_X4 g776(.A(new_n908), .B1(new_n612), .B2(new_n956), .C1(new_n959), .C2(new_n962), .ZN(G63));
  NAND2_X1  g777(.A1(G217), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT60), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n894), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n908), .B1(new_n966), .B2(new_n632), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n372), .A2(new_n376), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n967), .B1(new_n968), .B2(new_n966), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G66));
  AOI21_X1  g785(.A(new_n277), .B1(new_n547), .B2(G224), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n888), .A2(new_n873), .A3(new_n872), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n972), .B1(new_n974), .B2(new_n277), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n916), .B1(G898), .B2(new_n277), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n975), .B(new_n976), .Z(G69));
  NAND2_X1  g791(.A1(new_n239), .A2(new_n253), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n478), .B1(new_n349), .B2(new_n477), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(new_n980));
  XNOR2_X1  g794(.A(KEYINPUT123), .B(KEYINPUT124), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n829), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n666), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT62), .Z(new_n985));
  NAND4_X1  g799(.A1(new_n663), .A2(new_n682), .A3(new_n764), .A4(new_n869), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n985), .A2(new_n785), .A3(new_n792), .A4(new_n986), .ZN(new_n987));
  OR2_X1    g801(.A1(new_n987), .A2(G953), .ZN(new_n988));
  NAND3_X1  g802(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n982), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n425), .A2(G900), .A3(G953), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT125), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n791), .A2(KEYINPUT110), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n791), .A2(KEYINPUT110), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n785), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n833), .A2(new_n385), .A3(new_n737), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n783), .A2(new_n662), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n748), .A2(new_n751), .A3(new_n983), .A4(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n992), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n998), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n1000), .A2(new_n792), .A3(KEYINPUT125), .A4(new_n785), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n991), .B1(new_n1002), .B2(G953), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n990), .B1(new_n982), .B2(new_n1003), .ZN(G72));
  NAND3_X1  g818(.A1(new_n999), .A2(new_n1001), .A3(new_n973), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT63), .Z(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(KEYINPUT126), .ZN(new_n1009));
  INV_X1    g823(.A(new_n302), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT126), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1005), .A2(new_n1011), .A3(new_n1007), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1009), .A2(new_n1010), .A3(new_n293), .A4(new_n1012), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n1013), .A2(KEYINPUT127), .A3(new_n909), .ZN(new_n1014));
  AOI21_X1  g828(.A(KEYINPUT127), .B1(new_n1013), .B2(new_n909), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1007), .B1(new_n987), .B2(new_n974), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n302), .A3(new_n281), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1007), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n706), .A2(new_n707), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(new_n282), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n880), .B(new_n1020), .C1(new_n883), .C2(new_n844), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  NOR3_X1   g836(.A1(new_n1014), .A2(new_n1015), .A3(new_n1022), .ZN(G57));
endmodule


