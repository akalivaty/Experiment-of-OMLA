//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(KEYINPUT69), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(G567), .B2(new_n456), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(KEYINPUT69), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  INV_X1    g043(.A(G101), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  OAI22_X1  g047(.A1(new_n467), .A2(new_n468), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n465), .A2(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n466), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n473), .A2(new_n476), .ZN(G160));
  INV_X1    g052(.A(new_n467), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(new_n470), .ZN(new_n481));
  NAND2_X1  g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n466), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n479), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND3_X1  g063(.A1(new_n465), .A2(G126), .A3(G2105), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g067(.A1(new_n466), .A2(G138), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n465), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n465), .A2(new_n496), .A3(new_n493), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n495), .B2(new_n497), .ZN(G164));
  INV_X1    g073(.A(G62), .ZN(new_n499));
  OR2_X1    g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(G75), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT71), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(G75), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(G651), .B1(new_n502), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n500), .A2(new_n501), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT70), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n522), .A2(G88), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n515), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND3_X1  g103(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n529));
  INV_X1    g104(.A(new_n512), .ZN(new_n530));
  INV_X1    g105(.A(G51), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n522), .A2(new_n525), .ZN(new_n535));
  INV_X1    g110(.A(G89), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n539));
  OAI211_X1 g114(.A(new_n539), .B(new_n534), .C1(new_n535), .C2(new_n536), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n532), .B1(new_n538), .B2(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n518), .A2(new_n519), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT73), .B(G52), .Z(new_n546));
  AOI22_X1  g121(.A1(new_n545), .A2(G651), .B1(new_n512), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n522), .A2(G90), .A3(new_n525), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT74), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g125(.A(KEYINPUT74), .B1(new_n547), .B2(new_n548), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(G68), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G56), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n543), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n556), .A2(G651), .B1(G43), .B2(new_n512), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n522), .A2(G81), .A3(new_n525), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT75), .ZN(G176));
  XOR2_X1   g138(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n564));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n543), .B2(new_n569), .ZN(new_n570));
  AND2_X1   g145(.A1(G53), .A2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n571), .B1(new_n517), .B2(new_n516), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT9), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n524), .A2(new_n574), .A3(new_n571), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n570), .A2(G651), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n522), .A2(G91), .A3(new_n525), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G299));
  INV_X1    g153(.A(G168), .ZN(G286));
  OR2_X1    g154(.A1(new_n523), .A2(G74), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n512), .B2(G49), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n522), .A2(G87), .A3(new_n525), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n543), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(G48), .B2(new_n512), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n522), .A2(G86), .A3(new_n525), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G305));
  NAND2_X1  g164(.A1(new_n512), .A2(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n535), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(KEYINPUT78), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n594), .B(new_n590), .C1(new_n535), .C2(new_n591), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n597));
  INV_X1    g172(.A(G651), .ZN(new_n598));
  OR3_X1    g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n596), .B2(new_n598), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n593), .A2(new_n595), .A3(new_n601), .ZN(G290));
  NAND3_X1  g177(.A1(new_n522), .A2(G92), .A3(new_n525), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n522), .A2(KEYINPUT10), .A3(G92), .A4(new_n525), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n512), .A2(G54), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n523), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n598), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  MUX2_X1   g187(.A(new_n612), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g188(.A(new_n612), .B(G301), .S(G868), .Z(G321));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G299), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G280));
  XNOR2_X1  g192(.A(G280), .B(KEYINPUT79), .ZN(G297));
  AOI21_X1  g193(.A(new_n610), .B1(new_n605), .B2(new_n606), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n559), .A2(new_n615), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n612), .A2(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n465), .A2(new_n471), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  XOR2_X1   g203(.A(KEYINPUT80), .B(G2100), .Z(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n483), .A2(G123), .ZN(new_n632));
  NOR2_X1   g207(.A1(new_n466), .A2(G111), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(G135), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n632), .B1(new_n633), .B2(new_n634), .C1(new_n635), .C2(new_n467), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n631), .A3(new_n637), .ZN(G156));
  XOR2_X1   g213(.A(KEYINPUT15), .B(G2435), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2430), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT82), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  INV_X1    g231(.A(KEYINPUT18), .ZN(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2100), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2096), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT83), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT84), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n670), .A2(new_n672), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n673), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n675), .ZN(new_n678));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g255(.A1(new_n676), .A2(KEYINPUT20), .A3(new_n675), .ZN(new_n681));
  OAI221_X1 g256(.A(new_n677), .B1(new_n675), .B2(new_n673), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G1991), .B(G1996), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n686), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n687), .A2(new_n690), .A3(new_n688), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(G229));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G35), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G162), .B2(new_n695), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT29), .B(G2090), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n483), .A2(G128), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n466), .A2(G116), .ZN(new_n701));
  OAI21_X1  g276(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n702));
  INV_X1    g277(.A(G140), .ZN(new_n703));
  OAI221_X1 g278(.A(new_n700), .B1(new_n701), .B2(new_n702), .C1(new_n703), .C2(new_n467), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n695), .A2(G26), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G2067), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT92), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT26), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n478), .A2(G141), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n483), .A2(G129), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n471), .A2(G105), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n713), .A2(new_n714), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(new_n695), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n695), .B2(G32), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT27), .B(G1996), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n699), .B(new_n710), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT87), .B(G1348), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G4), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n619), .B2(new_n727), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n724), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n727), .A2(G5), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G171), .B2(new_n727), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G1961), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n727), .A2(G19), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n560), .B2(new_n727), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1341), .Z(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT30), .B(G28), .ZN(new_n737));
  OR2_X1    g312(.A1(KEYINPUT31), .A2(G11), .ZN(new_n738));
  NAND2_X1  g313(.A1(KEYINPUT31), .A2(G11), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n737), .A2(new_n695), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n636), .B2(new_n695), .ZN(new_n741));
  NOR2_X1   g316(.A1(G27), .A2(G29), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G164), .B2(G29), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G2078), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(G34), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G29), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n749), .A2(KEYINPUT91), .B1(G34), .B2(new_n747), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(KEYINPUT91), .B2(new_n749), .ZN(new_n751));
  INV_X1    g326(.A(G160), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n695), .ZN(new_n753));
  INV_X1    g328(.A(G2084), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n753), .A2(new_n754), .B1(G2078), .B2(new_n743), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n736), .A2(new_n746), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n727), .A2(G20), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT23), .ZN(new_n758));
  INV_X1    g333(.A(G299), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n727), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT94), .B(G1956), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n733), .A2(new_n756), .A3(new_n762), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n730), .B(new_n763), .C1(new_n726), .C2(new_n729), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n727), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n727), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1966), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n722), .A2(new_n723), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n754), .B2(new_n753), .ZN(new_n769));
  AND2_X1   g344(.A1(new_n695), .A2(G33), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(new_n466), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT89), .Z(new_n773));
  NAND3_X1  g348(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT25), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G139), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(new_n467), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT88), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n773), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n770), .B1(new_n781), .B2(G29), .ZN(new_n782));
  INV_X1    g357(.A(G2072), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n769), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n767), .B1(new_n786), .B2(KEYINPUT93), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(KEYINPUT93), .B2(new_n786), .ZN(new_n788));
  NOR2_X1   g363(.A1(G6), .A2(G16), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n587), .A2(new_n588), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(G16), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT32), .B(G1981), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT86), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(KEYINPUT86), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n727), .A2(G22), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G166), .B2(new_n727), .ZN(new_n797));
  INV_X1    g372(.A(G1971), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n727), .A2(G23), .ZN(new_n800));
  INV_X1    g375(.A(G288), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n727), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT33), .B(G1976), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n794), .A2(new_n795), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n483), .A2(G119), .ZN(new_n808));
  OR2_X1    g383(.A1(G95), .A2(G2105), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n809), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n810));
  INV_X1    g385(.A(G131), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n808), .B(new_n810), .C1(new_n811), .C2(new_n467), .ZN(new_n812));
  MUX2_X1   g387(.A(G25), .B(new_n812), .S(G29), .Z(new_n813));
  XOR2_X1   g388(.A(KEYINPUT35), .B(G1991), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n727), .A2(G24), .ZN(new_n816));
  INV_X1    g391(.A(G290), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n727), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT85), .B(G1986), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n818), .B(new_n819), .Z(new_n820));
  NAND4_X1  g395(.A1(new_n806), .A2(new_n807), .A3(new_n815), .A4(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT36), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT36), .ZN(new_n823));
  AOI211_X1 g398(.A(new_n764), .B(new_n788), .C1(new_n822), .C2(new_n823), .ZN(G311));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n788), .A2(new_n764), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(G150));
  NAND3_X1  g402(.A1(new_n522), .A2(G93), .A3(new_n525), .ZN(new_n828));
  OAI21_X1  g403(.A(G67), .B1(new_n518), .B2(new_n519), .ZN(new_n829));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n831), .A2(G651), .B1(G55), .B2(new_n512), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT96), .B(G860), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT37), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n619), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n559), .A2(new_n833), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n557), .A2(new_n558), .A3(new_n828), .A4(new_n832), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n840), .B(new_n843), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT39), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT97), .Z(new_n846));
  OAI21_X1  g421(.A(new_n835), .B1(new_n844), .B2(KEYINPUT39), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n837), .B1(new_n846), .B2(new_n847), .ZN(G145));
  INV_X1    g423(.A(KEYINPUT104), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT102), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n812), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n627), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n812), .B(KEYINPUT102), .ZN(new_n853));
  INV_X1    g428(.A(new_n627), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n856));
  INV_X1    g431(.A(G142), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n467), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n856), .B1(new_n467), .B2(new_n857), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n863));
  INV_X1    g438(.A(new_n483), .ZN(new_n864));
  INV_X1    g439(.A(G130), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n852), .A2(new_n855), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n867), .B1(new_n852), .B2(new_n855), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n720), .A2(G164), .ZN(new_n872));
  INV_X1    g447(.A(new_n497), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n496), .B1(new_n465), .B2(new_n493), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n719), .B1(new_n875), .B2(new_n492), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n704), .B(KEYINPUT99), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n781), .A2(KEYINPUT100), .ZN(new_n880));
  INV_X1    g455(.A(new_n878), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n881), .A2(new_n876), .A3(new_n872), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT100), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n773), .A2(new_n780), .A3(new_n884), .ZN(new_n885));
  AOI22_X1  g460(.A1(new_n879), .A2(new_n882), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n871), .B(KEYINPUT103), .C1(new_n883), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n880), .A2(new_n885), .ZN(new_n888));
  INV_X1    g463(.A(new_n882), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n881), .B1(new_n872), .B2(new_n876), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n870), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n892), .A2(KEYINPUT103), .A3(new_n868), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n869), .B2(new_n870), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n891), .A2(new_n893), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n887), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n487), .B(G160), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT98), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n636), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n849), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n887), .A2(new_n901), .A3(new_n897), .A4(KEYINPUT104), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(KEYINPUT105), .B(G37), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n898), .B2(new_n902), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g485(.A1(G305), .A2(new_n526), .A3(new_n515), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n522), .A2(G88), .A3(new_n525), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n588), .B(new_n587), .C1(new_n912), .C2(new_n514), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n911), .A2(new_n913), .A3(G288), .ZN(new_n914));
  AOI21_X1  g489(.A(G288), .B1(new_n911), .B2(new_n913), .ZN(new_n915));
  OAI21_X1  g490(.A(G290), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n801), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n911), .A2(new_n913), .A3(G288), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n817), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n921), .A2(KEYINPUT109), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n923), .B1(new_n924), .B2(new_n922), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT42), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n610), .B1(new_n576), .B2(new_n577), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n607), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT41), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n619), .A2(G299), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT106), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n928), .B1(G299), .B2(new_n619), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n612), .A2(new_n759), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n607), .B2(new_n927), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n931), .A2(new_n934), .A3(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n623), .B(new_n843), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n932), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT107), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n943), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n924), .A2(new_n947), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n926), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n946), .B1(new_n926), .B2(new_n948), .ZN(new_n950));
  OAI21_X1  g525(.A(G868), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(G868), .B2(new_n834), .ZN(G295));
  OAI21_X1  g527(.A(new_n951), .B1(G868), .B2(new_n834), .ZN(G331));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  INV_X1    g530(.A(new_n551), .ZN(new_n956));
  AND4_X1   g531(.A1(new_n558), .A2(new_n557), .A3(new_n828), .A4(new_n832), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n558), .A2(new_n557), .B1(new_n828), .B2(new_n832), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n549), .B(new_n956), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n841), .B(new_n842), .C1(new_n550), .C2(new_n551), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n959), .A2(G168), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G168), .B1(new_n959), .B2(new_n960), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n939), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n960), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(G286), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n959), .A2(G168), .A3(new_n960), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(new_n932), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n916), .A2(new_n920), .A3(KEYINPUT108), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n963), .A2(new_n923), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G37), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n935), .A2(new_n937), .ZN(new_n972));
  AOI22_X1  g547(.A1(new_n972), .A2(KEYINPUT106), .B1(new_n932), .B2(new_n933), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n973), .A2(new_n938), .B1(new_n965), .B2(new_n966), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n961), .A2(new_n962), .A3(new_n944), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT108), .B1(new_n916), .B2(new_n920), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n916), .A2(new_n920), .A3(KEYINPUT108), .ZN(new_n977));
  OAI22_X1  g552(.A1(new_n974), .A2(new_n975), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n955), .B1(new_n971), .B2(new_n978), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n965), .A2(new_n966), .B1(new_n972), .B2(new_n934), .ZN(new_n980));
  OAI22_X1  g555(.A1(new_n980), .A2(new_n975), .B1(new_n977), .B2(new_n976), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n969), .A2(new_n981), .A3(new_n906), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n954), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(KEYINPUT110), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n969), .A2(new_n981), .A3(new_n986), .A4(new_n906), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(KEYINPUT43), .A3(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n978), .A2(new_n969), .A3(new_n955), .A4(new_n970), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n989), .A2(KEYINPUT44), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n988), .A2(KEYINPUT111), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT111), .B1(new_n988), .B2(new_n990), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n984), .B1(new_n991), .B2(new_n992), .ZN(G397));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(G164), .B2(G1384), .ZN(new_n995));
  INV_X1    g570(.A(new_n473), .ZN(new_n996));
  INV_X1    g571(.A(new_n476), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT112), .B(G40), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n995), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OR3_X1    g577(.A1(new_n1002), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT46), .B1(new_n1002), .B2(G1996), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n704), .B(G2067), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1005), .A2(new_n719), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1003), .A2(new_n1004), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1002), .A2(G1996), .A3(new_n719), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT113), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n719), .A2(G1996), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1012), .A2(new_n1005), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1011), .B1(new_n1001), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n812), .B(new_n814), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n1015), .A2(KEYINPUT114), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(KEYINPUT114), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1016), .A2(new_n1001), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  OR2_X1    g594(.A1(G290), .A2(G1986), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1020), .A2(new_n1002), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(KEYINPUT48), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1009), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n814), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n812), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1014), .A2(new_n1025), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n704), .A2(G2067), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1002), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1023), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G8), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n495), .A2(new_n497), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n489), .A2(new_n491), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1384), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT45), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n473), .A2(new_n476), .A3(new_n998), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n995), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n798), .ZN(new_n1037));
  INV_X1    g612(.A(G1384), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n875), .B2(new_n492), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1000), .B1(new_n1039), .B2(KEYINPUT50), .ZN(new_n1040));
  INV_X1    g615(.A(G2090), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1033), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1030), .B1(new_n1037), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1047), .B(new_n1030), .C1(new_n515), .C2(new_n526), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1045), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1981), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n586), .A2(G651), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1052), .B1(new_n1053), .B2(KEYINPUT116), .ZN(new_n1054));
  NOR2_X1   g629(.A1(G305), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G305), .A2(new_n1054), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(KEYINPUT49), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT49), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1057), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n1055), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1030), .B1(new_n1035), .B2(new_n1033), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1058), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1035), .A2(new_n1033), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G8), .ZN(new_n1066));
  INV_X1    g641(.A(G1976), .ZN(new_n1067));
  NOR2_X1   g642(.A1(G288), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT52), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(G288), .B2(new_n1067), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1062), .B(new_n1070), .C1(new_n1067), .C2(G288), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1064), .A2(new_n1072), .ZN(new_n1073));
  AND3_X1   g648(.A1(new_n1033), .A2(KEYINPUT115), .A3(new_n1042), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT115), .B1(new_n1033), .B2(new_n1042), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1040), .B(new_n1041), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1037), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(G8), .A3(new_n1050), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1040), .B(new_n754), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1079));
  INV_X1    g654(.A(G1966), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1036), .A2(new_n1080), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1030), .B(G286), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1051), .A2(new_n1073), .A3(new_n1078), .A4(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT63), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT117), .B1(new_n1064), .B2(new_n1072), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1072), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(new_n1088), .A3(new_n1063), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  AOI211_X1 g665(.A(new_n1030), .B(new_n1049), .C1(new_n1076), .C2(new_n1037), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1092), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1077), .A2(G8), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n1049), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1090), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1085), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1063), .A2(new_n1067), .A3(new_n801), .ZN(new_n1099));
  NOR2_X1   g674(.A1(G305), .A2(G1981), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1100), .B(KEYINPUT118), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1066), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1102), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1087), .B(new_n1063), .C1(new_n1045), .C2(new_n1050), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1040), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1105));
  INV_X1    g680(.A(G1961), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1108), .A2(G2078), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n995), .A2(new_n1034), .A3(new_n1035), .A4(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n995), .A2(new_n1034), .A3(new_n745), .A4(new_n1035), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n1108), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1107), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(G171), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1104), .A2(new_n1114), .A3(new_n1091), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1079), .A2(new_n1081), .A3(G168), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1116), .A2(new_n1117), .A3(G8), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1092), .A2(G286), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1119), .A2(G8), .A3(new_n1116), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1118), .B1(new_n1120), .B2(KEYINPUT51), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1115), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g698(.A(KEYINPUT62), .B(new_n1118), .C1(KEYINPUT51), .C2(new_n1120), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1098), .B(new_n1103), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1107), .A2(KEYINPUT123), .ZN(new_n1126));
  AND3_X1   g701(.A1(G160), .A2(G40), .A3(new_n1109), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(new_n995), .A3(new_n1034), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1127), .A2(new_n995), .A3(new_n1034), .A4(KEYINPUT124), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1130), .A2(new_n1131), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1105), .A2(new_n1133), .A3(new_n1106), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1126), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1114), .B1(new_n1135), .B2(G171), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1104), .A2(new_n1091), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1120), .A2(KEYINPUT51), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1118), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1138), .A2(new_n1139), .A3(new_n1142), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT56), .B(G2072), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1036), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(G1956), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n1150));
  OAI21_X1  g725(.A(G299), .B1(KEYINPUT119), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(KEYINPUT119), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1151), .B(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1149), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1144), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1105), .A2(new_n725), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1035), .A2(new_n1033), .A3(new_n709), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n1160), .B(KEYINPUT120), .Z(new_n1161));
  NOR4_X1   g736(.A1(new_n1159), .A2(new_n1161), .A3(KEYINPUT60), .A4(new_n612), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT58), .B(G1341), .Z(new_n1163));
  NAND2_X1  g738(.A1(new_n1065), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(new_n1036), .B2(G1996), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1165), .A2(new_n1166), .A3(new_n560), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1166), .B1(new_n1165), .B2(new_n560), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1158), .A2(new_n1162), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1156), .A2(new_n1157), .A3(KEYINPUT61), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1156), .A2(new_n1157), .A3(KEYINPUT122), .A4(KEYINPUT61), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1176), .A2(new_n612), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1159), .A2(new_n1161), .A3(new_n619), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT60), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1170), .A2(new_n1175), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1157), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1181), .B1(new_n1177), .B2(new_n1156), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1143), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1135), .A2(KEYINPUT125), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1126), .A2(new_n1132), .A3(new_n1185), .A4(new_n1134), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1184), .A2(G171), .A3(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1113), .A2(G171), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1188), .A2(new_n1137), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1187), .A2(KEYINPUT126), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT126), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1125), .B1(new_n1183), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(G290), .A2(G1986), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1002), .B1(new_n1020), .B2(new_n1194), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1019), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1029), .B1(new_n1193), .B2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g772(.A1(new_n463), .A2(G227), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n655), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1200), .B1(new_n692), .B2(new_n693), .ZN(new_n1201));
  OAI211_X1 g775(.A(new_n1201), .B(new_n909), .C1(new_n979), .C2(new_n983), .ZN(G225));
  INV_X1    g776(.A(G225), .ZN(G308));
endmodule


