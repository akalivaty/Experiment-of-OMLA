

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U547 ( .A1(n754), .A2(n753), .ZN(n692) );
  INV_X1 U548 ( .A(n692), .ZN(n708) );
  AND2_X2 U549 ( .A1(n534), .A2(G2104), .ZN(n867) );
  NAND2_X1 U550 ( .A1(n692), .A2(G1996), .ZN(n666) );
  XNOR2_X1 U551 ( .A(KEYINPUT26), .B(KEYINPUT90), .ZN(n509) );
  XNOR2_X1 U552 ( .A(n666), .B(n509), .ZN(n668) );
  XNOR2_X1 U553 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X1 U554 ( .A1(n671), .A2(n927), .ZN(n673) );
  AND2_X1 U555 ( .A1(n721), .A2(n720), .ZN(n724) );
  OR2_X1 U556 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U557 ( .A(KEYINPUT80), .B(n665), .Z(n753) );
  OR2_X1 U558 ( .A1(n750), .A2(n749), .ZN(n751) );
  NOR2_X1 U559 ( .A1(G651), .A2(n608), .ZN(n626) );
  NOR2_X1 U560 ( .A1(G651), .A2(G543), .ZN(n618) );
  NAND2_X1 U561 ( .A1(n618), .A2(G89), .ZN(n510) );
  XNOR2_X1 U562 ( .A(KEYINPUT4), .B(n510), .ZN(n513) );
  XOR2_X1 U563 ( .A(G543), .B(KEYINPUT0), .Z(n608) );
  INV_X1 U564 ( .A(G651), .ZN(n515) );
  NOR2_X1 U565 ( .A1(n608), .A2(n515), .ZN(n622) );
  NAND2_X1 U566 ( .A1(n622), .A2(G76), .ZN(n511) );
  XOR2_X1 U567 ( .A(KEYINPUT73), .B(n511), .Z(n512) );
  NAND2_X1 U568 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U569 ( .A(n514), .B(KEYINPUT5), .ZN(n521) );
  NOR2_X1 U570 ( .A1(G543), .A2(n515), .ZN(n516) );
  XOR2_X1 U571 ( .A(KEYINPUT1), .B(n516), .Z(n619) );
  NAND2_X1 U572 ( .A1(G63), .A2(n619), .ZN(n518) );
  NAND2_X1 U573 ( .A1(G51), .A2(n626), .ZN(n517) );
  NAND2_X1 U574 ( .A1(n518), .A2(n517), .ZN(n519) );
  XOR2_X1 U575 ( .A(KEYINPUT6), .B(n519), .Z(n520) );
  NAND2_X1 U576 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U577 ( .A(n522), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U578 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U579 ( .A1(G85), .A2(n618), .ZN(n524) );
  NAND2_X1 U580 ( .A1(G72), .A2(n622), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n524), .A2(n523), .ZN(n528) );
  NAND2_X1 U582 ( .A1(G60), .A2(n619), .ZN(n526) );
  NAND2_X1 U583 ( .A1(G47), .A2(n626), .ZN(n525) );
  NAND2_X1 U584 ( .A1(n526), .A2(n525), .ZN(n527) );
  OR2_X1 U585 ( .A1(n528), .A2(n527), .ZN(G290) );
  AND2_X1 U586 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U587 ( .A(G57), .ZN(G237) );
  INV_X1 U588 ( .A(G132), .ZN(G219) );
  INV_X1 U589 ( .A(G82), .ZN(G220) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n863) );
  NAND2_X1 U591 ( .A1(G113), .A2(n863), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n529), .B(KEYINPUT64), .ZN(n532) );
  INV_X1 U593 ( .A(G2105), .ZN(n534) );
  NAND2_X1 U594 ( .A1(G101), .A2(n867), .ZN(n530) );
  XOR2_X1 U595 ( .A(KEYINPUT23), .B(n530), .Z(n531) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n664) );
  NOR2_X1 U597 ( .A1(G2105), .A2(G2104), .ZN(n533) );
  XOR2_X1 U598 ( .A(KEYINPUT17), .B(n533), .Z(n852) );
  NAND2_X1 U599 ( .A1(G137), .A2(n852), .ZN(n536) );
  NOR2_X2 U600 ( .A1(G2104), .A2(n534), .ZN(n864) );
  NAND2_X1 U601 ( .A1(G125), .A2(n864), .ZN(n535) );
  NAND2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n662) );
  NOR2_X1 U603 ( .A1(n664), .A2(n662), .ZN(G160) );
  NAND2_X1 U604 ( .A1(G7), .A2(G661), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n537), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U606 ( .A(G223), .ZN(n809) );
  NAND2_X1 U607 ( .A1(n809), .A2(G567), .ZN(n538) );
  XOR2_X1 U608 ( .A(KEYINPUT11), .B(n538), .Z(G234) );
  XNOR2_X1 U609 ( .A(KEYINPUT13), .B(KEYINPUT71), .ZN(n544) );
  NAND2_X1 U610 ( .A1(G81), .A2(n618), .ZN(n539) );
  XNOR2_X1 U611 ( .A(n539), .B(KEYINPUT12), .ZN(n540) );
  XNOR2_X1 U612 ( .A(n540), .B(KEYINPUT70), .ZN(n542) );
  NAND2_X1 U613 ( .A1(G68), .A2(n622), .ZN(n541) );
  NAND2_X1 U614 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U615 ( .A(n544), .B(n543), .ZN(n547) );
  NAND2_X1 U616 ( .A1(n619), .A2(G56), .ZN(n545) );
  XOR2_X1 U617 ( .A(KEYINPUT14), .B(n545), .Z(n546) );
  NOR2_X1 U618 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U619 ( .A(n548), .B(KEYINPUT72), .ZN(n550) );
  NAND2_X1 U620 ( .A1(G43), .A2(n626), .ZN(n549) );
  NAND2_X1 U621 ( .A1(n550), .A2(n549), .ZN(n927) );
  INV_X1 U622 ( .A(G860), .ZN(n596) );
  OR2_X1 U623 ( .A1(n927), .A2(n596), .ZN(G153) );
  NAND2_X1 U624 ( .A1(n619), .A2(G64), .ZN(n551) );
  XOR2_X1 U625 ( .A(KEYINPUT65), .B(n551), .Z(n553) );
  NAND2_X1 U626 ( .A1(n626), .A2(G52), .ZN(n552) );
  NAND2_X1 U627 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U628 ( .A(KEYINPUT66), .B(n554), .ZN(n560) );
  NAND2_X1 U629 ( .A1(n618), .A2(G90), .ZN(n555) );
  XOR2_X1 U630 ( .A(KEYINPUT67), .B(n555), .Z(n557) );
  NAND2_X1 U631 ( .A1(n622), .A2(G77), .ZN(n556) );
  NAND2_X1 U632 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U633 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U634 ( .A1(n560), .A2(n559), .ZN(G171) );
  INV_X1 U635 ( .A(G171), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G868), .A2(G301), .ZN(n569) );
  NAND2_X1 U637 ( .A1(G92), .A2(n618), .ZN(n562) );
  NAND2_X1 U638 ( .A1(G79), .A2(n622), .ZN(n561) );
  NAND2_X1 U639 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U640 ( .A1(G66), .A2(n619), .ZN(n564) );
  NAND2_X1 U641 ( .A1(G54), .A2(n626), .ZN(n563) );
  NAND2_X1 U642 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U643 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U644 ( .A(KEYINPUT15), .B(n567), .Z(n924) );
  OR2_X1 U645 ( .A1(n924), .A2(G868), .ZN(n568) );
  NAND2_X1 U646 ( .A1(n569), .A2(n568), .ZN(G284) );
  NAND2_X1 U647 ( .A1(G91), .A2(n618), .ZN(n571) );
  NAND2_X1 U648 ( .A1(G78), .A2(n622), .ZN(n570) );
  NAND2_X1 U649 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U650 ( .A(KEYINPUT68), .B(n572), .ZN(n575) );
  NAND2_X1 U651 ( .A1(G65), .A2(n619), .ZN(n573) );
  XNOR2_X1 U652 ( .A(KEYINPUT69), .B(n573), .ZN(n574) );
  NOR2_X1 U653 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U654 ( .A1(n626), .A2(G53), .ZN(n576) );
  NAND2_X1 U655 ( .A1(n577), .A2(n576), .ZN(G299) );
  NOR2_X1 U656 ( .A1(G868), .A2(G299), .ZN(n579) );
  INV_X1 U657 ( .A(G868), .ZN(n638) );
  NOR2_X1 U658 ( .A1(G286), .A2(n638), .ZN(n578) );
  NOR2_X1 U659 ( .A1(n579), .A2(n578), .ZN(G297) );
  NAND2_X1 U660 ( .A1(n596), .A2(G559), .ZN(n580) );
  NAND2_X1 U661 ( .A1(n580), .A2(n924), .ZN(n581) );
  XNOR2_X1 U662 ( .A(n581), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U663 ( .A1(G868), .A2(n927), .ZN(n584) );
  NAND2_X1 U664 ( .A1(G868), .A2(n924), .ZN(n582) );
  NOR2_X1 U665 ( .A1(G559), .A2(n582), .ZN(n583) );
  NOR2_X1 U666 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U667 ( .A(KEYINPUT74), .B(n585), .ZN(G282) );
  NAND2_X1 U668 ( .A1(G123), .A2(n864), .ZN(n586) );
  XNOR2_X1 U669 ( .A(n586), .B(KEYINPUT18), .ZN(n588) );
  NAND2_X1 U670 ( .A1(n863), .A2(G111), .ZN(n587) );
  NAND2_X1 U671 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U672 ( .A1(G99), .A2(n867), .ZN(n590) );
  BUF_X1 U673 ( .A(n852), .Z(n869) );
  NAND2_X1 U674 ( .A1(G135), .A2(n869), .ZN(n589) );
  NAND2_X1 U675 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U676 ( .A1(n592), .A2(n591), .ZN(n987) );
  XNOR2_X1 U677 ( .A(n987), .B(G2096), .ZN(n594) );
  INV_X1 U678 ( .A(G2100), .ZN(n593) );
  NAND2_X1 U679 ( .A1(n594), .A2(n593), .ZN(G156) );
  NAND2_X1 U680 ( .A1(G559), .A2(n924), .ZN(n595) );
  XOR2_X1 U681 ( .A(n927), .B(n595), .Z(n636) );
  NAND2_X1 U682 ( .A1(n596), .A2(n636), .ZN(n604) );
  NAND2_X1 U683 ( .A1(G93), .A2(n618), .ZN(n598) );
  NAND2_X1 U684 ( .A1(G80), .A2(n622), .ZN(n597) );
  NAND2_X1 U685 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U686 ( .A1(G67), .A2(n619), .ZN(n599) );
  XNOR2_X1 U687 ( .A(KEYINPUT75), .B(n599), .ZN(n600) );
  NOR2_X1 U688 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U689 ( .A1(n626), .A2(G55), .ZN(n602) );
  NAND2_X1 U690 ( .A1(n603), .A2(n602), .ZN(n639) );
  XNOR2_X1 U691 ( .A(n604), .B(n639), .ZN(G145) );
  NAND2_X1 U692 ( .A1(G49), .A2(n626), .ZN(n606) );
  NAND2_X1 U693 ( .A1(G74), .A2(G651), .ZN(n605) );
  NAND2_X1 U694 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U695 ( .A1(n619), .A2(n607), .ZN(n610) );
  NAND2_X1 U696 ( .A1(n608), .A2(G87), .ZN(n609) );
  NAND2_X1 U697 ( .A1(n610), .A2(n609), .ZN(G288) );
  NAND2_X1 U698 ( .A1(G88), .A2(n618), .ZN(n612) );
  NAND2_X1 U699 ( .A1(G75), .A2(n622), .ZN(n611) );
  NAND2_X1 U700 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U701 ( .A1(n619), .A2(G62), .ZN(n613) );
  XOR2_X1 U702 ( .A(KEYINPUT76), .B(n613), .Z(n614) );
  NOR2_X1 U703 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U704 ( .A1(n626), .A2(G50), .ZN(n616) );
  NAND2_X1 U705 ( .A1(n617), .A2(n616), .ZN(G303) );
  INV_X1 U706 ( .A(G303), .ZN(G166) );
  NAND2_X1 U707 ( .A1(G86), .A2(n618), .ZN(n621) );
  NAND2_X1 U708 ( .A1(G61), .A2(n619), .ZN(n620) );
  NAND2_X1 U709 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U710 ( .A1(n622), .A2(G73), .ZN(n623) );
  XOR2_X1 U711 ( .A(KEYINPUT2), .B(n623), .Z(n624) );
  NOR2_X1 U712 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U713 ( .A1(n626), .A2(G48), .ZN(n627) );
  NAND2_X1 U714 ( .A1(n628), .A2(n627), .ZN(G305) );
  XNOR2_X1 U715 ( .A(KEYINPUT19), .B(KEYINPUT78), .ZN(n630) );
  XNOR2_X1 U716 ( .A(G288), .B(KEYINPUT77), .ZN(n629) );
  XNOR2_X1 U717 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U718 ( .A(G290), .B(n631), .ZN(n633) );
  INV_X1 U719 ( .A(G299), .ZN(n932) );
  XNOR2_X1 U720 ( .A(n932), .B(G166), .ZN(n632) );
  XNOR2_X1 U721 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U722 ( .A(n634), .B(G305), .ZN(n635) );
  XNOR2_X1 U723 ( .A(n635), .B(n639), .ZN(n883) );
  XOR2_X1 U724 ( .A(n883), .B(n636), .Z(n637) );
  NOR2_X1 U725 ( .A1(n638), .A2(n637), .ZN(n641) );
  NOR2_X1 U726 ( .A1(G868), .A2(n639), .ZN(n640) );
  NOR2_X1 U727 ( .A1(n641), .A2(n640), .ZN(G295) );
  NAND2_X1 U728 ( .A1(G2078), .A2(G2084), .ZN(n642) );
  XOR2_X1 U729 ( .A(KEYINPUT20), .B(n642), .Z(n643) );
  NAND2_X1 U730 ( .A1(G2090), .A2(n643), .ZN(n644) );
  XNOR2_X1 U731 ( .A(KEYINPUT21), .B(n644), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n645), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U733 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U734 ( .A1(G220), .A2(G219), .ZN(n646) );
  XOR2_X1 U735 ( .A(KEYINPUT22), .B(n646), .Z(n647) );
  NOR2_X1 U736 ( .A1(G218), .A2(n647), .ZN(n648) );
  NAND2_X1 U737 ( .A1(G96), .A2(n648), .ZN(n815) );
  NAND2_X1 U738 ( .A1(G2106), .A2(n815), .ZN(n652) );
  NAND2_X1 U739 ( .A1(G69), .A2(G120), .ZN(n649) );
  NOR2_X1 U740 ( .A1(G237), .A2(n649), .ZN(n650) );
  NAND2_X1 U741 ( .A1(G108), .A2(n650), .ZN(n816) );
  NAND2_X1 U742 ( .A1(G567), .A2(n816), .ZN(n651) );
  NAND2_X1 U743 ( .A1(n652), .A2(n651), .ZN(n817) );
  NAND2_X1 U744 ( .A1(G483), .A2(G661), .ZN(n653) );
  NOR2_X1 U745 ( .A1(n817), .A2(n653), .ZN(n812) );
  NAND2_X1 U746 ( .A1(n812), .A2(G36), .ZN(G176) );
  NAND2_X1 U747 ( .A1(n864), .A2(G126), .ZN(n656) );
  NAND2_X1 U748 ( .A1(G102), .A2(n867), .ZN(n654) );
  XOR2_X1 U749 ( .A(KEYINPUT79), .B(n654), .Z(n655) );
  NAND2_X1 U750 ( .A1(n656), .A2(n655), .ZN(n660) );
  NAND2_X1 U751 ( .A1(G114), .A2(n863), .ZN(n658) );
  NAND2_X1 U752 ( .A1(G138), .A2(n852), .ZN(n657) );
  NAND2_X1 U753 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U754 ( .A1(n660), .A2(n659), .ZN(G164) );
  XOR2_X1 U755 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n718) );
  NOR2_X1 U756 ( .A1(G164), .A2(G1384), .ZN(n754) );
  INV_X1 U757 ( .A(G40), .ZN(n661) );
  OR2_X1 U758 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U759 ( .A1(n708), .A2(G1341), .ZN(n667) );
  NAND2_X1 U760 ( .A1(n668), .A2(n667), .ZN(n670) );
  INV_X1 U761 ( .A(KEYINPUT91), .ZN(n669) );
  NOR2_X1 U762 ( .A1(n673), .A2(n924), .ZN(n672) );
  XNOR2_X1 U763 ( .A(n672), .B(KEYINPUT93), .ZN(n680) );
  NAND2_X1 U764 ( .A1(n673), .A2(n924), .ZN(n678) );
  NAND2_X1 U765 ( .A1(G1348), .A2(n708), .ZN(n675) );
  NAND2_X1 U766 ( .A1(n692), .A2(G2067), .ZN(n674) );
  NAND2_X1 U767 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U768 ( .A(KEYINPUT92), .B(n676), .ZN(n677) );
  NAND2_X1 U769 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U770 ( .A1(n680), .A2(n679), .ZN(n686) );
  NAND2_X1 U771 ( .A1(G2072), .A2(n692), .ZN(n681) );
  XNOR2_X1 U772 ( .A(n681), .B(KEYINPUT88), .ZN(n682) );
  XNOR2_X1 U773 ( .A(n682), .B(KEYINPUT27), .ZN(n684) );
  XNOR2_X1 U774 ( .A(G1956), .B(KEYINPUT89), .ZN(n961) );
  NOR2_X1 U775 ( .A1(n961), .A2(n692), .ZN(n683) );
  NOR2_X1 U776 ( .A1(n684), .A2(n683), .ZN(n687) );
  NAND2_X1 U777 ( .A1(n932), .A2(n687), .ZN(n685) );
  NAND2_X1 U778 ( .A1(n686), .A2(n685), .ZN(n690) );
  NOR2_X1 U779 ( .A1(n932), .A2(n687), .ZN(n688) );
  XOR2_X1 U780 ( .A(n688), .B(KEYINPUT28), .Z(n689) );
  NAND2_X1 U781 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U782 ( .A(n691), .B(KEYINPUT29), .ZN(n696) );
  NAND2_X1 U783 ( .A1(G1961), .A2(n708), .ZN(n694) );
  XOR2_X1 U784 ( .A(G2078), .B(KEYINPUT25), .Z(n906) );
  NAND2_X1 U785 ( .A1(n692), .A2(n906), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n694), .A2(n693), .ZN(n700) );
  NOR2_X1 U787 ( .A1(G301), .A2(n700), .ZN(n695) );
  NOR2_X1 U788 ( .A1(n696), .A2(n695), .ZN(n706) );
  NAND2_X1 U789 ( .A1(G8), .A2(n708), .ZN(n741) );
  NOR2_X1 U790 ( .A1(G1966), .A2(n741), .ZN(n719) );
  NOR2_X1 U791 ( .A1(G2084), .A2(n708), .ZN(n722) );
  NOR2_X1 U792 ( .A1(n719), .A2(n722), .ZN(n697) );
  NAND2_X1 U793 ( .A1(G8), .A2(n697), .ZN(n698) );
  XNOR2_X1 U794 ( .A(KEYINPUT30), .B(n698), .ZN(n699) );
  NOR2_X1 U795 ( .A1(G168), .A2(n699), .ZN(n703) );
  NAND2_X1 U796 ( .A1(G301), .A2(n700), .ZN(n701) );
  XOR2_X1 U797 ( .A(KEYINPUT94), .B(n701), .Z(n702) );
  NOR2_X1 U798 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U799 ( .A(n704), .B(KEYINPUT31), .ZN(n705) );
  NOR2_X1 U800 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U801 ( .A(n707), .B(KEYINPUT95), .ZN(n721) );
  NAND2_X1 U802 ( .A1(n721), .A2(G286), .ZN(n715) );
  NOR2_X1 U803 ( .A1(G2090), .A2(n708), .ZN(n709) );
  XNOR2_X1 U804 ( .A(KEYINPUT97), .B(n709), .ZN(n712) );
  NOR2_X1 U805 ( .A1(G1971), .A2(n741), .ZN(n710) );
  NOR2_X1 U806 ( .A1(G166), .A2(n710), .ZN(n711) );
  NAND2_X1 U807 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U808 ( .A(n713), .B(KEYINPUT98), .ZN(n714) );
  NAND2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n716), .A2(G8), .ZN(n717) );
  XNOR2_X1 U811 ( .A(n718), .B(n717), .ZN(n727) );
  INV_X1 U812 ( .A(n719), .ZN(n720) );
  NAND2_X1 U813 ( .A1(G8), .A2(n722), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U815 ( .A(KEYINPUT96), .B(n725), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n737) );
  NOR2_X1 U817 ( .A1(G2090), .A2(G303), .ZN(n728) );
  NAND2_X1 U818 ( .A1(G8), .A2(n728), .ZN(n729) );
  NAND2_X1 U819 ( .A1(n737), .A2(n729), .ZN(n730) );
  XNOR2_X1 U820 ( .A(n730), .B(KEYINPUT100), .ZN(n731) );
  NAND2_X1 U821 ( .A1(n731), .A2(n741), .ZN(n735) );
  NOR2_X1 U822 ( .A1(G1981), .A2(G305), .ZN(n732) );
  XOR2_X1 U823 ( .A(n732), .B(KEYINPUT24), .Z(n733) );
  OR2_X1 U824 ( .A1(n741), .A2(n733), .ZN(n734) );
  NAND2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n752) );
  NOR2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n739) );
  NOR2_X1 U827 ( .A1(G1971), .A2(G303), .ZN(n736) );
  NOR2_X1 U828 ( .A1(n739), .A2(n736), .ZN(n936) );
  AND2_X1 U829 ( .A1(n936), .A2(n737), .ZN(n746) );
  NAND2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n935) );
  INV_X1 U831 ( .A(n741), .ZN(n738) );
  NAND2_X1 U832 ( .A1(n935), .A2(n738), .ZN(n744) );
  XOR2_X1 U833 ( .A(G1981), .B(G305), .Z(n943) );
  INV_X1 U834 ( .A(n943), .ZN(n743) );
  NAND2_X1 U835 ( .A1(n739), .A2(KEYINPUT33), .ZN(n740) );
  NOR2_X1 U836 ( .A1(n741), .A2(n740), .ZN(n742) );
  OR2_X1 U837 ( .A1(n743), .A2(n742), .ZN(n747) );
  OR2_X1 U838 ( .A1(n744), .A2(n747), .ZN(n745) );
  NOR2_X1 U839 ( .A1(n746), .A2(n745), .ZN(n750) );
  INV_X1 U840 ( .A(n747), .ZN(n748) );
  AND2_X1 U841 ( .A1(n748), .A2(KEYINPUT33), .ZN(n749) );
  NOR2_X1 U842 ( .A1(n752), .A2(n751), .ZN(n768) );
  INV_X1 U843 ( .A(n753), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n804) );
  XNOR2_X1 U845 ( .A(G1986), .B(G290), .ZN(n926) );
  NAND2_X1 U846 ( .A1(n804), .A2(n926), .ZN(n766) );
  NAND2_X1 U847 ( .A1(G104), .A2(n867), .ZN(n757) );
  NAND2_X1 U848 ( .A1(G140), .A2(n869), .ZN(n756) );
  NAND2_X1 U849 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U850 ( .A(KEYINPUT34), .B(n758), .ZN(n764) );
  NAND2_X1 U851 ( .A1(n863), .A2(G116), .ZN(n759) );
  XOR2_X1 U852 ( .A(KEYINPUT81), .B(n759), .Z(n761) );
  NAND2_X1 U853 ( .A1(n864), .A2(G128), .ZN(n760) );
  NAND2_X1 U854 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U855 ( .A(KEYINPUT35), .B(n762), .Z(n763) );
  NOR2_X1 U856 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U857 ( .A(KEYINPUT36), .B(n765), .ZN(n878) );
  XNOR2_X1 U858 ( .A(G2067), .B(KEYINPUT37), .ZN(n801) );
  NOR2_X1 U859 ( .A1(n878), .A2(n801), .ZN(n985) );
  NAND2_X1 U860 ( .A1(n804), .A2(n985), .ZN(n798) );
  NAND2_X1 U861 ( .A1(n766), .A2(n798), .ZN(n767) );
  NOR2_X1 U862 ( .A1(n768), .A2(n767), .ZN(n790) );
  NAND2_X1 U863 ( .A1(G119), .A2(n864), .ZN(n770) );
  NAND2_X1 U864 ( .A1(G131), .A2(n869), .ZN(n769) );
  NAND2_X1 U865 ( .A1(n770), .A2(n769), .ZN(n774) );
  NAND2_X1 U866 ( .A1(G107), .A2(n863), .ZN(n772) );
  NAND2_X1 U867 ( .A1(G95), .A2(n867), .ZN(n771) );
  NAND2_X1 U868 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U869 ( .A1(n774), .A2(n773), .ZN(n860) );
  XOR2_X1 U870 ( .A(KEYINPUT82), .B(G1991), .Z(n907) );
  NOR2_X1 U871 ( .A1(n860), .A2(n907), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n863), .A2(G117), .ZN(n775) );
  XOR2_X1 U873 ( .A(KEYINPUT83), .B(n775), .Z(n777) );
  NAND2_X1 U874 ( .A1(n864), .A2(G129), .ZN(n776) );
  NAND2_X1 U875 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U876 ( .A(KEYINPUT84), .B(n778), .ZN(n782) );
  NAND2_X1 U877 ( .A1(G105), .A2(n867), .ZN(n779) );
  XNOR2_X1 U878 ( .A(n779), .B(KEYINPUT85), .ZN(n780) );
  XNOR2_X1 U879 ( .A(n780), .B(KEYINPUT38), .ZN(n781) );
  NOR2_X1 U880 ( .A1(n782), .A2(n781), .ZN(n784) );
  NAND2_X1 U881 ( .A1(n869), .A2(G141), .ZN(n783) );
  NAND2_X1 U882 ( .A1(n784), .A2(n783), .ZN(n875) );
  AND2_X1 U883 ( .A1(G1996), .A2(n875), .ZN(n785) );
  NOR2_X1 U884 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U885 ( .A(KEYINPUT86), .B(n787), .ZN(n997) );
  XNOR2_X1 U886 ( .A(n804), .B(KEYINPUT87), .ZN(n788) );
  NOR2_X1 U887 ( .A1(n997), .A2(n788), .ZN(n794) );
  INV_X1 U888 ( .A(n794), .ZN(n789) );
  NAND2_X1 U889 ( .A1(n790), .A2(n789), .ZN(n807) );
  NOR2_X1 U890 ( .A1(G1996), .A2(n875), .ZN(n995) );
  NOR2_X1 U891 ( .A1(G1986), .A2(G290), .ZN(n791) );
  AND2_X1 U892 ( .A1(n860), .A2(n907), .ZN(n991) );
  NOR2_X1 U893 ( .A1(n791), .A2(n991), .ZN(n792) );
  XOR2_X1 U894 ( .A(KEYINPUT101), .B(n792), .Z(n793) );
  NOR2_X1 U895 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U896 ( .A(n795), .B(KEYINPUT102), .ZN(n796) );
  NOR2_X1 U897 ( .A1(n995), .A2(n796), .ZN(n797) );
  XNOR2_X1 U898 ( .A(n797), .B(KEYINPUT39), .ZN(n799) );
  NAND2_X1 U899 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U900 ( .A(KEYINPUT103), .B(n800), .Z(n802) );
  NAND2_X1 U901 ( .A1(n878), .A2(n801), .ZN(n988) );
  NAND2_X1 U902 ( .A1(n802), .A2(n988), .ZN(n803) );
  NAND2_X1 U903 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U904 ( .A(n805), .B(KEYINPUT104), .ZN(n806) );
  NAND2_X1 U905 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U906 ( .A(n808), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U907 ( .A1(n809), .A2(G2106), .ZN(n810) );
  XNOR2_X1 U908 ( .A(n810), .B(KEYINPUT106), .ZN(G217) );
  AND2_X1 U909 ( .A1(G15), .A2(G2), .ZN(n811) );
  NAND2_X1 U910 ( .A1(G661), .A2(n811), .ZN(G259) );
  NAND2_X1 U911 ( .A1(G3), .A2(G1), .ZN(n813) );
  NAND2_X1 U912 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U913 ( .A(KEYINPUT107), .B(n814), .Z(G188) );
  XOR2_X1 U914 ( .A(G96), .B(KEYINPUT108), .Z(G221) );
  NOR2_X1 U915 ( .A1(n816), .A2(n815), .ZN(G325) );
  XNOR2_X1 U916 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  XOR2_X1 U917 ( .A(KEYINPUT110), .B(n817), .Z(G319) );
  XOR2_X1 U918 ( .A(KEYINPUT42), .B(G2090), .Z(n819) );
  XNOR2_X1 U919 ( .A(G2078), .B(G2084), .ZN(n818) );
  XNOR2_X1 U920 ( .A(n819), .B(n818), .ZN(n820) );
  XOR2_X1 U921 ( .A(n820), .B(G2100), .Z(n822) );
  XNOR2_X1 U922 ( .A(G2067), .B(G2072), .ZN(n821) );
  XNOR2_X1 U923 ( .A(n822), .B(n821), .ZN(n826) );
  XOR2_X1 U924 ( .A(G2096), .B(KEYINPUT43), .Z(n824) );
  XNOR2_X1 U925 ( .A(KEYINPUT111), .B(G2678), .ZN(n823) );
  XNOR2_X1 U926 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U927 ( .A(n826), .B(n825), .Z(G227) );
  XNOR2_X1 U928 ( .A(G1981), .B(KEYINPUT112), .ZN(n836) );
  XOR2_X1 U929 ( .A(G1986), .B(G1966), .Z(n828) );
  XNOR2_X1 U930 ( .A(G1961), .B(G1956), .ZN(n827) );
  XNOR2_X1 U931 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U932 ( .A(G1991), .B(G1976), .Z(n830) );
  XNOR2_X1 U933 ( .A(G1996), .B(G1971), .ZN(n829) );
  XNOR2_X1 U934 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U935 ( .A(n832), .B(n831), .Z(n834) );
  XNOR2_X1 U936 ( .A(G2474), .B(KEYINPUT41), .ZN(n833) );
  XNOR2_X1 U937 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U938 ( .A(n836), .B(n835), .ZN(G229) );
  NAND2_X1 U939 ( .A1(G112), .A2(n863), .ZN(n837) );
  XNOR2_X1 U940 ( .A(n837), .B(KEYINPUT114), .ZN(n841) );
  XOR2_X1 U941 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n839) );
  NAND2_X1 U942 ( .A1(G124), .A2(n864), .ZN(n838) );
  XNOR2_X1 U943 ( .A(n839), .B(n838), .ZN(n840) );
  NAND2_X1 U944 ( .A1(n841), .A2(n840), .ZN(n845) );
  NAND2_X1 U945 ( .A1(G100), .A2(n867), .ZN(n843) );
  NAND2_X1 U946 ( .A1(G136), .A2(n869), .ZN(n842) );
  NAND2_X1 U947 ( .A1(n843), .A2(n842), .ZN(n844) );
  NOR2_X1 U948 ( .A1(n845), .A2(n844), .ZN(G162) );
  XOR2_X1 U949 ( .A(n987), .B(G162), .Z(n847) );
  XNOR2_X1 U950 ( .A(G160), .B(G164), .ZN(n846) );
  XNOR2_X1 U951 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U952 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n849) );
  XNOR2_X1 U953 ( .A(KEYINPUT117), .B(KEYINPUT116), .ZN(n848) );
  XNOR2_X1 U954 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U955 ( .A(n851), .B(n850), .Z(n862) );
  NAND2_X1 U956 ( .A1(G103), .A2(n867), .ZN(n854) );
  NAND2_X1 U957 ( .A1(G139), .A2(n852), .ZN(n853) );
  NAND2_X1 U958 ( .A1(n854), .A2(n853), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G115), .A2(n863), .ZN(n856) );
  NAND2_X1 U960 ( .A1(G127), .A2(n864), .ZN(n855) );
  NAND2_X1 U961 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U962 ( .A(KEYINPUT47), .B(n857), .Z(n858) );
  NOR2_X1 U963 ( .A1(n859), .A2(n858), .ZN(n980) );
  XNOR2_X1 U964 ( .A(n860), .B(n980), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(n880) );
  NAND2_X1 U966 ( .A1(G118), .A2(n863), .ZN(n866) );
  NAND2_X1 U967 ( .A1(G130), .A2(n864), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n874) );
  NAND2_X1 U969 ( .A1(n867), .A2(G106), .ZN(n868) );
  XOR2_X1 U970 ( .A(KEYINPUT115), .B(n868), .Z(n871) );
  NAND2_X1 U971 ( .A1(n869), .A2(G142), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U973 ( .A(n872), .B(KEYINPUT45), .Z(n873) );
  NOR2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n876) );
  XNOR2_X1 U975 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U976 ( .A(n878), .B(n877), .Z(n879) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n881) );
  NOR2_X1 U978 ( .A1(G37), .A2(n881), .ZN(G395) );
  XNOR2_X1 U979 ( .A(n924), .B(G301), .ZN(n882) );
  XNOR2_X1 U980 ( .A(n882), .B(n927), .ZN(n885) );
  XNOR2_X1 U981 ( .A(G286), .B(n883), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n886) );
  NOR2_X1 U983 ( .A1(G37), .A2(n886), .ZN(G397) );
  XOR2_X1 U984 ( .A(KEYINPUT105), .B(G2451), .Z(n888) );
  XNOR2_X1 U985 ( .A(G2446), .B(G2427), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n895) );
  XOR2_X1 U987 ( .A(G2438), .B(G2435), .Z(n890) );
  XNOR2_X1 U988 ( .A(G2443), .B(G2430), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U990 ( .A(n891), .B(G2454), .Z(n893) );
  XNOR2_X1 U991 ( .A(G1341), .B(G1348), .ZN(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n896) );
  NAND2_X1 U994 ( .A1(n896), .A2(G14), .ZN(n902) );
  NAND2_X1 U995 ( .A1(n902), .A2(G319), .ZN(n899) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n897) );
  XNOR2_X1 U997 ( .A(KEYINPUT49), .B(n897), .ZN(n898) );
  NOR2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n901) );
  NOR2_X1 U999 ( .A1(G395), .A2(G397), .ZN(n900) );
  NAND2_X1 U1000 ( .A1(n901), .A2(n900), .ZN(G225) );
  XOR2_X1 U1001 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  INV_X1 U1003 ( .A(G120), .ZN(G236) );
  INV_X1 U1004 ( .A(G69), .ZN(G235) );
  INV_X1 U1005 ( .A(G108), .ZN(G238) );
  INV_X1 U1006 ( .A(n902), .ZN(G401) );
  XNOR2_X1 U1007 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n1002) );
  XNOR2_X1 U1008 ( .A(G1996), .B(G32), .ZN(n904) );
  XNOR2_X1 U1009 ( .A(G33), .B(G2072), .ZN(n903) );
  NOR2_X1 U1010 ( .A1(n904), .A2(n903), .ZN(n913) );
  XOR2_X1 U1011 ( .A(G2067), .B(G26), .Z(n905) );
  NAND2_X1 U1012 ( .A1(n905), .A2(G28), .ZN(n911) );
  XOR2_X1 U1013 ( .A(n906), .B(G27), .Z(n909) );
  XNOR2_X1 U1014 ( .A(n907), .B(G25), .ZN(n908) );
  NAND2_X1 U1015 ( .A1(n909), .A2(n908), .ZN(n910) );
  NOR2_X1 U1016 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1017 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1018 ( .A(n914), .B(KEYINPUT53), .ZN(n917) );
  XOR2_X1 U1019 ( .A(G2084), .B(KEYINPUT54), .Z(n915) );
  XNOR2_X1 U1020 ( .A(G34), .B(n915), .ZN(n916) );
  NAND2_X1 U1021 ( .A1(n917), .A2(n916), .ZN(n919) );
  XNOR2_X1 U1022 ( .A(G35), .B(G2090), .ZN(n918) );
  NOR2_X1 U1023 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1024 ( .A(n1002), .B(n920), .Z(n922) );
  INV_X1 U1025 ( .A(G29), .ZN(n921) );
  NAND2_X1 U1026 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1027 ( .A1(n923), .A2(G11), .ZN(n979) );
  XNOR2_X1 U1028 ( .A(G16), .B(KEYINPUT56), .ZN(n949) );
  XOR2_X1 U1029 ( .A(n924), .B(G1348), .Z(n925) );
  NOR2_X1 U1030 ( .A1(n926), .A2(n925), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(G301), .B(G1961), .ZN(n929) );
  XNOR2_X1 U1032 ( .A(n927), .B(G1341), .ZN(n928) );
  NOR2_X1 U1033 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(n932), .B(G1956), .ZN(n934) );
  NAND2_X1 U1036 ( .A1(G1971), .A2(G303), .ZN(n933) );
  NAND2_X1 U1037 ( .A1(n934), .A2(n933), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1040 ( .A(KEYINPUT121), .B(n939), .ZN(n940) );
  NOR2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(KEYINPUT122), .B(n942), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(G168), .B(G1966), .ZN(n944) );
  NAND2_X1 U1044 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1045 ( .A(KEYINPUT57), .B(n945), .ZN(n946) );
  NAND2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n977) );
  INV_X1 U1048 ( .A(G16), .ZN(n975) );
  XNOR2_X1 U1049 ( .A(G1971), .B(G22), .ZN(n951) );
  XNOR2_X1 U1050 ( .A(G23), .B(G1976), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n953) );
  XOR2_X1 U1052 ( .A(G1986), .B(G24), .Z(n952) );
  NAND2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n955) );
  XOR2_X1 U1054 ( .A(KEYINPUT58), .B(KEYINPUT124), .Z(n954) );
  XNOR2_X1 U1055 ( .A(n955), .B(n954), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(G1961), .B(G5), .ZN(n957) );
  XNOR2_X1 U1057 ( .A(G21), .B(G1966), .ZN(n956) );
  NOR2_X1 U1058 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1059 ( .A1(n959), .A2(n958), .ZN(n971) );
  XOR2_X1 U1060 ( .A(G1348), .B(KEYINPUT59), .Z(n960) );
  XNOR2_X1 U1061 ( .A(G4), .B(n960), .ZN(n968) );
  XOR2_X1 U1062 ( .A(G1341), .B(G19), .Z(n963) );
  XNOR2_X1 U1063 ( .A(n961), .B(G20), .ZN(n962) );
  NAND2_X1 U1064 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1065 ( .A(G6), .B(G1981), .ZN(n964) );
  NOR2_X1 U1066 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1067 ( .A(n966), .B(KEYINPUT123), .ZN(n967) );
  NOR2_X1 U1068 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1069 ( .A(n969), .B(KEYINPUT60), .Z(n970) );
  NOR2_X1 U1070 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1071 ( .A(KEYINPUT61), .B(n972), .Z(n973) );
  XNOR2_X1 U1072 ( .A(KEYINPUT125), .B(n973), .ZN(n974) );
  NAND2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n1007) );
  XOR2_X1 U1076 ( .A(G2072), .B(n980), .Z(n982) );
  XOR2_X1 U1077 ( .A(G164), .B(G2078), .Z(n981) );
  NOR2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1079 ( .A(KEYINPUT50), .B(n983), .Z(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n993) );
  XOR2_X1 U1081 ( .A(G2084), .B(G160), .Z(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n1000) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1088 ( .A(KEYINPUT51), .B(n996), .Z(n998) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(KEYINPUT52), .B(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(G29), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(KEYINPUT120), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(n1008), .B(KEYINPUT62), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(KEYINPUT126), .B(n1009), .ZN(G150) );
  INV_X1 U1098 ( .A(G150), .ZN(G311) );
endmodule

