//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT31), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT67), .B1(new_n189), .B2(G134), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT67), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G137), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G134), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT11), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n190), .A2(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT66), .B(G131), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n189), .A2(KEYINPUT65), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G137), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT11), .A2(G134), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n196), .A2(new_n197), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  INV_X1    g019(.A(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G146), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n205), .B(new_n207), .C1(KEYINPUT1), .C2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(G134), .B1(new_n198), .B2(new_n200), .ZN(new_n210));
  INV_X1    g024(.A(new_n194), .ZN(new_n211));
  OAI21_X1  g025(.A(G131), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT1), .B1(new_n206), .B2(G146), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n206), .A2(G146), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n204), .A2(G143), .ZN(new_n215));
  OAI211_X1 g029(.A(G128), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AND4_X1   g030(.A1(new_n203), .A2(new_n209), .A3(new_n212), .A4(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n205), .A2(new_n207), .A3(KEYINPUT0), .A4(G128), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT0), .B(G128), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n190), .A2(new_n193), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n194), .A2(new_n195), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n202), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G131), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n221), .B1(new_n225), .B2(new_n203), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n188), .B1(new_n217), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT2), .ZN(new_n228));
  INV_X1    g042(.A(G113), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(KEYINPUT68), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(KEYINPUT2), .B2(G113), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n230), .A2(new_n232), .B1(KEYINPUT2), .B2(G113), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT69), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G119), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n238), .A3(G116), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n234), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n233), .A2(new_n239), .A3(new_n241), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n227), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n221), .ZN(new_n247));
  AND4_X1   g061(.A1(new_n197), .A2(new_n222), .A3(new_n202), .A4(new_n223), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n196), .B2(new_n202), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n247), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n216), .A2(new_n209), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n203), .A3(new_n212), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(KEYINPUT30), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n251), .A2(KEYINPUT70), .A3(KEYINPUT30), .A4(new_n253), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n246), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n234), .A2(new_n242), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n233), .B1(new_n239), .B2(new_n241), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n251), .A2(new_n261), .A3(new_n253), .ZN(new_n262));
  INV_X1    g076(.A(G237), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(G210), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT27), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G101), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n187), .B1(new_n258), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n256), .A2(new_n257), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n251), .A2(new_n253), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n261), .B1(new_n272), .B2(new_n188), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n269), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(KEYINPUT31), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n245), .B1(new_n217), .B2(new_n226), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(new_n262), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n217), .A2(new_n226), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT28), .B1(new_n280), .B2(new_n261), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT71), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n217), .A2(new_n226), .A3(new_n245), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n261), .B1(new_n251), .B2(new_n253), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT28), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n268), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n270), .A2(new_n276), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g104(.A1(G472), .A2(G902), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT32), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT31), .B1(new_n274), .B2(new_n275), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n187), .B(new_n269), .C1(new_n271), .C2(new_n273), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n268), .B1(new_n282), .B2(new_n287), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n294), .B(new_n291), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT74), .B(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n283), .B2(new_n284), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT73), .B1(new_n272), .B2(new_n245), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n281), .B1(new_n305), .B2(KEYINPUT28), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n289), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n301), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n283), .B1(new_n271), .B2(new_n273), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n310), .B1(new_n311), .B2(new_n268), .ZN(new_n312));
  OAI211_X1 g126(.A(KEYINPUT72), .B(new_n289), .C1(new_n258), .C2(new_n283), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n282), .A2(new_n287), .A3(new_n268), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n307), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n309), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n293), .A2(new_n299), .B1(new_n317), .B2(G472), .ZN(new_n318));
  XNOR2_X1  g132(.A(G125), .B(G140), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n320), .A2(KEYINPUT16), .A3(G140), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n319), .A2(KEYINPUT16), .B1(new_n321), .B2(KEYINPUT76), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT16), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(G125), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n322), .A2(G146), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n319), .A2(new_n204), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G110), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT69), .B(G119), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(G128), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n235), .A2(new_n208), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n333), .B2(new_n208), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n331), .B(new_n334), .C1(new_n336), .C2(new_n332), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n236), .A2(new_n238), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G128), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT24), .B(G110), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n339), .A2(KEYINPUT77), .A3(new_n335), .A4(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n335), .B(new_n340), .C1(new_n333), .C2(new_n208), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n337), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT78), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n337), .A2(new_n347), .A3(new_n341), .A4(new_n344), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n330), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n334), .B1(new_n336), .B2(new_n332), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G110), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(KEYINPUT75), .A3(G110), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n336), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n357), .A2(new_n340), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT76), .A4(G125), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n324), .A2(G125), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n320), .A2(G140), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n327), .B(new_n359), .C1(new_n362), .C2(new_n323), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n204), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n328), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n356), .A2(new_n358), .A3(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT22), .B(G137), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n350), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n369), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n365), .A2(new_n358), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n354), .B2(new_n355), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n371), .B1(new_n349), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(new_n300), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT25), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n370), .A2(new_n374), .A3(KEYINPUT25), .A4(new_n300), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G217), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n300), .B2(G234), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n370), .A2(new_n374), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n381), .A2(G902), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n318), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n388));
  INV_X1    g202(.A(G104), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT3), .B1(new_n389), .B2(G107), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n389), .A2(G107), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n396), .A3(G101), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n395), .A2(G101), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n390), .A2(new_n393), .A3(new_n399), .A4(new_n394), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT4), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n247), .B(new_n397), .C1(new_n398), .C2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n248), .A2(new_n250), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n389), .A2(G107), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n392), .A2(G104), .ZN(new_n405));
  OAI21_X1  g219(.A(G101), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n216), .A2(new_n400), .A3(new_n406), .A4(new_n209), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n400), .A2(new_n406), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n252), .A2(new_n410), .A3(KEYINPUT10), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n402), .A2(new_n403), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n216), .A2(new_n209), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n400), .A2(new_n406), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n407), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n225), .A2(new_n203), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n416), .A2(KEYINPUT12), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(KEYINPUT12), .B1(new_n416), .B2(new_n417), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n412), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G110), .B(G140), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n264), .A2(G227), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n402), .A2(new_n409), .A3(new_n411), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n417), .ZN(new_n426));
  INV_X1    g240(.A(new_n423), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n412), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(G902), .B1(new_n424), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G469), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n388), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n412), .A2(new_n427), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n420), .A2(new_n423), .B1(new_n432), .B2(new_n426), .ZN(new_n433));
  OAI211_X1 g247(.A(KEYINPUT81), .B(G469), .C1(new_n433), .C2(G902), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n418), .A2(new_n419), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n412), .A2(new_n427), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n427), .B1(new_n426), .B2(new_n412), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n430), .B(new_n300), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n431), .A2(new_n434), .A3(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT9), .B(G234), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT79), .ZN(new_n442));
  INV_X1    g256(.A(G902), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G221), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT80), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT82), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n440), .A2(KEYINPUT82), .A3(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n206), .A2(G128), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n208), .A2(G143), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT94), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G128), .B(G143), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(KEYINPUT94), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n459), .A3(G134), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT94), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT94), .B1(new_n453), .B2(new_n454), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n192), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT95), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT95), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n460), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G122), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G116), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n392), .B1(new_n469), .B2(KEYINPUT14), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n240), .A2(G122), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n470), .B(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n465), .A2(new_n467), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n442), .A2(G217), .A3(new_n264), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n458), .A2(KEYINPUT13), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n478), .B(G134), .C1(KEYINPUT13), .C2(new_n453), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n472), .B(G107), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n479), .A2(new_n480), .A3(new_n463), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n475), .A2(new_n477), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT96), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT96), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n475), .A2(new_n485), .A3(new_n477), .A4(new_n482), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n475), .A2(new_n482), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n476), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n300), .ZN(new_n490));
  INV_X1    g304(.A(G478), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n490), .B(new_n492), .Z(new_n493));
  XNOR2_X1  g307(.A(G113), .B(G122), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(new_n389), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n263), .A2(new_n264), .A3(G214), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n206), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n263), .A2(new_n264), .A3(G143), .A4(G214), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT18), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(new_n249), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n362), .A2(G146), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n329), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n499), .ZN(new_n506));
  INV_X1    g320(.A(new_n501), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(KEYINPUT88), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT88), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n499), .B2(new_n501), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n505), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n197), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n499), .A2(KEYINPUT17), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n364), .A2(new_n328), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT90), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n364), .A2(new_n328), .A3(KEYINPUT90), .A4(new_n514), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n506), .A2(new_n197), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n499), .A2(new_n513), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n495), .B(new_n512), .C1(new_n517), .C2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n495), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n521), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT19), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n362), .A2(KEYINPUT89), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT89), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT19), .B1(new_n319), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n204), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n526), .A2(new_n328), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n525), .B1(new_n532), .B2(new_n511), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n524), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G475), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n443), .ZN(new_n536));
  OAI211_X1 g350(.A(KEYINPUT91), .B(KEYINPUT20), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n524), .B2(new_n533), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT20), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n524), .A2(new_n533), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT92), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT20), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n542), .B(new_n544), .C1(new_n543), .C2(new_n536), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n537), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n512), .B1(new_n517), .B2(new_n523), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n547), .A2(new_n525), .ZN(new_n548));
  INV_X1    g362(.A(new_n524), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n443), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  XOR2_X1   g364(.A(KEYINPUT93), .B(G475), .Z(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n493), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(G210), .B1(G237), .B2(G902), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT86), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n216), .A2(new_n320), .A3(new_n209), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n218), .B(G125), .C1(new_n219), .C2(new_n220), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n264), .A2(G224), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n239), .A2(KEYINPUT5), .A3(new_n241), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n562), .B(G113), .C1(KEYINPUT5), .C2(new_n239), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n563), .A2(new_n244), .A3(new_n410), .ZN(new_n564));
  XNOR2_X1  g378(.A(G110), .B(G122), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n397), .B1(new_n259), .B2(new_n260), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n398), .A2(new_n401), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT6), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n565), .B(KEYINPUT83), .Z(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(KEYINPUT6), .A3(new_n571), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n561), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n563), .A2(new_n244), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n414), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT84), .A3(new_n564), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n565), .B(KEYINPUT8), .Z(new_n579));
  AOI21_X1  g393(.A(new_n410), .B1(new_n563), .B2(new_n244), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT85), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n559), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n556), .A2(new_n557), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n559), .A2(KEYINPUT7), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n568), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n443), .B1(new_n583), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n555), .B1(new_n575), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n568), .A2(KEYINPUT6), .B1(new_n570), .B2(new_n571), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n570), .A2(KEYINPUT6), .A3(new_n571), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n560), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n568), .A2(new_n588), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n578), .A2(new_n582), .ZN(new_n596));
  AOI21_X1  g410(.A(G902), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n594), .A2(new_n597), .A3(new_n554), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n591), .A2(KEYINPUT87), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT87), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n594), .A2(new_n597), .A3(new_n600), .A4(new_n554), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n264), .A2(G952), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(G234), .B2(G237), .ZN(new_n603));
  AOI211_X1 g417(.A(new_n264), .B(new_n300), .C1(G234), .C2(G237), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT21), .B(G898), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G214), .B1(G237), .B2(G902), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n599), .A2(new_n601), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n553), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n387), .A2(new_n452), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  AOI21_X1  g427(.A(new_n554), .B1(new_n594), .B2(new_n597), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n608), .B1(new_n614), .B2(KEYINPUT97), .ZN(new_n615));
  INV_X1    g429(.A(new_n554), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n575), .B2(new_n590), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT97), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n618), .A3(new_n598), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n606), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n301), .A2(new_n491), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n475), .A2(KEYINPUT98), .A3(new_n477), .A4(new_n482), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n488), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT98), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n483), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT33), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n484), .A2(new_n488), .A3(new_n630), .A4(new_n486), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n624), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n632), .A2(new_n633), .B1(new_n491), .B2(new_n490), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n629), .A2(new_n631), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n623), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT99), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n546), .A2(new_n552), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n622), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n477), .B1(new_n475), .B2(new_n482), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n475), .A2(new_n477), .A3(new_n482), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n641), .B1(new_n642), .B2(KEYINPUT98), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n483), .A2(new_n627), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n630), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n631), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n633), .B(new_n623), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n490), .A2(new_n491), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n632), .A2(new_n633), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n639), .B(new_n622), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n621), .B1(new_n640), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(G472), .B1(new_n290), .B2(new_n301), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n291), .B1(new_n297), .B2(new_n298), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n386), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n452), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT34), .B(G104), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  INV_X1    g475(.A(new_n606), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n615), .A2(new_n619), .A3(new_n552), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n490), .B(new_n492), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n539), .A2(new_n540), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n537), .A2(new_n541), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n657), .A2(new_n452), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT35), .B(G107), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  NAND2_X1  g485(.A1(new_n350), .A2(new_n366), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n371), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n674), .A2(new_n384), .ZN(new_n675));
  INV_X1    g489(.A(new_n381), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n377), .B2(new_n378), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n656), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n611), .A2(new_n679), .A3(new_n452), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  NAND2_X1  g496(.A1(new_n293), .A2(new_n299), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n317), .A2(G472), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n678), .A2(new_n620), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n604), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n688), .A2(new_n603), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n552), .A2(new_n689), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n690), .A2(new_n664), .A3(new_n666), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n452), .A2(new_n685), .A3(new_n686), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT101), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n619), .B(new_n615), .C1(new_n675), .C2(new_n677), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n318), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT101), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n695), .A2(new_n696), .A3(new_n452), .A4(new_n691), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G128), .ZN(G30));
  XNOR2_X1  g513(.A(new_n689), .B(KEYINPUT39), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n452), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT40), .Z(new_n702));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n703));
  INV_X1    g517(.A(G472), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n305), .A2(new_n268), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(G902), .ZN(new_n706));
  INV_X1    g520(.A(new_n311), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n268), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n704), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n703), .B1(new_n683), .B2(new_n710), .ZN(new_n711));
  AOI211_X1 g525(.A(KEYINPUT102), .B(new_n709), .C1(new_n293), .C2(new_n299), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n678), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n598), .A2(KEYINPUT87), .ZN(new_n716));
  INV_X1    g530(.A(new_n555), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n717), .B1(new_n594), .B2(new_n597), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n601), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n719), .B(KEYINPUT38), .Z(new_n720));
  AND4_X1   g534(.A1(new_n639), .A2(new_n720), .A3(new_n664), .A4(new_n607), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n702), .A2(new_n715), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G143), .ZN(G45));
  OAI211_X1 g537(.A(new_n639), .B(new_n689), .C1(new_n649), .C2(new_n650), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n452), .A3(new_n685), .A4(new_n686), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G146), .ZN(G48));
  OAI21_X1  g541(.A(new_n639), .B1(new_n649), .B2(new_n650), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT100), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n651), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n437), .A2(new_n438), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n430), .B1(new_n731), .B2(new_n300), .ZN(new_n732));
  INV_X1    g546(.A(new_n445), .ZN(new_n733));
  INV_X1    g547(.A(new_n439), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n730), .A2(new_n387), .A3(new_n621), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT41), .B(G113), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  AOI22_X1  g552(.A1(new_n379), .A2(new_n381), .B1(new_n384), .B2(new_n383), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n685), .A2(new_n668), .A3(new_n739), .A4(new_n735), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G116), .ZN(G18));
  NOR2_X1   g555(.A1(new_n318), .A2(new_n678), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n735), .A2(new_n619), .A3(new_n662), .A4(new_n615), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n553), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  NOR2_X1   g560(.A1(new_n306), .A2(new_n268), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n291), .B1(new_n747), .B2(new_n297), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n739), .A2(new_n654), .A3(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n639), .A2(new_n664), .A3(new_n619), .A4(new_n615), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT103), .ZN(new_n752));
  NOR4_X1   g566(.A1(new_n732), .A2(new_n734), .A3(new_n733), .A4(new_n606), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n749), .A2(new_n751), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n739), .A2(new_n753), .A3(new_n654), .A4(new_n748), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT103), .B1(new_n755), .B2(new_n750), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  NAND2_X1  g572(.A1(new_n654), .A2(new_n748), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n678), .ZN(new_n760));
  INV_X1    g574(.A(new_n735), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n620), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n725), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  OAI21_X1  g578(.A(G469), .B1(new_n433), .B2(G902), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(KEYINPUT104), .A3(new_n439), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT104), .B1(new_n765), .B2(new_n439), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n445), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n719), .A2(new_n607), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n387), .A2(new_n725), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT42), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n387), .A2(KEYINPUT42), .A3(new_n725), .A4(new_n771), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  NAND4_X1  g591(.A1(new_n771), .A2(new_n685), .A3(new_n739), .A4(new_n691), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT105), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT105), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n387), .A2(new_n780), .A3(new_n691), .A4(new_n771), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G134), .ZN(G36));
  NAND2_X1  g597(.A1(new_n424), .A2(new_n428), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT106), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n430), .B1(new_n784), .B2(new_n785), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(G469), .A2(G902), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n734), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n789), .A2(KEYINPUT46), .A3(new_n790), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n733), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n700), .ZN(new_n796));
  XOR2_X1   g610(.A(new_n796), .B(KEYINPUT107), .Z(new_n797));
  INV_X1    g611(.A(new_n638), .ZN(new_n798));
  OR3_X1    g612(.A1(new_n798), .A2(KEYINPUT43), .A3(new_n639), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT43), .B1(new_n798), .B2(new_n639), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n799), .A2(new_n656), .A3(new_n714), .A4(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT44), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n770), .B(KEYINPUT108), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n797), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  XNOR2_X1  g619(.A(new_n795), .B(KEYINPUT47), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n685), .A2(new_n739), .A3(new_n770), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n725), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G140), .ZN(G42));
  INV_X1    g623(.A(new_n770), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n735), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n799), .A2(new_n603), .A3(new_n800), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n387), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT48), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n602), .B(KEYINPUT116), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n713), .A2(new_n739), .A3(new_n603), .A4(new_n812), .ZN(new_n819));
  INV_X1    g633(.A(new_n730), .ZN(new_n820));
  INV_X1    g634(.A(new_n762), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n799), .A2(new_n603), .A3(new_n749), .A4(new_n800), .ZN(new_n822));
  OAI221_X1 g636(.A(new_n818), .B1(new_n819), .B2(new_n820), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n816), .B1(new_n817), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n735), .A2(new_n608), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT114), .Z(new_n826));
  NOR3_X1   g640(.A1(new_n822), .A2(new_n720), .A3(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT50), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n813), .A2(new_n678), .A3(new_n759), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n819), .A2(new_n639), .A3(new_n638), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n803), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n822), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n732), .A2(new_n734), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT109), .Z(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n447), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n834), .B1(new_n806), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT51), .ZN(new_n839));
  OAI221_X1 g653(.A(new_n824), .B1(new_n817), .B2(new_n823), .C1(new_n832), .C2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n832), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n828), .A2(KEYINPUT115), .A3(new_n831), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n838), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n840), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n726), .A2(new_n763), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n445), .B(new_n689), .C1(new_n767), .C2(new_n768), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n849), .A2(new_n750), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n850), .B(new_n678), .C1(new_n711), .C2(new_n712), .ZN(new_n851));
  AND4_X1   g665(.A1(KEYINPUT52), .A2(new_n698), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n851), .A2(new_n726), .A3(new_n763), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(new_n853), .B2(new_n698), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n736), .A2(new_n757), .A3(new_n740), .A4(new_n745), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n771), .A2(new_n725), .A3(new_n760), .ZN(new_n858));
  INV_X1    g672(.A(new_n742), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n493), .A2(new_n666), .A3(new_n690), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n452), .A2(new_n810), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n858), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n862), .B1(new_n781), .B2(new_n779), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n634), .A2(new_n637), .A3(new_n639), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n864), .A2(new_n553), .ZN(new_n865));
  INV_X1    g679(.A(new_n610), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n657), .A3(new_n452), .A4(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n867), .A2(new_n612), .A3(new_n680), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n857), .A2(new_n863), .A3(new_n776), .A4(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n847), .B1(new_n855), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  INV_X1    g685(.A(new_n698), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n851), .A2(new_n726), .A3(new_n763), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n853), .A2(KEYINPUT52), .A3(new_n698), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n862), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n868), .A2(new_n877), .A3(new_n782), .A4(KEYINPUT53), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NOR4_X1   g693(.A1(new_n318), .A2(new_n769), .A3(new_n770), .A4(new_n386), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT42), .B1(new_n880), .B2(new_n725), .ZN(new_n881));
  INV_X1    g695(.A(new_n775), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT112), .B1(new_n883), .B2(new_n856), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n387), .A2(new_n735), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n653), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n745), .A2(new_n740), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT112), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n889), .A3(new_n757), .A4(new_n776), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n876), .A2(new_n879), .A3(new_n884), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n870), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(KEYINPUT54), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n893), .A2(KEYINPUT113), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n868), .A2(new_n877), .A3(new_n782), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n895), .A2(new_n883), .A3(new_n856), .ZN(new_n896));
  INV_X1    g710(.A(new_n847), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(new_n876), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n876), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n898), .A2(KEYINPUT111), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(KEYINPUT111), .B2(new_n898), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT54), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n893), .A2(KEYINPUT113), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n846), .A2(new_n894), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n905), .B1(G952), .B2(G953), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n836), .B(KEYINPUT49), .Z(new_n907));
  NOR4_X1   g721(.A1(new_n720), .A2(new_n386), .A3(new_n446), .A4(new_n608), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n798), .A2(new_n639), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n907), .A2(new_n713), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n906), .A2(new_n910), .ZN(G75));
  NOR2_X1   g725(.A1(new_n264), .A2(G952), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n884), .A2(new_n890), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n878), .B1(new_n874), .B2(new_n875), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n899), .A2(new_n847), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(new_n300), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT56), .B1(new_n916), .B2(new_n616), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n592), .A2(new_n593), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n560), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT55), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n916), .A2(new_n555), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n920), .B(KEYINPUT119), .ZN(new_n923));
  XOR2_X1   g737(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n912), .B(new_n921), .C1(new_n922), .C2(new_n925), .ZN(G51));
  XNOR2_X1  g740(.A(new_n892), .B(KEYINPUT54), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n790), .B(KEYINPUT57), .Z(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT120), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n927), .A2(KEYINPUT120), .A3(new_n928), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n731), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n916), .A2(new_n787), .A3(new_n788), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n912), .B1(new_n933), .B2(new_n934), .ZN(G54));
  INV_X1    g749(.A(new_n912), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n916), .A2(KEYINPUT58), .A3(G475), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(new_n542), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n542), .B2(new_n937), .ZN(G60));
  NAND3_X1  g753(.A1(new_n894), .A2(new_n903), .A3(new_n904), .ZN(new_n940));
  NAND2_X1  g754(.A1(G478), .A2(G902), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT59), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n635), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n927), .A2(new_n635), .A3(new_n942), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n943), .A2(new_n912), .A3(new_n944), .ZN(G63));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT123), .ZN(new_n947));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT121), .Z(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT60), .Z(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n870), .B2(new_n891), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n947), .B1(new_n952), .B2(new_n383), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n912), .B1(new_n952), .B2(new_n674), .ZN(new_n954));
  INV_X1    g768(.A(new_n383), .ZN(new_n955));
  OAI211_X1 g769(.A(KEYINPUT123), .B(new_n955), .C1(new_n915), .C2(new_n951), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT61), .A4(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n955), .B1(new_n915), .B2(new_n951), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT61), .B1(new_n954), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n959), .B2(KEYINPUT122), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  AOI211_X1 g775(.A(new_n961), .B(KEYINPUT61), .C1(new_n954), .C2(new_n958), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n946), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n892), .A2(new_n674), .A3(new_n950), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n936), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n952), .A2(new_n383), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n961), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n959), .A2(KEYINPUT122), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT124), .A4(new_n957), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n963), .A2(new_n971), .ZN(G66));
  INV_X1    g786(.A(G224), .ZN(new_n973));
  OAI21_X1  g787(.A(G953), .B1(new_n605), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n857), .A2(new_n868), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n976), .B2(G953), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n918), .B1(G898), .B2(new_n264), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(G69));
  NAND3_X1  g793(.A1(new_n387), .A2(new_n865), .A3(new_n810), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n804), .B(new_n808), .C1(new_n701), .C2(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n698), .A2(new_n848), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n722), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT62), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n984), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT125), .ZN(new_n988));
  AOI21_X1  g802(.A(G953), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n271), .A2(new_n227), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n528), .A2(new_n530), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n990), .B(new_n991), .Z(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n264), .B1(G227), .B2(G900), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n797), .A2(new_n387), .A3(new_n751), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n808), .A2(new_n776), .A3(new_n782), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n804), .A2(new_n996), .A3(new_n997), .A4(new_n982), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n264), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n687), .A2(G953), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT126), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n992), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  OR3_X1    g816(.A1(new_n994), .A2(new_n995), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n995), .B1(new_n994), .B2(new_n1002), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(G72));
  NAND3_X1  g819(.A1(new_n986), .A2(new_n976), .A3(new_n988), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  AOI21_X1  g822(.A(new_n708), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1008), .B1(new_n998), .B2(new_n975), .ZN(new_n1010));
  AND3_X1   g824(.A1(new_n1010), .A2(new_n311), .A3(new_n289), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n312), .B(new_n313), .C1(new_n258), .C2(new_n269), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n902), .A2(new_n1008), .A3(new_n1012), .ZN(new_n1013));
  NOR4_X1   g827(.A1(new_n1009), .A2(new_n1011), .A3(new_n1013), .A4(new_n912), .ZN(G57));
endmodule


