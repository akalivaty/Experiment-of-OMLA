

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  XNOR2_X1 U323 ( .A(n439), .B(KEYINPUT65), .ZN(n577) );
  XOR2_X1 U324 ( .A(G85GAT), .B(KEYINPUT73), .Z(n378) );
  NOR2_X1 U325 ( .A1(n578), .A2(n406), .ZN(n407) );
  XNOR2_X1 U326 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U327 ( .A(G43GAT), .B(G134GAT), .Z(n382) );
  XNOR2_X1 U328 ( .A(n457), .B(n456), .ZN(n458) );
  AND2_X1 U329 ( .A1(G226GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U330 ( .A(n295), .B(G183GAT), .Z(n292) );
  INV_X1 U331 ( .A(KEYINPUT25), .ZN(n464) );
  INV_X1 U332 ( .A(n569), .ZN(n400) );
  XNOR2_X1 U333 ( .A(n465), .B(n464), .ZN(n470) );
  AND2_X1 U334 ( .A1(n401), .A2(n400), .ZN(n402) );
  NAND2_X1 U335 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U336 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U337 ( .A(n366), .B(n291), .ZN(n306) );
  NOR2_X1 U338 ( .A1(n589), .A2(n476), .ZN(n477) );
  XNOR2_X1 U339 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U340 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n369) );
  XNOR2_X1 U341 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U342 ( .A(n582), .B(n369), .ZN(n562) );
  INV_X1 U343 ( .A(G43GAT), .ZN(n480) );
  XNOR2_X1 U344 ( .A(n316), .B(n315), .ZN(n507) );
  XNOR2_X1 U345 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n483) );
  XNOR2_X1 U346 ( .A(n480), .B(KEYINPUT40), .ZN(n481) );
  XNOR2_X1 U347 ( .A(n484), .B(n483), .ZN(G1351GAT) );
  XNOR2_X1 U348 ( .A(n482), .B(n481), .ZN(G1330GAT) );
  XOR2_X1 U349 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n294) );
  XNOR2_X1 U350 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U352 ( .A(G169GAT), .B(G176GAT), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n292), .B(n296), .ZN(n307) );
  XNOR2_X1 U354 ( .A(G99GAT), .B(G71GAT), .ZN(n297) );
  XNOR2_X1 U355 ( .A(n297), .B(G120GAT), .ZN(n354) );
  XOR2_X1 U356 ( .A(KEYINPUT20), .B(n354), .Z(n299) );
  NAND2_X1 U357 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U358 ( .A(n299), .B(n298), .ZN(n302) );
  XNOR2_X1 U359 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n300) );
  XOR2_X1 U360 ( .A(G113GAT), .B(KEYINPUT0), .Z(n432) );
  XNOR2_X1 U361 ( .A(n300), .B(n432), .ZN(n301) );
  XOR2_X1 U362 ( .A(n302), .B(n301), .Z(n304) );
  XOR2_X1 U363 ( .A(G15GAT), .B(G127GAT), .Z(n328) );
  XNOR2_X1 U364 ( .A(n382), .B(n328), .ZN(n303) );
  XNOR2_X1 U365 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U366 ( .A(n307), .B(n305), .ZN(n479) );
  XOR2_X1 U367 ( .A(G92GAT), .B(G64GAT), .Z(n366) );
  XOR2_X1 U368 ( .A(n308), .B(KEYINPUT95), .Z(n316) );
  XOR2_X1 U369 ( .A(G211GAT), .B(KEYINPUT21), .Z(n310) );
  XNOR2_X1 U370 ( .A(G197GAT), .B(G218GAT), .ZN(n309) );
  XNOR2_X1 U371 ( .A(n310), .B(n309), .ZN(n446) );
  XNOR2_X1 U372 ( .A(n446), .B(KEYINPUT94), .ZN(n314) );
  XNOR2_X1 U373 ( .A(G204GAT), .B(KEYINPUT96), .ZN(n312) );
  XOR2_X1 U374 ( .A(G36GAT), .B(G8GAT), .Z(n339) );
  INV_X1 U375 ( .A(n339), .ZN(n311) );
  XNOR2_X1 U376 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U377 ( .A(G211GAT), .B(G155GAT), .Z(n318) );
  XNOR2_X1 U378 ( .A(G22GAT), .B(G78GAT), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n332) );
  XOR2_X1 U380 ( .A(G57GAT), .B(KEYINPUT13), .Z(n357) );
  XOR2_X1 U381 ( .A(KEYINPUT14), .B(n357), .Z(n320) );
  NAND2_X1 U382 ( .A1(G231GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U384 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n322) );
  XNOR2_X1 U385 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n321) );
  XNOR2_X1 U386 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U387 ( .A(n324), .B(n323), .Z(n330) );
  XOR2_X1 U388 ( .A(G64GAT), .B(G71GAT), .Z(n326) );
  XNOR2_X1 U389 ( .A(G1GAT), .B(G183GAT), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U391 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U392 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n332), .B(n331), .ZN(n586) );
  XOR2_X1 U394 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n371) );
  XOR2_X1 U395 ( .A(KEYINPUT69), .B(G1GAT), .Z(n334) );
  XNOR2_X1 U396 ( .A(G169GAT), .B(G113GAT), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U398 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n336) );
  XNOR2_X1 U399 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n338), .B(n337), .ZN(n350) );
  XOR2_X1 U402 ( .A(G15GAT), .B(G197GAT), .Z(n341) );
  XOR2_X1 U403 ( .A(G141GAT), .B(G22GAT), .Z(n443) );
  XNOR2_X1 U404 ( .A(n443), .B(n339), .ZN(n340) );
  XNOR2_X1 U405 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U406 ( .A(n342), .B(G50GAT), .Z(n348) );
  XNOR2_X1 U407 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n343), .B(KEYINPUT7), .ZN(n393) );
  XOR2_X1 U409 ( .A(n393), .B(KEYINPUT30), .Z(n345) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U411 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n346), .B(G43GAT), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X2 U414 ( .A(n350), .B(n349), .ZN(n578) );
  XOR2_X1 U415 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n356) );
  XOR2_X1 U416 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n352) );
  XNOR2_X1 U417 ( .A(G176GAT), .B(KEYINPUT75), .ZN(n351) );
  XNOR2_X1 U418 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U420 ( .A(n356), .B(n355), .Z(n361) );
  XOR2_X1 U421 ( .A(n357), .B(n378), .Z(n359) );
  NAND2_X1 U422 ( .A1(G230GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U423 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U424 ( .A(n361), .B(n360), .ZN(n368) );
  XNOR2_X1 U425 ( .A(G148GAT), .B(KEYINPUT71), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n362), .B(KEYINPUT72), .ZN(n363) );
  XOR2_X1 U427 ( .A(n363), .B(G204GAT), .Z(n365) );
  XNOR2_X1 U428 ( .A(G78GAT), .B(G106GAT), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n453) );
  XNOR2_X1 U430 ( .A(n453), .B(n366), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n582) );
  NAND2_X1 U432 ( .A1(n578), .A2(n562), .ZN(n370) );
  XOR2_X1 U433 ( .A(n371), .B(n370), .Z(n372) );
  NOR2_X1 U434 ( .A1(n586), .A2(n372), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n373), .B(KEYINPUT114), .ZN(n401) );
  XOR2_X1 U436 ( .A(KEYINPUT79), .B(KEYINPUT66), .Z(n375) );
  XNOR2_X1 U437 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n374) );
  XNOR2_X1 U438 ( .A(n375), .B(n374), .ZN(n399) );
  INV_X1 U439 ( .A(n378), .ZN(n376) );
  XNOR2_X1 U440 ( .A(G50GAT), .B(G162GAT), .ZN(n377) );
  INV_X1 U441 ( .A(n377), .ZN(n447) );
  NAND2_X1 U442 ( .A1(n376), .A2(n447), .ZN(n380) );
  NAND2_X1 U443 ( .A1(n378), .A2(n377), .ZN(n379) );
  NAND2_X1 U444 ( .A1(n380), .A2(n379), .ZN(n384) );
  NAND2_X1 U445 ( .A1(G232GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n384), .B(n383), .ZN(n392) );
  XOR2_X1 U447 ( .A(KEYINPUT78), .B(KEYINPUT76), .Z(n386) );
  XNOR2_X1 U448 ( .A(G99GAT), .B(G218GAT), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U450 ( .A(G92GAT), .B(G106GAT), .Z(n388) );
  XNOR2_X1 U451 ( .A(G36GAT), .B(G190GAT), .ZN(n387) );
  XNOR2_X1 U452 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U453 ( .A(n390), .B(n389), .Z(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n393), .B(KEYINPUT77), .ZN(n395) );
  INV_X1 U456 ( .A(KEYINPUT10), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n569) );
  XOR2_X1 U459 ( .A(KEYINPUT47), .B(n402), .Z(n409) );
  INV_X1 U460 ( .A(n586), .ZN(n474) );
  XNOR2_X1 U461 ( .A(n400), .B(KEYINPUT36), .ZN(n589) );
  NOR2_X1 U462 ( .A1(n474), .A2(n589), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n403), .B(KEYINPUT45), .ZN(n404) );
  NAND2_X1 U464 ( .A1(n404), .A2(n582), .ZN(n405) );
  XOR2_X1 U465 ( .A(n405), .B(KEYINPUT115), .Z(n406) );
  XNOR2_X1 U466 ( .A(n407), .B(KEYINPUT116), .ZN(n408) );
  NOR2_X1 U467 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U468 ( .A(KEYINPUT48), .B(n410), .ZN(n542) );
  NOR2_X1 U469 ( .A1(n507), .A2(n542), .ZN(n412) );
  XNOR2_X1 U470 ( .A(KEYINPUT124), .B(KEYINPUT54), .ZN(n411) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n438) );
  XNOR2_X1 U472 ( .A(KEYINPUT3), .B(KEYINPUT86), .ZN(n413) );
  XNOR2_X1 U473 ( .A(n413), .B(G155GAT), .ZN(n414) );
  XOR2_X1 U474 ( .A(n414), .B(KEYINPUT87), .Z(n416) );
  XNOR2_X1 U475 ( .A(KEYINPUT2), .B(KEYINPUT85), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n416), .B(n415), .ZN(n452) );
  XOR2_X1 U477 ( .A(KEYINPUT77), .B(G148GAT), .Z(n418) );
  XNOR2_X1 U478 ( .A(G141GAT), .B(G127GAT), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U480 ( .A(G85GAT), .B(G162GAT), .Z(n420) );
  XNOR2_X1 U481 ( .A(G29GAT), .B(G134GAT), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U483 ( .A(n422), .B(n421), .ZN(n436) );
  XOR2_X1 U484 ( .A(G57GAT), .B(KEYINPUT1), .Z(n424) );
  XNOR2_X1 U485 ( .A(G1GAT), .B(G120GAT), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U487 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n426) );
  XNOR2_X1 U488 ( .A(KEYINPUT92), .B(KEYINPUT6), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U490 ( .A(n428), .B(n427), .Z(n434) );
  XOR2_X1 U491 ( .A(KEYINPUT93), .B(KEYINPUT4), .Z(n430) );
  NAND2_X1 U492 ( .A1(G225GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n452), .B(n437), .ZN(n504) );
  NAND2_X1 U498 ( .A1(n438), .A2(n504), .ZN(n439) );
  XOR2_X1 U499 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n441) );
  XNOR2_X1 U500 ( .A(KEYINPUT90), .B(KEYINPUT88), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U502 ( .A(n442), .B(KEYINPUT24), .Z(n445) );
  XNOR2_X1 U503 ( .A(n443), .B(KEYINPUT89), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n451) );
  XOR2_X1 U505 ( .A(n447), .B(n446), .Z(n449) );
  NAND2_X1 U506 ( .A1(G228GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U508 ( .A(n451), .B(n450), .Z(n455) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(n466) );
  NAND2_X1 U511 ( .A1(n577), .A2(n466), .ZN(n457) );
  INV_X1 U512 ( .A(KEYINPUT55), .ZN(n456) );
  NOR2_X1 U513 ( .A1(n479), .A2(n458), .ZN(n573) );
  NAND2_X1 U514 ( .A1(n573), .A2(n562), .ZN(n461) );
  XOR2_X1 U515 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n459) );
  XNOR2_X1 U516 ( .A(n459), .B(G176GAT), .ZN(n460) );
  XNOR2_X1 U517 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  XNOR2_X1 U518 ( .A(n479), .B(KEYINPUT84), .ZN(n462) );
  XOR2_X1 U519 ( .A(n466), .B(KEYINPUT28), .Z(n536) );
  INV_X1 U520 ( .A(n504), .ZN(n530) );
  XOR2_X1 U521 ( .A(n507), .B(KEYINPUT27), .Z(n468) );
  NAND2_X1 U522 ( .A1(n530), .A2(n468), .ZN(n558) );
  NOR2_X1 U523 ( .A1(n536), .A2(n558), .ZN(n543) );
  NAND2_X1 U524 ( .A1(n462), .A2(n543), .ZN(n473) );
  INV_X1 U525 ( .A(n479), .ZN(n544) );
  INV_X1 U526 ( .A(n507), .ZN(n533) );
  NAND2_X1 U527 ( .A1(n544), .A2(n533), .ZN(n463) );
  NAND2_X1 U528 ( .A1(n466), .A2(n463), .ZN(n465) );
  NOR2_X1 U529 ( .A1(n544), .A2(n466), .ZN(n467) );
  XNOR2_X1 U530 ( .A(KEYINPUT26), .B(n467), .ZN(n576) );
  NAND2_X1 U531 ( .A1(n576), .A2(n468), .ZN(n469) );
  NAND2_X1 U532 ( .A1(n471), .A2(n504), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n473), .A2(n472), .ZN(n489) );
  NAND2_X1 U534 ( .A1(n474), .A2(n489), .ZN(n475) );
  XOR2_X1 U535 ( .A(KEYINPUT101), .B(n475), .Z(n476) );
  XNOR2_X1 U536 ( .A(KEYINPUT37), .B(n477), .ZN(n529) );
  NAND2_X1 U537 ( .A1(n578), .A2(n582), .ZN(n492) );
  NOR2_X1 U538 ( .A1(n529), .A2(n492), .ZN(n478) );
  XOR2_X1 U539 ( .A(KEYINPUT38), .B(n478), .Z(n510) );
  NOR2_X1 U540 ( .A1(n510), .A2(n479), .ZN(n482) );
  NAND2_X1 U541 ( .A1(n569), .A2(n573), .ZN(n484) );
  NAND2_X1 U542 ( .A1(n586), .A2(n573), .ZN(n486) );
  XNOR2_X1 U543 ( .A(G183GAT), .B(KEYINPUT126), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(G1350GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n494) );
  NAND2_X1 U546 ( .A1(n586), .A2(n400), .ZN(n487) );
  XNOR2_X1 U547 ( .A(n487), .B(KEYINPUT81), .ZN(n488) );
  XNOR2_X1 U548 ( .A(n488), .B(KEYINPUT16), .ZN(n490) );
  NAND2_X1 U549 ( .A1(n490), .A2(n489), .ZN(n491) );
  XOR2_X1 U550 ( .A(KEYINPUT97), .B(n491), .Z(n514) );
  NOR2_X1 U551 ( .A1(n492), .A2(n514), .ZN(n499) );
  NAND2_X1 U552 ( .A1(n499), .A2(n530), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U554 ( .A(G1GAT), .B(n495), .Z(G1324GAT) );
  NAND2_X1 U555 ( .A1(n533), .A2(n499), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n496), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U557 ( .A(G15GAT), .B(KEYINPUT35), .Z(n498) );
  NAND2_X1 U558 ( .A1(n499), .A2(n544), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(G1326GAT) );
  XOR2_X1 U560 ( .A(G22GAT), .B(KEYINPUT99), .Z(n501) );
  NAND2_X1 U561 ( .A1(n499), .A2(n536), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n501), .B(n500), .ZN(G1327GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT100), .B(KEYINPUT39), .Z(n503) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT102), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(n506) );
  NOR2_X1 U566 ( .A1(n510), .A2(n504), .ZN(n505) );
  XOR2_X1 U567 ( .A(n506), .B(n505), .Z(G1328GAT) );
  NOR2_X1 U568 ( .A1(n507), .A2(n510), .ZN(n508) );
  XOR2_X1 U569 ( .A(G36GAT), .B(n508), .Z(G1329GAT) );
  INV_X1 U570 ( .A(n536), .ZN(n509) );
  NOR2_X1 U571 ( .A1(n510), .A2(n509), .ZN(n512) );
  XNOR2_X1 U572 ( .A(G50GAT), .B(KEYINPUT103), .ZN(n511) );
  XNOR2_X1 U573 ( .A(n512), .B(n511), .ZN(G1331GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n516) );
  INV_X1 U575 ( .A(n578), .ZN(n513) );
  NAND2_X1 U576 ( .A1(n562), .A2(n513), .ZN(n528) );
  NOR2_X1 U577 ( .A1(n528), .A2(n514), .ZN(n524) );
  NAND2_X1 U578 ( .A1(n524), .A2(n530), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(n518) );
  XOR2_X1 U580 ( .A(G57GAT), .B(KEYINPUT42), .Z(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U582 ( .A(KEYINPUT104), .B(n519), .Z(G1332GAT) );
  XOR2_X1 U583 ( .A(G64GAT), .B(KEYINPUT107), .Z(n521) );
  NAND2_X1 U584 ( .A1(n524), .A2(n533), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(G1333GAT) );
  NAND2_X1 U586 ( .A1(n524), .A2(n544), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT108), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G71GAT), .B(n523), .ZN(G1334GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n526) );
  NAND2_X1 U590 ( .A1(n524), .A2(n536), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U592 ( .A(G78GAT), .B(n527), .Z(G1335GAT) );
  XNOR2_X1 U593 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n532) );
  NOR2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n530), .A2(n537), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(G1336GAT) );
  NAND2_X1 U597 ( .A1(n533), .A2(n537), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n544), .ZN(n535) );
  XNOR2_X1 U600 ( .A(n535), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(KEYINPUT111), .ZN(n541) );
  XOR2_X1 U602 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n539) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1339GAT) );
  NAND2_X1 U606 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U607 ( .A1(n542), .A2(n545), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n553), .A2(n578), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n546), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .Z(n548) );
  NAND2_X1 U611 ( .A1(n553), .A2(n562), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(G1341GAT) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n552) );
  XOR2_X1 U614 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n550) );
  NAND2_X1 U615 ( .A1(n553), .A2(n586), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U619 ( .A1(n553), .A2(n569), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  INV_X1 U621 ( .A(n542), .ZN(n556) );
  NAND2_X1 U622 ( .A1(n556), .A2(n576), .ZN(n557) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(n570) );
  NAND2_X1 U624 ( .A1(n578), .A2(n570), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G141GAT), .B(n559), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT121), .B(KEYINPUT120), .Z(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n566) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n564) );
  NAND2_X1 U630 ( .A1(n562), .A2(n570), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n586), .A2(n570), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT122), .ZN(n568) );
  XNOR2_X1 U635 ( .A(G155GAT), .B(n568), .ZN(G1346GAT) );
  XOR2_X1 U636 ( .A(G162GAT), .B(KEYINPUT123), .Z(n572) );
  NAND2_X1 U637 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(G1347GAT) );
  XOR2_X1 U639 ( .A(G169GAT), .B(KEYINPUT125), .Z(n575) );
  NAND2_X1 U640 ( .A1(n573), .A2(n578), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1348GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n588) );
  INV_X1 U644 ( .A(n588), .ZN(n585) );
  NAND2_X1 U645 ( .A1(n585), .A2(n578), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  OR2_X1 U649 ( .A1(n588), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

