//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1264, new_n1265, new_n1266,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n202), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n209), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  OR3_X1    g0019(.A1(new_n209), .A2(KEYINPUT64), .A3(G13), .ZN(new_n220));
  OAI21_X1  g0020(.A(KEYINPUT64), .B1(new_n209), .B2(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n203), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n219), .B(new_n224), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G50), .B(G68), .Z(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND2_X1  g0045(.A1(new_n202), .A2(G20), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n226), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G77), .ZN(new_n248));
  INV_X1    g0048(.A(G50), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n226), .A2(new_n250), .ZN(new_n251));
  OAI221_X1 g0051(.A(new_n246), .B1(new_n247), .B2(new_n248), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n225), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT11), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n252), .A2(KEYINPUT11), .A3(new_n254), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT69), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n202), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT12), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n257), .A2(KEYINPUT69), .A3(new_n258), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT66), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(new_n264), .B2(new_n254), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n263), .A2(KEYINPUT66), .A3(new_n225), .A4(new_n253), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n262), .A2(G20), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G68), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n261), .A2(new_n266), .A3(new_n267), .A4(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G169), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n275), .A2(KEYINPUT70), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT13), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(G1), .A2(G13), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n262), .A2(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G274), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n284), .B1(new_n281), .B2(new_n282), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n283), .A2(G238), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G226), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n291), .A2(G232), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n289), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G97), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n281), .A2(new_n282), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n277), .B(new_n288), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(new_n294), .B2(new_n295), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n285), .A2(new_n287), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n286), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n211), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT13), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n276), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT14), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n298), .A2(new_n303), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n304), .A2(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI211_X1 g0108(.A(KEYINPUT14), .B(new_n276), .C1(new_n298), .C2(new_n303), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n274), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n261), .A2(new_n266), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n298), .A2(new_n303), .A3(G190), .ZN(new_n312));
  AND2_X1   g0112(.A1(new_n267), .A2(new_n273), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n306), .A2(G200), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(G20), .A2(G77), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT15), .B(G87), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT8), .B(G58), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n316), .B1(new_n317), .B2(new_n247), .C1(new_n251), .C2(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n319), .A2(new_n254), .B1(new_n248), .B2(new_n264), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n272), .A2(G77), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n297), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n289), .A2(G232), .A3(new_n291), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n206), .B2(new_n289), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G33), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n329), .A2(new_n211), .A3(new_n291), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n323), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n283), .A2(G244), .B1(new_n285), .B2(new_n287), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n322), .B1(new_n333), .B2(G190), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n331), .A2(new_n332), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G200), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n335), .A2(new_n275), .B1(new_n320), .B2(new_n321), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n307), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n334), .A2(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n310), .A2(new_n315), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G200), .ZN(new_n341));
  NOR2_X1   g0141(.A1(G222), .A2(G1698), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n291), .A2(G223), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n289), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(new_n323), .C1(G77), .C2(new_n289), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n283), .A2(G226), .B1(new_n285), .B2(new_n287), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n341), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n345), .A2(new_n346), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n347), .B1(G190), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT10), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g0151(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n352));
  NOR2_X1   g0152(.A1(G20), .A2(G33), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G150), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n352), .B(new_n354), .C1(new_n247), .C2(new_n318), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n254), .B1(new_n249), .B2(new_n264), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT9), .ZN(new_n357));
  INV_X1    g0157(.A(new_n254), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(KEYINPUT65), .A3(new_n263), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT65), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n264), .B2(new_n254), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n359), .A2(new_n361), .A3(G50), .A4(new_n271), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n356), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n357), .B1(new_n356), .B2(new_n362), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n364), .A2(new_n365), .A3(KEYINPUT67), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT67), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n356), .A2(new_n362), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT9), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n367), .B1(new_n369), .B2(new_n363), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n351), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n363), .ZN(new_n373));
  AOI211_X1 g0173(.A(new_n372), .B(new_n350), .C1(new_n373), .C2(new_n349), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n349), .B1(new_n364), .B2(new_n365), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT68), .B1(new_n375), .B2(KEYINPUT10), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n371), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n348), .A2(G169), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n348), .A2(new_n307), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n368), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n340), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT17), .ZN(new_n382));
  INV_X1    g0182(.A(new_n318), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n264), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n359), .A2(new_n361), .A3(new_n271), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n384), .B1(new_n385), .B2(new_n383), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  OR2_X1    g0187(.A1(G223), .A2(G1698), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n290), .A2(G1698), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n327), .A2(new_n388), .A3(new_n328), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G87), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n323), .ZN(new_n393));
  INV_X1    g0193(.A(G190), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n283), .A2(G232), .B1(new_n285), .B2(new_n287), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n297), .A2(G232), .A3(new_n286), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n300), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n297), .B1(new_n390), .B2(new_n391), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n341), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n327), .A2(new_n328), .A3(KEYINPUT73), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(G20), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n327), .B2(KEYINPUT73), .ZN(new_n405));
  AOI21_X1  g0205(.A(G20), .B1(new_n327), .B2(new_n328), .ZN(new_n406));
  XOR2_X1   g0206(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n407));
  OAI22_X1  g0207(.A1(new_n402), .A2(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G68), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT72), .ZN(new_n410));
  INV_X1    g0210(.A(G159), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n410), .B1(new_n251), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n353), .A2(KEYINPUT72), .A3(G159), .ZN(new_n413));
  XNOR2_X1  g0213(.A(G58), .B(G68), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n412), .A2(new_n413), .B1(new_n414), .B2(G20), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT16), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n406), .B2(new_n403), .ZN(new_n417));
  XNOR2_X1  g0217(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n329), .A2(new_n418), .A3(new_n226), .ZN(new_n419));
  OAI211_X1 g0219(.A(KEYINPUT16), .B(new_n415), .C1(new_n417), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n254), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n387), .B(new_n401), .C1(new_n416), .C2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT74), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(G58), .A2(G68), .ZN(new_n425));
  NOR2_X1   g0225(.A1(G58), .A2(G68), .ZN(new_n426));
  OAI21_X1  g0226(.A(G20), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n413), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT72), .B1(new_n353), .B2(G159), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n430), .B1(new_n408), .B2(G68), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n254), .B(new_n420), .C1(new_n431), .C2(KEYINPUT16), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n432), .A2(KEYINPUT74), .A3(new_n387), .A4(new_n401), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n382), .B1(new_n424), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n422), .A2(new_n382), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n432), .A2(new_n387), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n393), .A2(new_n395), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(G169), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n439), .B2(new_n307), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT18), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n438), .A2(new_n444), .A3(new_n441), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n381), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(G116), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT76), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n250), .B2(G1), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n262), .A2(KEYINPUT76), .A3(G33), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n269), .A2(new_n270), .A3(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n262), .A2(new_n450), .A3(G13), .A4(G20), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT83), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n450), .A2(G20), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n254), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT84), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n254), .A2(KEYINPUT84), .A3(new_n459), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(G20), .B1(G33), .B2(G283), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT75), .B(G97), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(G33), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT20), .B1(new_n464), .B2(new_n467), .ZN(new_n468));
  AOI221_X4 g0268(.A(new_n461), .B1(new_n450), .B2(G20), .C1(new_n253), .C2(new_n225), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT84), .B1(new_n254), .B2(new_n459), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n467), .B(KEYINPUT20), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n458), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n262), .B(G45), .C1(new_n278), .C2(KEYINPUT5), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT78), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G41), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n478), .A2(KEYINPUT78), .A3(new_n262), .A4(G45), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n477), .A2(G41), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n476), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G270), .A3(new_n297), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n326), .A2(G33), .ZN(new_n485));
  OAI21_X1  g0285(.A(G303), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n327), .A2(new_n328), .A3(G264), .A4(G1698), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n327), .A2(new_n328), .A3(G257), .A4(new_n291), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n323), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n480), .B1(new_n474), .B2(new_n475), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(new_n285), .A3(new_n479), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n483), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(KEYINPUT82), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT82), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n483), .A2(new_n490), .A3(new_n495), .A4(new_n492), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n473), .B1(new_n497), .B2(G190), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n341), .B2(new_n497), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n493), .A2(new_n307), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n473), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  AND4_X1   g0302(.A1(G169), .A2(new_n473), .A3(new_n494), .A4(new_n496), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(KEYINPUT21), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n473), .A2(new_n494), .A3(G169), .A4(new_n496), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT85), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT21), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n499), .B(new_n504), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n211), .A2(new_n291), .ZN(new_n512));
  INV_X1    g0312(.A(G244), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G1698), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n327), .A2(new_n512), .A3(new_n328), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G116), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n297), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n262), .A2(new_n284), .A3(G45), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n213), .B1(new_n279), .B2(G1), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n297), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT79), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT79), .ZN(new_n523));
  NOR2_X1   g0323(.A1(G238), .A2(G1698), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n524), .B1(new_n513), .B2(G1698), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n525), .A2(new_n289), .B1(G33), .B2(G116), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n523), .B(new_n520), .C1(new_n526), .C2(new_n297), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n522), .A2(new_n527), .A3(new_n307), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT80), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n522), .A2(new_n527), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n275), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n522), .A2(new_n527), .A3(KEYINPUT80), .A4(new_n307), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n327), .A2(new_n328), .A3(new_n226), .A4(G68), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n205), .A2(KEYINPUT75), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT75), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G97), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n247), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n534), .B1(new_n538), .B2(KEYINPUT19), .ZN(new_n539));
  NAND3_X1  g0339(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n540), .A2(new_n226), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G87), .A2(G107), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(new_n466), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n254), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n317), .A2(new_n264), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n264), .A2(new_n254), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n452), .A2(new_n453), .ZN(new_n547));
  INV_X1    g0347(.A(new_n317), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n544), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n530), .A2(new_n532), .A3(new_n533), .A4(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n546), .A2(G87), .A3(new_n547), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT81), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n546), .A2(KEYINPUT81), .A3(G87), .A4(new_n547), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n556), .A2(new_n544), .A3(new_n545), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n531), .A2(G200), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n522), .A2(new_n527), .A3(G190), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n551), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n327), .A2(new_n328), .A3(G244), .A4(new_n291), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT4), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G250), .A2(G1698), .ZN(new_n565));
  NAND2_X1  g0365(.A1(KEYINPUT4), .A2(G244), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n565), .B1(new_n566), .B2(G1698), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n289), .A2(new_n567), .B1(G33), .B2(G283), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n323), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n482), .A2(G257), .A3(new_n297), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n492), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(new_n394), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n226), .B1(new_n484), .B2(new_n485), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n418), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT73), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n484), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n577), .B(new_n404), .C1(new_n329), .C2(new_n576), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n206), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(new_n535), .B2(new_n537), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G97), .A2(G107), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT6), .B1(new_n207), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(G20), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n353), .A2(G77), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n254), .B1(new_n579), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n264), .A2(new_n205), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n546), .A2(new_n547), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(new_n205), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n573), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n323), .B1(new_n491), .B2(new_n479), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n476), .A2(new_n479), .A3(new_n481), .ZN(new_n595));
  AOI22_X1  g0395(.A1(G257), .A2(new_n594), .B1(new_n595), .B2(new_n285), .ZN(new_n596));
  AOI21_X1  g0396(.A(KEYINPUT77), .B1(new_n569), .B2(new_n323), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT77), .ZN(new_n598));
  AOI211_X1 g0398(.A(new_n598), .B(new_n297), .C1(new_n564), .C2(new_n568), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n596), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G200), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n587), .A2(new_n591), .B1(new_n572), .B2(new_n275), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n596), .B(new_n307), .C1(new_n597), .C2(new_n599), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n593), .A2(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g0404(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n327), .A2(new_n328), .A3(new_n226), .A4(G87), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n289), .A2(new_n605), .A3(new_n226), .A4(G87), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n516), .A2(G20), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT23), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n226), .B2(G107), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT24), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT24), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n608), .A2(new_n609), .A3(new_n617), .A4(new_n614), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n358), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n263), .A2(G107), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT25), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n206), .B2(new_n589), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n327), .A2(new_n328), .A3(G257), .A4(G1698), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n327), .A2(new_n328), .A3(G250), .A4(new_n291), .ZN(new_n626));
  AND2_X1   g0426(.A1(KEYINPUT87), .A2(G294), .ZN(new_n627));
  NOR2_X1   g0427(.A1(KEYINPUT87), .A2(G294), .ZN(new_n628));
  OAI21_X1  g0428(.A(G33), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n625), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n297), .B1(new_n630), .B2(KEYINPUT88), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT88), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n625), .A2(new_n626), .A3(new_n632), .A4(new_n629), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n631), .A2(new_n633), .B1(G264), .B2(new_n594), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n492), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n275), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n307), .A3(new_n492), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n624), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(G200), .B1(new_n634), .B2(new_n492), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n630), .A2(KEYINPUT88), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n323), .A3(new_n633), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n594), .A2(G264), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n394), .A2(new_n641), .A3(new_n492), .A4(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n623), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n561), .A2(new_n604), .A3(new_n638), .A4(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n449), .A2(new_n511), .A3(new_n645), .ZN(G372));
  OAI211_X1 g0446(.A(new_n504), .B(new_n638), .C1(new_n509), .C2(new_n510), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT19), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n466), .B2(new_n247), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n466), .A2(new_n542), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n534), .B(new_n649), .C1(new_n650), .C2(new_n541), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n651), .A2(new_n254), .B1(new_n264), .B2(new_n317), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n520), .B1(new_n526), .B2(new_n297), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G200), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n559), .A2(new_n652), .A3(new_n556), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n275), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n528), .A2(new_n550), .A3(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n408), .A2(G107), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n659), .A2(new_n584), .A3(new_n585), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n590), .B1(new_n660), .B2(new_n254), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n596), .A2(G190), .A3(new_n570), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n571), .A2(new_n492), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n570), .A2(new_n598), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n569), .A2(KEYINPUT77), .A3(new_n323), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n661), .B(new_n662), .C1(new_n666), .C2(new_n341), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n572), .A2(new_n275), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n603), .A2(new_n592), .A3(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n644), .A2(new_n658), .A3(new_n667), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT89), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT89), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n604), .A2(new_n672), .A3(new_n644), .A4(new_n658), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n647), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n602), .A2(new_n603), .A3(new_n655), .A4(new_n657), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n657), .B1(new_n675), .B2(KEYINPUT26), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n603), .A2(new_n592), .A3(new_n668), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n561), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n676), .B1(new_n678), .B2(KEYINPUT26), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n448), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT90), .ZN(new_n682));
  INV_X1    g0482(.A(new_n380), .ZN(new_n683));
  INV_X1    g0483(.A(new_n315), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n337), .A2(new_n338), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n310), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n437), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n446), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n683), .B1(new_n688), .B2(new_n377), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n682), .A2(new_n689), .ZN(G369));
  OAI21_X1  g0490(.A(new_n501), .B1(new_n505), .B2(new_n507), .ZN(new_n691));
  INV_X1    g0491(.A(new_n510), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(new_n508), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n262), .A2(new_n226), .A3(G13), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  INV_X1    g0496(.A(G213), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G343), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n473), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n693), .A2(new_n499), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n693), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT91), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n638), .A2(new_n699), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT92), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n638), .B(new_n644), .C1(new_n623), .C2(new_n699), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n705), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n693), .A2(new_n700), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n638), .B2(new_n700), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n711), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n222), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n650), .A2(new_n450), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n717), .A2(new_n262), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n229), .B2(new_n717), .ZN(new_n720));
  XOR2_X1   g0520(.A(new_n720), .B(KEYINPUT28), .Z(new_n721));
  AOI21_X1  g0521(.A(new_n700), .B1(new_n674), .B2(new_n679), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT26), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n677), .A2(new_n725), .A3(new_n560), .A4(new_n551), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n655), .A2(new_n657), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT26), .B1(new_n727), .B2(new_n669), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n726), .A2(new_n657), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n670), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n647), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n700), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n723), .ZN(new_n733));
  INV_X1    g0533(.A(G330), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n570), .A2(new_n492), .A3(new_n571), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n522), .A2(new_n527), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n500), .A2(new_n735), .A3(new_n634), .A4(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n572), .A2(new_n531), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n740), .A2(KEYINPUT30), .A3(new_n500), .A4(new_n634), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n635), .A2(new_n600), .A3(new_n307), .A4(new_n653), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n739), .B(new_n741), .C1(new_n497), .C2(new_n742), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT31), .B1(new_n743), .B2(new_n700), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AND4_X1   g0546(.A1(new_n638), .A2(new_n561), .A3(new_n604), .A4(new_n644), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n747), .A2(new_n693), .A3(new_n499), .A4(new_n699), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n734), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n724), .A2(new_n733), .A3(new_n749), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT93), .Z(new_n751));
  OAI21_X1  g0551(.A(new_n721), .B1(new_n751), .B2(G1), .ZN(G364));
  INV_X1    g0552(.A(new_n717), .ZN(new_n753));
  INV_X1    g0553(.A(G13), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n262), .B1(new_n755), .B2(G45), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n758));
  XOR2_X1   g0558(.A(new_n758), .B(KEYINPUT94), .Z(new_n759));
  OR2_X1    g0559(.A1(new_n703), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n759), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n225), .B1(G20), .B2(new_n275), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT95), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n716), .A2(new_n289), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n279), .B2(new_n229), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(new_n241), .B2(new_n279), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n716), .A2(new_n329), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n769), .A2(G355), .B1(new_n450), .B2(new_n716), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n764), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n394), .ZN(new_n773));
  AND2_X1   g0573(.A1(new_n773), .A2(G326), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n226), .A2(new_n394), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n341), .A2(G179), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n289), .B(new_n774), .C1(G303), .C2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n307), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n226), .A2(G190), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G179), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G322), .A2(new_n782), .B1(new_n786), .B2(G329), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n780), .A2(new_n783), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n783), .A2(new_n776), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G311), .A2(new_n789), .B1(new_n791), .B2(G283), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n226), .B1(new_n784), .B2(G190), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n627), .A2(new_n628), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n772), .A2(G190), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n794), .A2(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n779), .A2(new_n787), .A3(new_n792), .A4(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G58), .A2(new_n782), .B1(new_n789), .B2(G77), .ZN(new_n801));
  INV_X1    g0601(.A(new_n773), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n249), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT96), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n778), .A2(G87), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n289), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G107), .B2(new_n791), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n793), .A2(new_n205), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(new_n797), .B2(G68), .ZN(new_n809));
  OAI21_X1  g0609(.A(KEYINPUT32), .B1(new_n785), .B2(new_n411), .ZN(new_n810));
  OR3_X1    g0610(.A1(new_n785), .A2(KEYINPUT32), .A3(new_n411), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n807), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n800), .B1(new_n804), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n771), .B1(new_n813), .B2(new_n762), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n757), .B1(new_n760), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n705), .B1(G330), .B2(new_n703), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(new_n816), .B2(new_n757), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT97), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  NAND2_X1  g0619(.A1(new_n339), .A2(new_n699), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n820), .B1(new_n674), .B2(new_n679), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n685), .A2(new_n700), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n334), .A2(new_n336), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n322), .A2(new_n700), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n823), .B1(new_n826), .B2(new_n685), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n822), .B1(new_n722), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n749), .ZN(new_n829));
  OR2_X1    g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n757), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n828), .B2(new_n829), .ZN(new_n832));
  INV_X1    g0632(.A(new_n827), .ZN(new_n833));
  NOR2_X1   g0633(.A1(G13), .A2(G33), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n762), .A2(new_n834), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n757), .B1(new_n248), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT98), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n289), .B(new_n808), .C1(G294), .C2(new_n782), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G116), .A2(new_n789), .B1(new_n786), .B2(G311), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G107), .A2(new_n778), .B1(new_n791), .B2(G87), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G283), .A2(new_n797), .B1(new_n773), .B2(G303), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(KEYINPUT99), .B(G143), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n782), .A2(new_n844), .B1(new_n789), .B2(G159), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  INV_X1    g0646(.A(G150), .ZN(new_n847));
  INV_X1    g0647(.A(new_n797), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n845), .B1(new_n802), .B2(new_n846), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT34), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n289), .B1(new_n777), .B2(new_n249), .ZN(new_n852));
  INV_X1    g0652(.A(G132), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n790), .A2(new_n202), .B1(new_n785), .B2(new_n853), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n852), .B(new_n854), .C1(G58), .C2(new_n794), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n849), .A2(new_n850), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n843), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n838), .B1(new_n858), .B2(new_n762), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n830), .A2(new_n832), .B1(new_n835), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G384));
  NAND2_X1  g0661(.A1(new_n227), .A2(G116), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n581), .A2(new_n583), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n863), .B2(KEYINPUT35), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(KEYINPUT35), .B2(new_n863), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT36), .ZN(new_n866));
  OAI21_X1  g0666(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n228), .A2(new_n867), .B1(G50), .B2(new_n202), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(G1), .A3(new_n754), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT100), .Z(new_n871));
  NAND2_X1  g0671(.A1(new_n274), .A2(new_n700), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n310), .A2(new_n315), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n872), .B1(new_n310), .B2(new_n315), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n823), .B(KEYINPUT101), .Z(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n821), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT102), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n202), .B1(new_n574), .B2(KEYINPUT7), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n406), .A2(new_n418), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n430), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n883), .A2(KEYINPUT16), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n387), .B1(new_n884), .B2(new_n421), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n698), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n437), .B2(new_n446), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n698), .B(KEYINPUT103), .Z(new_n889));
  NAND2_X1  g0689(.A1(new_n438), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n442), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n424), .A2(new_n433), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n885), .B1(new_n441), .B2(new_n698), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n424), .A3(new_n433), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n892), .A2(new_n894), .B1(new_n896), .B2(KEYINPUT37), .ZN(new_n897));
  OR3_X1    g0697(.A1(new_n887), .A2(new_n888), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n888), .B1(new_n887), .B2(new_n897), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI211_X1 g0700(.A(KEYINPUT102), .B(new_n876), .C1(new_n821), .C2(new_n877), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n880), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n446), .A2(new_n889), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n902), .A2(KEYINPUT104), .A3(new_n904), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n310), .A2(new_n700), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT39), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n887), .A2(new_n897), .A3(new_n888), .ZN(new_n909));
  INV_X1    g0709(.A(new_n890), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n443), .A2(new_n910), .A3(new_n445), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n358), .B1(new_n883), .B2(KEYINPUT16), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT16), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n202), .B1(new_n575), .B2(new_n578), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n913), .B1(new_n914), .B2(new_n430), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n386), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT74), .B1(new_n916), .B2(new_n401), .ZN(new_n917));
  INV_X1    g0717(.A(new_n433), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT17), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(KEYINPUT105), .A3(new_n435), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT105), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n434), .B2(new_n436), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n911), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n422), .B1(new_n910), .B2(new_n442), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT37), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT38), .B1(new_n892), .B2(new_n894), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n909), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n907), .B(new_n908), .C1(new_n927), .C2(KEYINPUT39), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n905), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT104), .B1(new_n902), .B2(new_n904), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT106), .ZN(new_n932));
  INV_X1    g0732(.A(new_n928), .ZN(new_n933));
  AOI22_X1  g0733(.A1(new_n878), .A2(new_n879), .B1(new_n898), .B2(new_n899), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n903), .B1(new_n934), .B2(new_n901), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n935), .B2(KEYINPUT104), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n902), .A2(new_n904), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT104), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n932), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n931), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n448), .B1(new_n724), .B2(new_n733), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n689), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n941), .B(new_n943), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n511), .A2(new_n645), .A3(new_n700), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n739), .A2(new_n741), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n742), .A2(new_n497), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n700), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT31), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n827), .B(new_n876), .C1(new_n945), .C2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT40), .B1(new_n927), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(KEYINPUT40), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n900), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n449), .B1(new_n748), .B2(new_n746), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(G330), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n944), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n262), .B2(new_n755), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n944), .A2(new_n961), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n871), .B1(new_n963), .B2(new_n964), .ZN(G367));
  OAI21_X1  g0765(.A(new_n604), .B1(new_n661), .B2(new_n699), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n677), .A2(new_n700), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n711), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n557), .A2(new_n699), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n658), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n657), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n969), .B(new_n973), .Z(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n975));
  INV_X1    g0775(.A(new_n713), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n968), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(KEYINPUT42), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n669), .B1(new_n966), .B2(new_n638), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n699), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n977), .A2(KEYINPUT42), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n975), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT107), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n974), .B(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(new_n968), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n714), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT44), .Z(new_n988));
  NOR2_X1   g0788(.A1(new_n714), .A2(new_n986), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(new_n711), .Z(new_n992));
  NOR2_X1   g0792(.A1(new_n709), .A2(new_n712), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n976), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n705), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n751), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n751), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT108), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n717), .B(KEYINPUT41), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n756), .B(KEYINPUT109), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1000), .B1(new_n999), .B2(new_n1001), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n985), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n972), .A2(new_n759), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n766), .A2(new_n237), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n763), .B1(new_n222), .B2(new_n317), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n289), .B1(new_n777), .B2(new_n201), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1011), .B1(G68), .B2(new_n794), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G150), .A2(new_n782), .B1(new_n791), .B2(G77), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G50), .A2(new_n789), .B1(new_n786), .B2(G137), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n773), .A2(new_n844), .B1(new_n797), .B2(G159), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n289), .B1(new_n786), .B2(G317), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n466), .B2(new_n790), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT111), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n778), .A2(G116), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT46), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n1021), .A2(new_n1022), .B1(new_n795), .B2(new_n848), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G107), .B2(new_n794), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1020), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT110), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT110), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n773), .A2(G311), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G303), .A2(new_n782), .B1(new_n789), .B2(G283), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1016), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT47), .Z(new_n1034));
  INV_X1    g0834(.A(new_n762), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n831), .B1(new_n1009), .B2(new_n1010), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1008), .B1(new_n1036), .B2(KEYINPUT112), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(KEYINPUT112), .B2(new_n1036), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1007), .A2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT113), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(G387));
  NOR2_X1   g0841(.A1(new_n997), .A2(new_n753), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n751), .B2(new_n995), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n769), .A2(new_n718), .B1(new_n206), .B2(new_n716), .ZN(new_n1044));
  AOI211_X1 g0844(.A(G45), .B(new_n718), .C1(G68), .C2(G77), .ZN(new_n1045));
  AOI21_X1  g0845(.A(KEYINPUT50), .B1(new_n383), .B2(new_n249), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n383), .A2(KEYINPUT50), .A3(new_n249), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n765), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n234), .A2(new_n279), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1044), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n764), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n757), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n329), .B1(new_n789), .B2(G68), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n794), .A2(new_n548), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(new_n848), .C2(new_n318), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n773), .A2(G159), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT114), .Z(new_n1058));
  OAI22_X1  g0858(.A1(new_n777), .A2(new_n248), .B1(new_n785), .B2(new_n847), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n781), .A2(new_n249), .B1(new_n790), .B2(new_n205), .ZN(new_n1060));
  NOR4_X1   g0860(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(G283), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n777), .A2(new_n795), .B1(new_n793), .B2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G317), .A2(new_n782), .B1(new_n789), .B2(G303), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n797), .A2(G311), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n773), .A2(G322), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1063), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT115), .Z(new_n1071));
  OR2_X1    g0871(.A1(new_n1071), .A2(KEYINPUT49), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n289), .B1(new_n786), .B2(G326), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n450), .B2(new_n790), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1074), .B1(new_n1071), .B2(KEYINPUT49), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1061), .B1(new_n1072), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1053), .B1(new_n1076), .B2(new_n1035), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n710), .B2(new_n761), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n995), .B2(new_n1003), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1043), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT116), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1043), .A2(KEYINPUT116), .A3(new_n1079), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(G393));
  AOI21_X1  g0884(.A(new_n753), .B1(new_n992), .B2(new_n997), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n997), .B2(new_n992), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n992), .A2(new_n1003), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n763), .B1(new_n222), .B2(new_n466), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n766), .A2(new_n244), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n831), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n802), .A2(new_n847), .B1(new_n781), .B2(new_n411), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT51), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n793), .A2(new_n248), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n289), .B1(new_n790), .B2(new_n212), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1093), .B(new_n1094), .C1(G50), .C2(new_n797), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n777), .A2(new_n202), .B1(new_n788), .B2(new_n318), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n786), .B2(new_n844), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1092), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n782), .A2(G311), .B1(G317), .B2(new_n773), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT52), .Z(new_n1100));
  AOI22_X1  g0900(.A1(G283), .A2(new_n778), .B1(new_n786), .B2(G322), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1101), .A2(KEYINPUT117), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(KEYINPUT117), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n289), .B1(new_n791), .B2(G107), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(G294), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n788), .A2(new_n1106), .B1(new_n793), .B2(new_n450), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G303), .B2(new_n797), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT118), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1098), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1090), .B1(new_n1110), .B2(new_n762), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n968), .B2(new_n759), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1086), .A2(new_n1087), .A3(new_n1112), .ZN(G390));
  INV_X1    g0913(.A(new_n877), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n822), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n876), .B1(new_n749), .B2(new_n827), .ZN(new_n1116));
  OAI211_X1 g0916(.A(G330), .B(new_n827), .C1(new_n945), .C2(new_n952), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(new_n875), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1115), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n875), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n731), .A2(new_n700), .A3(new_n833), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1121), .A2(KEYINPUT119), .A3(new_n877), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT119), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n670), .B1(new_n693), .B2(new_n638), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n699), .B(new_n827), .C1(new_n1124), .C2(new_n729), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n1125), .B2(new_n1114), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1120), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT120), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n1117), .B2(new_n875), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n749), .A2(KEYINPUT120), .A3(new_n827), .A4(new_n876), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1119), .B1(new_n1127), .B2(new_n1131), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n448), .B(G330), .C1(new_n945), .C2(new_n952), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(KEYINPUT121), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT121), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n749), .A2(new_n1135), .A3(new_n448), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1137), .A2(new_n689), .A3(new_n942), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n1132), .A2(new_n1138), .A3(KEYINPUT122), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT122), .B1(new_n1132), .B2(new_n1138), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n908), .B1(new_n927), .B2(KEYINPUT39), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n878), .A2(new_n906), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(KEYINPUT119), .B1(new_n1121), .B2(new_n877), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1125), .A2(new_n1123), .A3(new_n1114), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n876), .A3(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n927), .A2(new_n907), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1144), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1142), .A2(new_n1143), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n749), .A2(new_n827), .A3(new_n876), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1141), .A2(new_n1154), .ZN(new_n1155));
  OR2_X1    g0955(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1156), .B(new_n1151), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1155), .A2(new_n717), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1154), .A2(new_n1004), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1142), .A2(new_n834), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n836), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n831), .B1(new_n383), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n777), .A2(new_n847), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT53), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(G132), .A2(new_n782), .B1(new_n786), .B2(G125), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(KEYINPUT54), .B(G143), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1164), .B(new_n1165), .C1(new_n788), .C2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n329), .B1(new_n791), .B2(G50), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G128), .A2(new_n773), .B1(new_n797), .B2(G137), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(new_n411), .C2(new_n793), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G116), .A2(new_n782), .B1(new_n786), .B2(G294), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n202), .B2(new_n790), .C1(new_n466), .C2(new_n788), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1093), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G107), .A2(new_n797), .B1(new_n773), .B2(G283), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n805), .A2(new_n1173), .A3(new_n1174), .A4(new_n329), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n1167), .A2(new_n1170), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1162), .B1(new_n1176), .B2(new_n762), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1159), .B1(new_n1160), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1158), .A2(new_n1178), .ZN(G378));
  NAND2_X1  g0979(.A1(new_n377), .A2(new_n380), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(new_n368), .A3(new_n698), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n368), .A2(new_n698), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n377), .A2(new_n380), .A3(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1181), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1184), .B1(new_n1181), .B2(new_n1183), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n957), .B2(G330), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n734), .B(new_n1187), .C1(new_n954), .C2(new_n956), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n931), .B2(new_n940), .ZN(new_n1193));
  OAI21_X1  g0993(.A(KEYINPUT106), .B1(new_n929), .B2(new_n930), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n939), .A2(new_n932), .A3(new_n928), .A4(new_n905), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n1191), .A3(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1193), .A2(new_n1003), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1187), .A2(new_n834), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n757), .B1(new_n249), .B2(new_n836), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n848), .A2(new_n853), .B1(new_n793), .B2(new_n847), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1166), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G128), .A2(new_n782), .B1(new_n778), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n846), .B2(new_n788), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1200), .B(new_n1203), .C1(G125), .C2(new_n773), .ZN(new_n1204));
  XOR2_X1   g1004(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n1205));
  OR2_X1    g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n250), .B(new_n278), .C1(new_n790), .C2(new_n411), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G124), .B2(new_n786), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n329), .A2(new_n278), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1212), .B(new_n249), .C1(G33), .C2(G41), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1212), .B1(G77), .B2(new_n778), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n201), .B2(new_n790), .C1(new_n1062), .C2(new_n785), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT123), .Z(new_n1216));
  OAI22_X1  g1016(.A1(new_n781), .A2(new_n206), .B1(new_n788), .B2(new_n317), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G68), .B2(new_n794), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G97), .A2(new_n797), .B1(new_n773), .B2(G116), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1216), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1213), .B1(new_n1221), .B2(KEYINPUT58), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1211), .B(new_n1222), .C1(KEYINPUT58), .C2(new_n1221), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1198), .B(new_n1199), .C1(new_n1035), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1197), .A2(new_n1224), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1194), .A2(new_n1191), .A3(new_n1195), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1191), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT57), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n1157), .B2(new_n1138), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n753), .B1(new_n1228), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1193), .A2(new_n1196), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT122), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1153), .A2(new_n1120), .B1(new_n822), .B2(new_n1114), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1116), .B1(new_n1146), .B2(new_n1145), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(new_n1150), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1137), .A2(new_n689), .A3(new_n942), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1233), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1132), .A2(new_n1138), .A3(KEYINPUT122), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1154), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(new_n1237), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1229), .B1(new_n1232), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1225), .B1(new_n1231), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(G375));
  NAND2_X1  g1044(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1141), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1001), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n875), .A2(new_n834), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n831), .B1(G68), .B2(new_n1161), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n329), .B1(new_n791), .B2(G58), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1201), .A2(new_n797), .B1(G132), .B2(new_n773), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1250), .B(new_n1251), .C1(new_n249), .C2(new_n793), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G159), .A2(new_n778), .B1(new_n786), .B2(G128), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n846), .B2(new_n781), .C1(new_n847), .C2(new_n788), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G97), .A2(new_n778), .B1(new_n786), .B2(G303), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n206), .B2(new_n788), .C1(new_n1062), .C2(new_n781), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n289), .B1(new_n791), .B2(G77), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G116), .A2(new_n797), .B1(new_n773), .B2(G294), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1055), .A3(new_n1258), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1252), .A2(new_n1254), .B1(new_n1256), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1249), .B1(new_n1260), .B2(new_n762), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1132), .A2(new_n1003), .B1(new_n1248), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1247), .A2(new_n1262), .ZN(G381));
  INV_X1    g1063(.A(G378), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1082), .A2(new_n818), .A3(new_n1083), .ZN(new_n1265));
  NOR4_X1   g1065(.A1(G390), .A2(new_n1265), .A3(G384), .A4(G381), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1040), .A2(new_n1264), .A3(new_n1243), .A4(new_n1266), .ZN(G407));
  NOR2_X1   g1067(.A1(new_n697), .A2(G343), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1243), .A2(new_n1264), .A3(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(G407), .A2(G213), .A3(new_n1269), .ZN(G409));
  NAND2_X1  g1070(.A1(G393), .A2(G396), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1265), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(G390), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT113), .B1(new_n1271), .B2(new_n1265), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1273), .B1(G390), .B2(new_n1274), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1007), .A2(new_n1038), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1039), .B(new_n1273), .C1(G390), .C2(new_n1274), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(KEYINPUT61), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1197), .A2(new_n1224), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1157), .A2(new_n1138), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1228), .A2(new_n1001), .A3(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(G378), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT57), .B1(new_n1228), .B2(new_n1282), .ZN(new_n1286));
  OAI21_X1  g1086(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1237), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n717), .B1(new_n1232), .B2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1281), .C1(new_n1286), .C2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT125), .B1(new_n1243), .B2(G378), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1285), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT126), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1268), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1231), .A2(new_n1242), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1298), .A2(KEYINPUT125), .A3(G378), .A4(new_n1281), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1284), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT126), .B1(new_n1300), .B2(new_n1268), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT60), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n753), .B1(new_n1245), .B2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1246), .B2(new_n1302), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1262), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1305), .B(G384), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1296), .A2(new_n1301), .A3(KEYINPUT63), .A4(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1293), .A2(new_n1295), .A3(new_n1306), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1268), .A2(G2897), .ZN(new_n1311));
  XOR2_X1   g1111(.A(new_n1306), .B(new_n1311), .Z(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1268), .B2(new_n1300), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1280), .A2(new_n1307), .A3(new_n1310), .A4(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1296), .A2(new_n1301), .ZN(new_n1315));
  AOI21_X1  g1115(.A(KEYINPUT61), .B1(new_n1315), .B2(new_n1312), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1306), .A2(KEYINPUT62), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1296), .A2(new_n1301), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT62), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1308), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1316), .A2(new_n1321), .A3(KEYINPUT127), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1279), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT127), .B1(new_n1316), .B2(new_n1321), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1314), .B1(new_n1323), .B2(new_n1324), .ZN(G405));
  OAI22_X1  g1125(.A1(new_n1291), .A2(new_n1292), .B1(G378), .B2(new_n1243), .ZN(new_n1326));
  XNOR2_X1  g1126(.A(new_n1326), .B(new_n1306), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(new_n1279), .B(new_n1327), .ZN(G402));
endmodule


