

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(n541), .A2(n536), .ZN(n548) );
  OR2_X1 U553 ( .A1(n720), .A2(n719), .ZN(n518) );
  NOR2_X1 U554 ( .A1(n678), .A2(n883), .ZN(n648) );
  AND2_X1 U555 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U556 ( .A(n666), .B(KEYINPUT29), .ZN(n667) );
  NAND2_X1 U557 ( .A1(n615), .A2(n614), .ZN(n678) );
  INV_X1 U558 ( .A(KEYINPUT102), .ZN(n697) );
  NAND2_X1 U559 ( .A1(n721), .A2(n518), .ZN(n722) );
  NOR2_X1 U560 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U561 ( .A1(n571), .A2(n523), .ZN(n783) );
  NOR2_X1 U562 ( .A1(n571), .A2(G651), .ZN(n787) );
  NOR2_X1 U563 ( .A1(n555), .A2(n554), .ZN(G160) );
  INV_X1 U564 ( .A(G651), .ZN(n523) );
  NOR2_X1 U565 ( .A1(G543), .A2(n523), .ZN(n519) );
  XOR2_X1 U566 ( .A(KEYINPUT1), .B(n519), .Z(n782) );
  NAND2_X1 U567 ( .A1(G63), .A2(n782), .ZN(n521) );
  XOR2_X1 U568 ( .A(KEYINPUT0), .B(G543), .Z(n571) );
  NAND2_X1 U569 ( .A1(G51), .A2(n787), .ZN(n520) );
  NAND2_X1 U570 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U571 ( .A(KEYINPUT6), .B(n522), .ZN(n531) );
  NAND2_X1 U572 ( .A1(n783), .A2(G76), .ZN(n524) );
  XNOR2_X1 U573 ( .A(KEYINPUT70), .B(n524), .ZN(n528) );
  XOR2_X1 U574 ( .A(KEYINPUT4), .B(KEYINPUT69), .Z(n526) );
  NOR2_X1 U575 ( .A1(G543), .A2(G651), .ZN(n786) );
  NAND2_X1 U576 ( .A1(G89), .A2(n786), .ZN(n525) );
  XNOR2_X1 U577 ( .A(n526), .B(n525), .ZN(n527) );
  NAND2_X1 U578 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U579 ( .A(n529), .B(KEYINPUT5), .Z(n530) );
  NOR2_X1 U580 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U581 ( .A(KEYINPUT7), .B(n532), .Z(n534) );
  XOR2_X1 U582 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n533) );
  XNOR2_X1 U583 ( .A(n534), .B(n533), .ZN(G168) );
  XOR2_X1 U584 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  INV_X1 U585 ( .A(G2104), .ZN(n536) );
  NOR2_X2 U586 ( .A1(G2105), .A2(n536), .ZN(n990) );
  NAND2_X1 U587 ( .A1(G102), .A2(n990), .ZN(n535) );
  XNOR2_X1 U588 ( .A(n535), .B(KEYINPUT88), .ZN(n539) );
  INV_X1 U589 ( .A(G2105), .ZN(n541) );
  NAND2_X1 U590 ( .A1(G114), .A2(n548), .ZN(n537) );
  XOR2_X1 U591 ( .A(KEYINPUT87), .B(n537), .Z(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n545) );
  NOR2_X1 U593 ( .A1(G2105), .A2(G2104), .ZN(n540) );
  XOR2_X1 U594 ( .A(KEYINPUT17), .B(n540), .Z(n991) );
  NAND2_X1 U595 ( .A1(G138), .A2(n991), .ZN(n543) );
  NOR2_X1 U596 ( .A1(G2104), .A2(n541), .ZN(n987) );
  NAND2_X1 U597 ( .A1(G126), .A2(n987), .ZN(n542) );
  NAND2_X1 U598 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U599 ( .A1(n545), .A2(n544), .ZN(G164) );
  NAND2_X1 U600 ( .A1(G101), .A2(n990), .ZN(n547) );
  XOR2_X1 U601 ( .A(KEYINPUT64), .B(KEYINPUT23), .Z(n546) );
  XNOR2_X1 U602 ( .A(n547), .B(n546), .ZN(n551) );
  NAND2_X1 U603 ( .A1(G113), .A2(n548), .ZN(n549) );
  XOR2_X1 U604 ( .A(KEYINPUT65), .B(n549), .Z(n550) );
  NAND2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U606 ( .A1(G137), .A2(n991), .ZN(n553) );
  NAND2_X1 U607 ( .A1(G125), .A2(n987), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U609 ( .A1(G64), .A2(n782), .ZN(n557) );
  NAND2_X1 U610 ( .A1(G52), .A2(n787), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n557), .A2(n556), .ZN(n562) );
  NAND2_X1 U612 ( .A1(G77), .A2(n783), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G90), .A2(n786), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U615 ( .A(KEYINPUT9), .B(n560), .Z(n561) );
  NOR2_X1 U616 ( .A1(n562), .A2(n561), .ZN(G171) );
  NAND2_X1 U617 ( .A1(G62), .A2(n782), .ZN(n564) );
  NAND2_X1 U618 ( .A1(G75), .A2(n783), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U620 ( .A1(G88), .A2(n786), .ZN(n566) );
  NAND2_X1 U621 ( .A1(G50), .A2(n787), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U623 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U624 ( .A(KEYINPUT82), .B(n569), .Z(G303) );
  NAND2_X1 U625 ( .A1(G74), .A2(G651), .ZN(n570) );
  XNOR2_X1 U626 ( .A(n570), .B(KEYINPUT78), .ZN(n576) );
  NAND2_X1 U627 ( .A1(G49), .A2(n787), .ZN(n573) );
  NAND2_X1 U628 ( .A1(G87), .A2(n571), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U630 ( .A1(n782), .A2(n574), .ZN(n575) );
  NAND2_X1 U631 ( .A1(n576), .A2(n575), .ZN(G288) );
  NAND2_X1 U632 ( .A1(G73), .A2(n783), .ZN(n577) );
  XOR2_X1 U633 ( .A(KEYINPUT2), .B(n577), .Z(n584) );
  NAND2_X1 U634 ( .A1(n782), .A2(G61), .ZN(n578) );
  XNOR2_X1 U635 ( .A(KEYINPUT79), .B(n578), .ZN(n581) );
  NAND2_X1 U636 ( .A1(n786), .A2(G86), .ZN(n579) );
  XOR2_X1 U637 ( .A(KEYINPUT80), .B(n579), .Z(n580) );
  NOR2_X1 U638 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U639 ( .A(n582), .B(KEYINPUT81), .ZN(n583) );
  NOR2_X1 U640 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U641 ( .A1(n787), .A2(G48), .ZN(n585) );
  NAND2_X1 U642 ( .A1(n586), .A2(n585), .ZN(G305) );
  NAND2_X1 U643 ( .A1(G72), .A2(n783), .ZN(n588) );
  NAND2_X1 U644 ( .A1(G85), .A2(n786), .ZN(n587) );
  NAND2_X1 U645 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U646 ( .A1(G60), .A2(n782), .ZN(n590) );
  NAND2_X1 U647 ( .A1(G47), .A2(n787), .ZN(n589) );
  NAND2_X1 U648 ( .A1(n590), .A2(n589), .ZN(n591) );
  OR2_X1 U649 ( .A1(n592), .A2(n591), .ZN(G290) );
  NOR2_X1 U650 ( .A1(G164), .A2(G1384), .ZN(n615) );
  NAND2_X1 U651 ( .A1(G160), .A2(G40), .ZN(n613) );
  NOR2_X1 U652 ( .A1(n615), .A2(n613), .ZN(n749) );
  XNOR2_X1 U653 ( .A(n749), .B(KEYINPUT94), .ZN(n611) );
  NAND2_X1 U654 ( .A1(G141), .A2(n991), .ZN(n594) );
  NAND2_X1 U655 ( .A1(G129), .A2(n987), .ZN(n593) );
  NAND2_X1 U656 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U657 ( .A1(G105), .A2(n990), .ZN(n595) );
  XNOR2_X1 U658 ( .A(n595), .B(KEYINPUT38), .ZN(n596) );
  XNOR2_X1 U659 ( .A(n596), .B(KEYINPUT93), .ZN(n597) );
  NOR2_X1 U660 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U661 ( .A1(n548), .A2(G117), .ZN(n599) );
  NAND2_X1 U662 ( .A1(n600), .A2(n599), .ZN(n983) );
  NAND2_X1 U663 ( .A1(G1996), .A2(n983), .ZN(n610) );
  NAND2_X1 U664 ( .A1(G131), .A2(n991), .ZN(n601) );
  XNOR2_X1 U665 ( .A(n601), .B(KEYINPUT92), .ZN(n608) );
  NAND2_X1 U666 ( .A1(G95), .A2(n990), .ZN(n603) );
  NAND2_X1 U667 ( .A1(G119), .A2(n987), .ZN(n602) );
  NAND2_X1 U668 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U669 ( .A1(G107), .A2(n548), .ZN(n604) );
  XNOR2_X1 U670 ( .A(KEYINPUT91), .B(n604), .ZN(n605) );
  NOR2_X1 U671 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U672 ( .A1(n608), .A2(n607), .ZN(n1003) );
  NAND2_X1 U673 ( .A1(G1991), .A2(n1003), .ZN(n609) );
  NAND2_X1 U674 ( .A1(n610), .A2(n609), .ZN(n859) );
  NAND2_X1 U675 ( .A1(n611), .A2(n859), .ZN(n612) );
  XNOR2_X1 U676 ( .A(n612), .B(KEYINPUT95), .ZN(n742) );
  XOR2_X1 U677 ( .A(KEYINPUT96), .B(n613), .Z(n614) );
  INV_X1 U678 ( .A(n678), .ZN(n653) );
  NOR2_X1 U679 ( .A1(n653), .A2(G1961), .ZN(n616) );
  XOR2_X1 U680 ( .A(KEYINPUT98), .B(n616), .Z(n618) );
  XNOR2_X1 U681 ( .A(G2078), .B(KEYINPUT25), .ZN(n889) );
  NAND2_X1 U682 ( .A1(n653), .A2(n889), .ZN(n617) );
  NAND2_X1 U683 ( .A1(n618), .A2(n617), .ZN(n672) );
  NAND2_X1 U684 ( .A1(n672), .A2(G171), .ZN(n668) );
  NAND2_X1 U685 ( .A1(n653), .A2(G2072), .ZN(n619) );
  XNOR2_X1 U686 ( .A(n619), .B(KEYINPUT27), .ZN(n621) );
  AND2_X1 U687 ( .A1(G1956), .A2(n678), .ZN(n620) );
  NOR2_X1 U688 ( .A1(n621), .A2(n620), .ZN(n661) );
  NAND2_X1 U689 ( .A1(G65), .A2(n782), .ZN(n623) );
  NAND2_X1 U690 ( .A1(G53), .A2(n787), .ZN(n622) );
  NAND2_X1 U691 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U692 ( .A1(G78), .A2(n783), .ZN(n625) );
  NAND2_X1 U693 ( .A1(G91), .A2(n786), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U695 ( .A1(n627), .A2(n626), .ZN(n795) );
  NOR2_X1 U696 ( .A1(n661), .A2(n795), .ZN(n628) );
  XOR2_X1 U697 ( .A(n628), .B(KEYINPUT28), .Z(n665) );
  NAND2_X1 U698 ( .A1(G66), .A2(n782), .ZN(n630) );
  NAND2_X1 U699 ( .A1(G79), .A2(n783), .ZN(n629) );
  NAND2_X1 U700 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U701 ( .A1(G92), .A2(n786), .ZN(n632) );
  NAND2_X1 U702 ( .A1(G54), .A2(n787), .ZN(n631) );
  NAND2_X1 U703 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U705 ( .A(KEYINPUT15), .B(n635), .Z(n1012) );
  NAND2_X1 U706 ( .A1(n782), .A2(G56), .ZN(n636) );
  XOR2_X1 U707 ( .A(KEYINPUT14), .B(n636), .Z(n644) );
  NAND2_X1 U708 ( .A1(n786), .A2(G81), .ZN(n637) );
  XOR2_X1 U709 ( .A(KEYINPUT12), .B(n637), .Z(n640) );
  NAND2_X1 U710 ( .A1(n783), .A2(G68), .ZN(n638) );
  XOR2_X1 U711 ( .A(n638), .B(KEYINPUT66), .Z(n639) );
  XOR2_X1 U712 ( .A(KEYINPUT67), .B(n641), .Z(n642) );
  XNOR2_X1 U713 ( .A(n642), .B(KEYINPUT13), .ZN(n643) );
  NOR2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U715 ( .A1(n787), .A2(G43), .ZN(n645) );
  NAND2_X1 U716 ( .A1(n646), .A2(n645), .ZN(n1009) );
  XNOR2_X1 U717 ( .A(G1996), .B(KEYINPUT99), .ZN(n883) );
  INV_X1 U718 ( .A(KEYINPUT26), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n648), .B(n647), .ZN(n650) );
  NAND2_X1 U720 ( .A1(n678), .A2(G1341), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U722 ( .A1(n1009), .A2(n651), .ZN(n652) );
  OR2_X1 U723 ( .A1(n1012), .A2(n652), .ZN(n660) );
  NAND2_X1 U724 ( .A1(n652), .A2(n1012), .ZN(n658) );
  AND2_X1 U725 ( .A1(n653), .A2(G2067), .ZN(n654) );
  XOR2_X1 U726 ( .A(n654), .B(KEYINPUT100), .Z(n656) );
  NAND2_X1 U727 ( .A1(n678), .A2(G1348), .ZN(n655) );
  NAND2_X1 U728 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U729 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U730 ( .A1(n660), .A2(n659), .ZN(n663) );
  NAND2_X1 U731 ( .A1(n795), .A2(n661), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U733 ( .A1(n668), .A2(n667), .ZN(n677) );
  NAND2_X1 U734 ( .A1(G8), .A2(n678), .ZN(n719) );
  NOR2_X1 U735 ( .A1(G1966), .A2(n719), .ZN(n689) );
  NOR2_X1 U736 ( .A1(G2084), .A2(n678), .ZN(n686) );
  NOR2_X1 U737 ( .A1(n689), .A2(n686), .ZN(n669) );
  NAND2_X1 U738 ( .A1(G8), .A2(n669), .ZN(n670) );
  XNOR2_X1 U739 ( .A(KEYINPUT30), .B(n670), .ZN(n671) );
  NOR2_X1 U740 ( .A1(G168), .A2(n671), .ZN(n674) );
  NOR2_X1 U741 ( .A1(G171), .A2(n672), .ZN(n673) );
  NOR2_X1 U742 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U743 ( .A(KEYINPUT31), .B(n675), .Z(n676) );
  NAND2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n687) );
  NAND2_X1 U745 ( .A1(n687), .A2(G286), .ZN(n683) );
  NOR2_X1 U746 ( .A1(G1971), .A2(n719), .ZN(n680) );
  NOR2_X1 U747 ( .A1(G2090), .A2(n678), .ZN(n679) );
  NOR2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U749 ( .A1(n681), .A2(G303), .ZN(n682) );
  NAND2_X1 U750 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U751 ( .A1(n684), .A2(G8), .ZN(n685) );
  XNOR2_X1 U752 ( .A(n685), .B(KEYINPUT32), .ZN(n693) );
  NAND2_X1 U753 ( .A1(G8), .A2(n686), .ZN(n691) );
  INV_X1 U754 ( .A(n687), .ZN(n688) );
  NOR2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n713) );
  NOR2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n699) );
  NOR2_X1 U759 ( .A1(G303), .A2(G1971), .ZN(n694) );
  NOR2_X1 U760 ( .A1(n699), .A2(n694), .ZN(n916) );
  NAND2_X1 U761 ( .A1(n713), .A2(n916), .ZN(n696) );
  NAND2_X1 U762 ( .A1(G288), .A2(G1976), .ZN(n695) );
  XOR2_X1 U763 ( .A(KEYINPUT101), .B(n695), .Z(n915) );
  NAND2_X1 U764 ( .A1(n696), .A2(n915), .ZN(n698) );
  XNOR2_X1 U765 ( .A(n698), .B(n697), .ZN(n706) );
  INV_X1 U766 ( .A(n719), .ZN(n702) );
  INV_X1 U767 ( .A(KEYINPUT33), .ZN(n708) );
  NAND2_X1 U768 ( .A1(n702), .A2(n699), .ZN(n700) );
  NOR2_X1 U769 ( .A1(n708), .A2(n700), .ZN(n701) );
  XNOR2_X1 U770 ( .A(n701), .B(KEYINPUT103), .ZN(n707) );
  AND2_X1 U771 ( .A1(n702), .A2(n707), .ZN(n704) );
  XNOR2_X1 U772 ( .A(G1981), .B(G305), .ZN(n905) );
  INV_X1 U773 ( .A(n905), .ZN(n703) );
  AND2_X1 U774 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U775 ( .A1(n706), .A2(n705), .ZN(n712) );
  INV_X1 U776 ( .A(n707), .ZN(n709) );
  OR2_X1 U777 ( .A1(n709), .A2(n708), .ZN(n710) );
  OR2_X1 U778 ( .A1(n905), .A2(n710), .ZN(n711) );
  NAND2_X1 U779 ( .A1(n712), .A2(n711), .ZN(n723) );
  NOR2_X1 U780 ( .A1(G2090), .A2(G303), .ZN(n714) );
  NAND2_X1 U781 ( .A1(G8), .A2(n714), .ZN(n715) );
  NAND2_X1 U782 ( .A1(n713), .A2(n715), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n716), .A2(n719), .ZN(n721) );
  NOR2_X1 U784 ( .A1(G1981), .A2(G305), .ZN(n717) );
  XNOR2_X1 U785 ( .A(n717), .B(KEYINPUT97), .ZN(n718) );
  XNOR2_X1 U786 ( .A(n718), .B(KEYINPUT24), .ZN(n720) );
  OR2_X1 U787 ( .A1(n723), .A2(n722), .ZN(n735) );
  NAND2_X1 U788 ( .A1(n991), .A2(G140), .ZN(n724) );
  XOR2_X1 U789 ( .A(KEYINPUT89), .B(n724), .Z(n726) );
  NAND2_X1 U790 ( .A1(n990), .A2(G104), .ZN(n725) );
  NAND2_X1 U791 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U792 ( .A(KEYINPUT34), .B(n727), .ZN(n733) );
  NAND2_X1 U793 ( .A1(G116), .A2(n548), .ZN(n729) );
  NAND2_X1 U794 ( .A1(G128), .A2(n987), .ZN(n728) );
  NAND2_X1 U795 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U796 ( .A(KEYINPUT90), .B(n730), .Z(n731) );
  XNOR2_X1 U797 ( .A(KEYINPUT35), .B(n731), .ZN(n732) );
  NOR2_X1 U798 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U799 ( .A(KEYINPUT36), .B(n734), .ZN(n1006) );
  XNOR2_X1 U800 ( .A(G2067), .B(KEYINPUT37), .ZN(n739) );
  NOR2_X1 U801 ( .A1(n1006), .A2(n739), .ZN(n872) );
  NAND2_X1 U802 ( .A1(n749), .A2(n872), .ZN(n746) );
  NAND2_X1 U803 ( .A1(n735), .A2(n746), .ZN(n736) );
  NOR2_X1 U804 ( .A1(n742), .A2(n736), .ZN(n738) );
  XNOR2_X1 U805 ( .A(G1986), .B(G290), .ZN(n912) );
  NAND2_X1 U806 ( .A1(n912), .A2(n749), .ZN(n737) );
  NAND2_X1 U807 ( .A1(n738), .A2(n737), .ZN(n752) );
  NAND2_X1 U808 ( .A1(n1006), .A2(n739), .ZN(n869) );
  NOR2_X1 U809 ( .A1(G1996), .A2(n983), .ZN(n864) );
  NOR2_X1 U810 ( .A1(G1986), .A2(G290), .ZN(n740) );
  NOR2_X1 U811 ( .A1(G1991), .A2(n1003), .ZN(n860) );
  NOR2_X1 U812 ( .A1(n740), .A2(n860), .ZN(n741) );
  NOR2_X1 U813 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U814 ( .A1(n864), .A2(n743), .ZN(n744) );
  XNOR2_X1 U815 ( .A(KEYINPUT104), .B(n744), .ZN(n745) );
  XNOR2_X1 U816 ( .A(n745), .B(KEYINPUT39), .ZN(n747) );
  NAND2_X1 U817 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U818 ( .A1(n869), .A2(n748), .ZN(n750) );
  NAND2_X1 U819 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U820 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U821 ( .A(n753), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U822 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U823 ( .A(n795), .ZN(G299) );
  INV_X1 U824 ( .A(G120), .ZN(G236) );
  INV_X1 U825 ( .A(G69), .ZN(G235) );
  INV_X1 U826 ( .A(G108), .ZN(G238) );
  NAND2_X1 U827 ( .A1(G7), .A2(G661), .ZN(n754) );
  XNOR2_X1 U828 ( .A(n754), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U829 ( .A(G223), .ZN(n831) );
  NAND2_X1 U830 ( .A1(n831), .A2(G567), .ZN(n755) );
  XOR2_X1 U831 ( .A(KEYINPUT11), .B(n755), .Z(G234) );
  INV_X1 U832 ( .A(G860), .ZN(n781) );
  OR2_X1 U833 ( .A1(n1009), .A2(n781), .ZN(G153) );
  INV_X1 U834 ( .A(G171), .ZN(G301) );
  INV_X1 U835 ( .A(n1012), .ZN(n907) );
  INV_X1 U836 ( .A(G868), .ZN(n802) );
  NAND2_X1 U837 ( .A1(n907), .A2(n802), .ZN(n756) );
  XNOR2_X1 U838 ( .A(n756), .B(KEYINPUT68), .ZN(n758) );
  NAND2_X1 U839 ( .A1(G868), .A2(G301), .ZN(n757) );
  NAND2_X1 U840 ( .A1(n758), .A2(n757), .ZN(G284) );
  NAND2_X1 U841 ( .A1(G868), .A2(G286), .ZN(n760) );
  NAND2_X1 U842 ( .A1(G299), .A2(n802), .ZN(n759) );
  NAND2_X1 U843 ( .A1(n760), .A2(n759), .ZN(G297) );
  NAND2_X1 U844 ( .A1(n781), .A2(G559), .ZN(n761) );
  NAND2_X1 U845 ( .A1(n761), .A2(n1012), .ZN(n762) );
  XNOR2_X1 U846 ( .A(n762), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U847 ( .A1(G868), .A2(n1009), .ZN(n765) );
  NAND2_X1 U848 ( .A1(G868), .A2(n1012), .ZN(n763) );
  NOR2_X1 U849 ( .A1(G559), .A2(n763), .ZN(n764) );
  NOR2_X1 U850 ( .A1(n765), .A2(n764), .ZN(G282) );
  NAND2_X1 U851 ( .A1(G135), .A2(n991), .ZN(n766) );
  XNOR2_X1 U852 ( .A(n766), .B(KEYINPUT74), .ZN(n775) );
  NAND2_X1 U853 ( .A1(G123), .A2(n987), .ZN(n767) );
  XOR2_X1 U854 ( .A(KEYINPUT18), .B(n767), .Z(n768) );
  XNOR2_X1 U855 ( .A(n768), .B(KEYINPUT73), .ZN(n770) );
  NAND2_X1 U856 ( .A1(G99), .A2(n990), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n773) );
  NAND2_X1 U858 ( .A1(G111), .A2(n548), .ZN(n771) );
  XNOR2_X1 U859 ( .A(KEYINPUT75), .B(n771), .ZN(n772) );
  NOR2_X1 U860 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U862 ( .A(KEYINPUT76), .B(n776), .Z(n985) );
  XNOR2_X1 U863 ( .A(n985), .B(G2096), .ZN(n778) );
  INV_X1 U864 ( .A(G2100), .ZN(n777) );
  NAND2_X1 U865 ( .A1(n778), .A2(n777), .ZN(G156) );
  XNOR2_X1 U866 ( .A(n1009), .B(KEYINPUT77), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n1012), .A2(G559), .ZN(n779) );
  XNOR2_X1 U868 ( .A(n780), .B(n779), .ZN(n799) );
  NAND2_X1 U869 ( .A1(n781), .A2(n799), .ZN(n792) );
  NAND2_X1 U870 ( .A1(G67), .A2(n782), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G80), .A2(n783), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n791) );
  NAND2_X1 U873 ( .A1(G93), .A2(n786), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G55), .A2(n787), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U876 ( .A1(n791), .A2(n790), .ZN(n801) );
  XOR2_X1 U877 ( .A(n792), .B(n801), .Z(G145) );
  INV_X1 U878 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U879 ( .A(KEYINPUT19), .B(G288), .ZN(n798) );
  XNOR2_X1 U880 ( .A(n801), .B(G166), .ZN(n793) );
  XNOR2_X1 U881 ( .A(n793), .B(G305), .ZN(n794) );
  XNOR2_X1 U882 ( .A(n795), .B(n794), .ZN(n796) );
  XNOR2_X1 U883 ( .A(n796), .B(G290), .ZN(n797) );
  XNOR2_X1 U884 ( .A(n798), .B(n797), .ZN(n1010) );
  XOR2_X1 U885 ( .A(n1010), .B(n799), .Z(n800) );
  NOR2_X1 U886 ( .A1(n802), .A2(n800), .ZN(n804) );
  AND2_X1 U887 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U888 ( .A1(n804), .A2(n803), .ZN(G295) );
  NAND2_X1 U889 ( .A1(G2078), .A2(G2084), .ZN(n805) );
  XOR2_X1 U890 ( .A(KEYINPUT20), .B(n805), .Z(n806) );
  NAND2_X1 U891 ( .A1(G2090), .A2(n806), .ZN(n807) );
  XNOR2_X1 U892 ( .A(KEYINPUT21), .B(n807), .ZN(n808) );
  NAND2_X1 U893 ( .A1(n808), .A2(G2072), .ZN(G158) );
  XOR2_X1 U894 ( .A(KEYINPUT83), .B(G44), .Z(n809) );
  XNOR2_X1 U895 ( .A(KEYINPUT3), .B(n809), .ZN(G218) );
  NOR2_X1 U896 ( .A1(G235), .A2(G236), .ZN(n810) );
  XNOR2_X1 U897 ( .A(n810), .B(KEYINPUT85), .ZN(n811) );
  NOR2_X1 U898 ( .A1(G238), .A2(n811), .ZN(n812) );
  NAND2_X1 U899 ( .A1(G57), .A2(n812), .ZN(n960) );
  NAND2_X1 U900 ( .A1(n960), .A2(G567), .ZN(n818) );
  NAND2_X1 U901 ( .A1(G132), .A2(G82), .ZN(n813) );
  XNOR2_X1 U902 ( .A(n813), .B(KEYINPUT22), .ZN(n814) );
  XNOR2_X1 U903 ( .A(n814), .B(KEYINPUT84), .ZN(n815) );
  NOR2_X1 U904 ( .A1(G218), .A2(n815), .ZN(n816) );
  NAND2_X1 U905 ( .A1(G96), .A2(n816), .ZN(n961) );
  NAND2_X1 U906 ( .A1(n961), .A2(G2106), .ZN(n817) );
  NAND2_X1 U907 ( .A1(n818), .A2(n817), .ZN(n980) );
  NAND2_X1 U908 ( .A1(G483), .A2(G661), .ZN(n819) );
  NOR2_X1 U909 ( .A1(n980), .A2(n819), .ZN(n833) );
  NAND2_X1 U910 ( .A1(n833), .A2(G36), .ZN(n820) );
  XNOR2_X1 U911 ( .A(KEYINPUT86), .B(n820), .ZN(G176) );
  XOR2_X1 U912 ( .A(G2443), .B(G2454), .Z(n822) );
  XNOR2_X1 U913 ( .A(G1348), .B(G2435), .ZN(n821) );
  XNOR2_X1 U914 ( .A(n822), .B(n821), .ZN(n829) );
  XOR2_X1 U915 ( .A(KEYINPUT105), .B(G2446), .Z(n824) );
  XNOR2_X1 U916 ( .A(G1341), .B(G2430), .ZN(n823) );
  XNOR2_X1 U917 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U918 ( .A(n825), .B(G2451), .Z(n827) );
  XNOR2_X1 U919 ( .A(G2438), .B(G2427), .ZN(n826) );
  XNOR2_X1 U920 ( .A(n827), .B(n826), .ZN(n828) );
  XNOR2_X1 U921 ( .A(n829), .B(n828), .ZN(n830) );
  NAND2_X1 U922 ( .A1(n830), .A2(G14), .ZN(n1018) );
  XOR2_X1 U923 ( .A(KEYINPUT106), .B(n1018), .Z(G401) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U926 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n834), .A2(n833), .ZN(n835) );
  XOR2_X1 U929 ( .A(KEYINPUT107), .B(n835), .Z(G188) );
  NAND2_X1 U931 ( .A1(G112), .A2(n548), .ZN(n836) );
  XNOR2_X1 U932 ( .A(n836), .B(KEYINPUT110), .ZN(n840) );
  XOR2_X1 U933 ( .A(KEYINPUT109), .B(KEYINPUT44), .Z(n838) );
  NAND2_X1 U934 ( .A1(G124), .A2(n987), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n840), .A2(n839), .ZN(n844) );
  NAND2_X1 U937 ( .A1(G100), .A2(n990), .ZN(n842) );
  NAND2_X1 U938 ( .A1(G136), .A2(n991), .ZN(n841) );
  NAND2_X1 U939 ( .A1(n842), .A2(n841), .ZN(n843) );
  NOR2_X1 U940 ( .A1(n844), .A2(n843), .ZN(G162) );
  XNOR2_X1 U941 ( .A(KEYINPUT50), .B(KEYINPUT118), .ZN(n856) );
  NAND2_X1 U942 ( .A1(G115), .A2(n548), .ZN(n846) );
  NAND2_X1 U943 ( .A1(G127), .A2(n987), .ZN(n845) );
  NAND2_X1 U944 ( .A1(n846), .A2(n845), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n847), .B(KEYINPUT47), .ZN(n849) );
  NAND2_X1 U946 ( .A1(G139), .A2(n991), .ZN(n848) );
  NAND2_X1 U947 ( .A1(n849), .A2(n848), .ZN(n852) );
  NAND2_X1 U948 ( .A1(G103), .A2(n990), .ZN(n850) );
  XNOR2_X1 U949 ( .A(KEYINPUT111), .B(n850), .ZN(n851) );
  NOR2_X1 U950 ( .A1(n852), .A2(n851), .ZN(n984) );
  XNOR2_X1 U951 ( .A(G2072), .B(n984), .ZN(n854) );
  XNOR2_X1 U952 ( .A(G164), .B(G2078), .ZN(n853) );
  NAND2_X1 U953 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n875) );
  XNOR2_X1 U955 ( .A(G160), .B(G2084), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n857), .B(KEYINPUT115), .ZN(n858) );
  NOR2_X1 U957 ( .A1(n858), .A2(n985), .ZN(n862) );
  NOR2_X1 U958 ( .A1(n860), .A2(n859), .ZN(n861) );
  NAND2_X1 U959 ( .A1(n862), .A2(n861), .ZN(n868) );
  XOR2_X1 U960 ( .A(G2090), .B(G162), .Z(n863) );
  NOR2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U962 ( .A(KEYINPUT116), .B(n865), .Z(n866) );
  XOR2_X1 U963 ( .A(KEYINPUT51), .B(n866), .Z(n867) );
  NOR2_X1 U964 ( .A1(n868), .A2(n867), .ZN(n870) );
  NAND2_X1 U965 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U966 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U967 ( .A(n873), .B(KEYINPUT117), .ZN(n874) );
  NOR2_X1 U968 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U969 ( .A(KEYINPUT52), .B(n876), .ZN(n877) );
  INV_X1 U970 ( .A(KEYINPUT55), .ZN(n900) );
  NAND2_X1 U971 ( .A1(n877), .A2(n900), .ZN(n878) );
  NAND2_X1 U972 ( .A1(n878), .A2(G29), .ZN(n958) );
  XNOR2_X1 U973 ( .A(G2090), .B(G35), .ZN(n894) );
  XNOR2_X1 U974 ( .A(G25), .B(G1991), .ZN(n879) );
  XNOR2_X1 U975 ( .A(n879), .B(KEYINPUT119), .ZN(n888) );
  XNOR2_X1 U976 ( .A(G2067), .B(G26), .ZN(n881) );
  XNOR2_X1 U977 ( .A(G33), .B(G2072), .ZN(n880) );
  NOR2_X1 U978 ( .A1(n881), .A2(n880), .ZN(n882) );
  NAND2_X1 U979 ( .A1(G28), .A2(n882), .ZN(n886) );
  XOR2_X1 U980 ( .A(G32), .B(n883), .Z(n884) );
  XNOR2_X1 U981 ( .A(KEYINPUT120), .B(n884), .ZN(n885) );
  NOR2_X1 U982 ( .A1(n886), .A2(n885), .ZN(n887) );
  NAND2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n891) );
  XOR2_X1 U984 ( .A(G27), .B(n889), .Z(n890) );
  NOR2_X1 U985 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U986 ( .A(KEYINPUT53), .B(n892), .ZN(n893) );
  NOR2_X1 U987 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U988 ( .A(KEYINPUT121), .B(n895), .Z(n898) );
  XOR2_X1 U989 ( .A(KEYINPUT54), .B(G34), .Z(n896) );
  XNOR2_X1 U990 ( .A(G2084), .B(n896), .ZN(n897) );
  NAND2_X1 U991 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U992 ( .A(n900), .B(n899), .ZN(n902) );
  INV_X1 U993 ( .A(G29), .ZN(n901) );
  NAND2_X1 U994 ( .A1(n902), .A2(n901), .ZN(n903) );
  NAND2_X1 U995 ( .A1(G11), .A2(n903), .ZN(n956) );
  XNOR2_X1 U996 ( .A(G16), .B(KEYINPUT56), .ZN(n926) );
  XOR2_X1 U997 ( .A(G168), .B(G1966), .Z(n904) );
  NOR2_X1 U998 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U999 ( .A(KEYINPUT57), .B(n906), .Z(n924) );
  XNOR2_X1 U1000 ( .A(G301), .B(G1961), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(n907), .B(G1348), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1003 ( .A(KEYINPUT122), .B(n910), .ZN(n920) );
  XNOR2_X1 U1004 ( .A(G1956), .B(G299), .ZN(n911) );
  NOR2_X1 U1005 ( .A1(n912), .A2(n911), .ZN(n914) );
  NAND2_X1 U1006 ( .A1(G303), .A2(G1971), .ZN(n913) );
  NAND2_X1 U1007 ( .A1(n914), .A2(n913), .ZN(n918) );
  NAND2_X1 U1008 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1009 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1010 ( .A1(n920), .A2(n919), .ZN(n922) );
  XNOR2_X1 U1011 ( .A(G1341), .B(n1009), .ZN(n921) );
  NOR2_X1 U1012 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1013 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1014 ( .A1(n926), .A2(n925), .ZN(n954) );
  INV_X1 U1015 ( .A(G16), .ZN(n952) );
  XNOR2_X1 U1016 ( .A(G1971), .B(G22), .ZN(n928) );
  XNOR2_X1 U1017 ( .A(G23), .B(G1976), .ZN(n927) );
  NOR2_X1 U1018 ( .A1(n928), .A2(n927), .ZN(n930) );
  XOR2_X1 U1019 ( .A(G1986), .B(G24), .Z(n929) );
  NAND2_X1 U1020 ( .A1(n930), .A2(n929), .ZN(n932) );
  XOR2_X1 U1021 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n931) );
  XNOR2_X1 U1022 ( .A(n932), .B(n931), .ZN(n936) );
  XNOR2_X1 U1023 ( .A(G1966), .B(G21), .ZN(n934) );
  XNOR2_X1 U1024 ( .A(G1961), .B(G5), .ZN(n933) );
  NOR2_X1 U1025 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1026 ( .A1(n936), .A2(n935), .ZN(n949) );
  XOR2_X1 U1027 ( .A(G1348), .B(KEYINPUT59), .Z(n937) );
  XNOR2_X1 U1028 ( .A(G4), .B(n937), .ZN(n946) );
  XOR2_X1 U1029 ( .A(G1341), .B(G19), .Z(n938) );
  XNOR2_X1 U1030 ( .A(KEYINPUT123), .B(n938), .ZN(n940) );
  XNOR2_X1 U1031 ( .A(G6), .B(G1981), .ZN(n939) );
  NOR2_X1 U1032 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1033 ( .A(KEYINPUT124), .B(n941), .Z(n943) );
  XNOR2_X1 U1034 ( .A(G1956), .B(G20), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1036 ( .A(n944), .B(KEYINPUT125), .ZN(n945) );
  NOR2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1038 ( .A(KEYINPUT60), .B(n947), .Z(n948) );
  NOR2_X1 U1039 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1040 ( .A(KEYINPUT61), .B(n950), .ZN(n951) );
  NAND2_X1 U1041 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1042 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1043 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1044 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1045 ( .A(KEYINPUT62), .B(n959), .Z(G311) );
  XNOR2_X1 U1046 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1047 ( .A(G132), .ZN(G219) );
  INV_X1 U1048 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1049 ( .A1(n961), .A2(n960), .ZN(G325) );
  INV_X1 U1050 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1051 ( .A(G1986), .B(G1966), .ZN(n971) );
  XOR2_X1 U1052 ( .A(KEYINPUT108), .B(G1971), .Z(n963) );
  XNOR2_X1 U1053 ( .A(G1961), .B(G1956), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(n963), .B(n962), .ZN(n967) );
  XOR2_X1 U1055 ( .A(KEYINPUT41), .B(G1976), .Z(n965) );
  XNOR2_X1 U1056 ( .A(G1996), .B(G1991), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n965), .B(n964), .ZN(n966) );
  XOR2_X1 U1058 ( .A(n967), .B(n966), .Z(n969) );
  XNOR2_X1 U1059 ( .A(G1981), .B(G2474), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n969), .B(n968), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(n971), .B(n970), .ZN(G229) );
  XOR2_X1 U1062 ( .A(G2100), .B(G2096), .Z(n973) );
  XNOR2_X1 U1063 ( .A(G2072), .B(G2090), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(n973), .B(n972), .ZN(n977) );
  XOR2_X1 U1065 ( .A(G2678), .B(KEYINPUT42), .Z(n975) );
  XNOR2_X1 U1066 ( .A(G2067), .B(KEYINPUT43), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n975), .B(n974), .ZN(n976) );
  XOR2_X1 U1068 ( .A(n977), .B(n976), .Z(n979) );
  XNOR2_X1 U1069 ( .A(G2078), .B(G2084), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(n979), .B(n978), .ZN(G227) );
  INV_X1 U1071 ( .A(n980), .ZN(G319) );
  XOR2_X1 U1072 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n982) );
  XNOR2_X1 U1073 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n982), .B(n981), .ZN(n1002) );
  XNOR2_X1 U1075 ( .A(n984), .B(n983), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(n986), .B(n985), .ZN(n998) );
  NAND2_X1 U1077 ( .A1(G118), .A2(n548), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(G130), .A2(n987), .ZN(n988) );
  NAND2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n996) );
  NAND2_X1 U1080 ( .A1(G106), .A2(n990), .ZN(n993) );
  NAND2_X1 U1081 ( .A1(G142), .A2(n991), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1083 ( .A(KEYINPUT45), .B(n994), .Z(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1085 ( .A(n998), .B(n997), .Z(n1000) );
  XNOR2_X1 U1086 ( .A(G164), .B(G160), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(n1000), .B(n999), .ZN(n1001) );
  XNOR2_X1 U1088 ( .A(n1002), .B(n1001), .ZN(n1005) );
  XNOR2_X1 U1089 ( .A(n1003), .B(G162), .ZN(n1004) );
  XNOR2_X1 U1090 ( .A(n1005), .B(n1004), .ZN(n1007) );
  XOR2_X1 U1091 ( .A(n1007), .B(n1006), .Z(n1008) );
  NOR2_X1 U1092 ( .A1(G37), .A2(n1008), .ZN(G395) );
  XNOR2_X1 U1093 ( .A(n1010), .B(n1009), .ZN(n1011) );
  XNOR2_X1 U1094 ( .A(n1011), .B(G286), .ZN(n1014) );
  XOR2_X1 U1095 ( .A(n1012), .B(G171), .Z(n1013) );
  XNOR2_X1 U1096 ( .A(n1014), .B(n1013), .ZN(n1015) );
  NOR2_X1 U1097 ( .A1(G37), .A2(n1015), .ZN(G397) );
  XNOR2_X1 U1098 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n1017) );
  NOR2_X1 U1099 ( .A1(G229), .A2(G227), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(n1017), .B(n1016), .ZN(n1020) );
  NAND2_X1 U1101 ( .A1(G319), .A2(n1018), .ZN(n1019) );
  NOR2_X1 U1102 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  NOR2_X1 U1103 ( .A1(G395), .A2(G397), .ZN(n1021) );
  NAND2_X1 U1104 ( .A1(n1022), .A2(n1021), .ZN(G225) );
  INV_X1 U1105 ( .A(G225), .ZN(G308) );
  INV_X1 U1106 ( .A(G96), .ZN(G221) );
  INV_X1 U1107 ( .A(G57), .ZN(G237) );
endmodule

