//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT70), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G140), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT69), .B(G140), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(new_n192), .ZN(new_n195));
  INV_X1    g009(.A(G140), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n196), .A2(KEYINPUT69), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(KEYINPUT69), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n191), .B(G125), .C1(new_n197), .C2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(KEYINPUT19), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n192), .A2(G140), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT19), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n201), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT83), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n195), .A2(KEYINPUT16), .A3(new_n199), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n202), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT83), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n200), .A2(new_n213), .A3(new_n201), .A4(new_n205), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n207), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G953), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT68), .A2(G237), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT68), .A2(G237), .ZN(new_n218));
  OAI211_X1 g032(.A(G214), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT68), .B(G237), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n222), .A2(KEYINPUT81), .A3(G214), .A4(new_n216), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT82), .ZN(new_n224));
  INV_X1    g038(.A(G143), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n221), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  OR2_X1    g040(.A1(new_n219), .A2(new_n225), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(G143), .B1(new_n219), .B2(new_n220), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n224), .B1(new_n229), .B2(new_n223), .ZN(new_n230));
  OAI21_X1  g044(.A(G131), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n223), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT82), .ZN(new_n233));
  INV_X1    g047(.A(G131), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n233), .A2(new_n234), .A3(new_n227), .A4(new_n226), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n215), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(KEYINPUT18), .B(G131), .C1(new_n228), .C2(new_n230), .ZN(new_n237));
  NAND2_X1  g051(.A1(KEYINPUT18), .A2(G131), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n233), .A2(new_n227), .A3(new_n226), .A4(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n195), .A2(G146), .A3(new_n199), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n202), .A2(new_n203), .A3(new_n201), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n237), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n190), .B1(new_n236), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n237), .A2(new_n239), .A3(new_n242), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT17), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n231), .A2(new_n235), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n201), .B1(new_n208), .B2(new_n210), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n208), .A2(new_n201), .A3(new_n210), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(KEYINPUT71), .ZN(new_n250));
  OAI211_X1 g064(.A(KEYINPUT17), .B(G131), .C1(new_n228), .C2(new_n230), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n208), .A2(new_n201), .A3(new_n210), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n250), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n189), .B(new_n245), .C1(new_n247), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n244), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT20), .ZN(new_n258));
  NOR2_X1   g072(.A1(G475), .A2(G902), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT84), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT84), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n257), .A2(new_n262), .A3(new_n258), .A4(new_n259), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n257), .A2(new_n259), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT20), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n261), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G902), .ZN(new_n267));
  INV_X1    g081(.A(new_n256), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n231), .A2(new_n235), .A3(new_n246), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n269), .A2(new_n254), .A3(new_n250), .A4(new_n251), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n189), .B1(new_n270), .B2(new_n245), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n267), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G475), .ZN(new_n273));
  XNOR2_X1  g087(.A(G116), .B(G122), .ZN(new_n274));
  INV_X1    g088(.A(G107), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n276), .B(KEYINPUT85), .ZN(new_n277));
  XNOR2_X1  g091(.A(G128), .B(G143), .ZN(new_n278));
  INV_X1    g092(.A(G134), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT14), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n274), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G116), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n283), .A2(KEYINPUT14), .A3(G122), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(G107), .A3(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n277), .A2(new_n280), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n274), .B(new_n275), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n278), .A2(new_n279), .ZN(new_n288));
  INV_X1    g102(.A(G128), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G143), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(G143), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(KEYINPUT13), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(KEYINPUT13), .B2(new_n291), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n287), .B(new_n288), .C1(new_n293), .C2(new_n279), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n286), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT9), .B(G234), .ZN(new_n296));
  INV_X1    g110(.A(G217), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n296), .A2(new_n297), .A3(G953), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n286), .A2(new_n294), .A3(new_n298), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n267), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT15), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n304), .A2(KEYINPUT86), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(KEYINPUT86), .ZN(new_n306));
  OAI21_X1  g120(.A(G478), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n303), .B(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(G234), .A2(G237), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(G952), .A3(new_n216), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(G902), .A3(G953), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT21), .B(G898), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n312), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n266), .A2(new_n273), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT87), .ZN(new_n319));
  INV_X1    g133(.A(G469), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G140), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n216), .A2(G227), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n275), .A2(G104), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n188), .A2(G107), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT76), .B(G101), .Z(new_n329));
  OR2_X1    g143(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n275), .A2(G104), .ZN(new_n331));
  AND2_X1   g145(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n328), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G101), .B1(new_n327), .B2(new_n325), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT10), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n201), .A2(G143), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n225), .A2(G146), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(KEYINPUT1), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n341), .A3(G128), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n338), .B(new_n339), .C1(KEYINPUT1), .C2(new_n289), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n336), .A2(new_n337), .A3(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n334), .A2(new_n343), .A3(new_n342), .A4(new_n335), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT10), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT0), .A4(G128), .ZN(new_n350));
  INV_X1    g164(.A(new_n340), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT0), .B(G128), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G101), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(new_n328), .B2(new_n333), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n188), .A2(G107), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n330), .B2(new_n331), .ZN(new_n359));
  NAND2_X1  g173(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n326), .B1(new_n327), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(G101), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n334), .A3(KEYINPUT4), .ZN(new_n363));
  AND3_X1   g177(.A1(new_n357), .A2(KEYINPUT77), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT77), .B1(new_n357), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n349), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT11), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n367), .B1(new_n279), .B2(G137), .ZN(new_n368));
  INV_X1    g182(.A(G137), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(KEYINPUT11), .A3(G134), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n279), .A2(G137), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G131), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n368), .A2(new_n370), .A3(new_n234), .A4(new_n371), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(KEYINPUT66), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(KEYINPUT66), .B1(new_n373), .B2(new_n374), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n366), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n378), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n349), .B(new_n380), .C1(new_n364), .C2(new_n365), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n324), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n334), .A2(new_n335), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n344), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n347), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n373), .A2(new_n374), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT12), .ZN(new_n388));
  AOI22_X1  g202(.A1(new_n387), .A2(KEYINPUT12), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n389), .A2(new_n381), .A3(new_n324), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n320), .B(new_n267), .C1(new_n382), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(G469), .A2(G902), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n389), .A2(new_n381), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n323), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n379), .A2(new_n381), .A3(new_n324), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n391), .B(new_n392), .C1(new_n320), .C2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G221), .B1(new_n296), .B2(G902), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n398), .B(KEYINPUT74), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G214), .B1(G237), .B2(G902), .ZN(new_n401));
  XOR2_X1   g215(.A(new_n401), .B(KEYINPUT78), .Z(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G119), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G116), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n283), .A2(G119), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT2), .B(G113), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT65), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G113), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT2), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT2), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G113), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G116), .B(G119), .ZN(new_n417));
  AOI21_X1  g231(.A(KEYINPUT65), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n409), .B1(new_n411), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n355), .A2(new_n356), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n363), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G110), .B(G122), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n410), .B1(new_n407), .B2(new_n408), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n416), .A2(new_n417), .A3(KEYINPUT65), .ZN(new_n424));
  INV_X1    g238(.A(new_n405), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT5), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n412), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT5), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n423), .A2(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(new_n334), .A3(new_n335), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n421), .A2(new_n422), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n428), .A2(KEYINPUT79), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n427), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n428), .A2(KEYINPUT79), .ZN(new_n434));
  OAI22_X1  g248(.A1(new_n433), .A2(new_n434), .B1(new_n411), .B2(new_n418), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n336), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n422), .B(KEYINPUT8), .Z(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n429), .B2(new_n383), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n342), .A2(new_n192), .A3(new_n343), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n350), .B(G125), .C1(new_n351), .C2(new_n352), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n216), .A2(G224), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT7), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT7), .A4(new_n443), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n431), .A2(new_n439), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n267), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT80), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n421), .A2(new_n430), .ZN(new_n452));
  INV_X1    g266(.A(new_n422), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT6), .A3(new_n431), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(new_n456), .A3(new_n453), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n442), .B(new_n443), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n448), .A2(KEYINPUT80), .A3(new_n267), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n451), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G210), .B1(G237), .B2(G902), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n451), .A2(new_n459), .A3(new_n462), .A4(new_n460), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n397), .A2(new_n400), .A3(new_n403), .A4(new_n466), .ZN(new_n467));
  OR3_X1    g281(.A1(new_n318), .A2(new_n319), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G472), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n386), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n353), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n472), .A3(new_n375), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n369), .A2(G134), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n371), .A3(KEYINPUT64), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n475), .B(G131), .C1(KEYINPUT64), .C2(new_n474), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n345), .A2(new_n374), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(KEYINPUT30), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT30), .ZN(new_n479));
  AND4_X1   g293(.A1(new_n374), .A2(new_n476), .A3(new_n343), .A4(new_n342), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n353), .B1(new_n374), .B2(new_n373), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(new_n419), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT67), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n419), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(KEYINPUT67), .B(new_n409), .C1(new_n411), .C2(new_n418), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n473), .A2(new_n477), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n222), .A2(new_n216), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(G210), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT27), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT27), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(new_n492), .A3(G210), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT26), .B(G101), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n494), .B1(new_n491), .B2(new_n493), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n488), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT29), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT28), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n487), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n480), .B1(new_n378), .B2(new_n472), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n485), .A2(new_n486), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n480), .A2(new_n481), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n503), .A2(new_n505), .B1(new_n506), .B2(new_n419), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n502), .B1(new_n507), .B2(new_n501), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n499), .B(new_n500), .C1(new_n508), .C2(new_n498), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n473), .A2(new_n477), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n504), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n501), .B1(new_n511), .B2(new_n487), .ZN(new_n512));
  INV_X1    g326(.A(new_n502), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n498), .A2(new_n500), .ZN(new_n515));
  AOI21_X1  g329(.A(G902), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n469), .B1(new_n509), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n483), .A2(new_n497), .A3(new_n487), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT31), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n483), .A2(new_n497), .A3(KEYINPUT31), .A4(new_n487), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n520), .A2(new_n521), .B1(new_n508), .B2(new_n498), .ZN(new_n522));
  NOR2_X1   g336(.A1(G472), .A2(G902), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT32), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n520), .A2(new_n521), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n508), .A2(new_n498), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT32), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n523), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n517), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n297), .B1(G234), .B2(new_n267), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n289), .A2(KEYINPUT23), .A3(G119), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n404), .A2(G128), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n404), .A2(G128), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n534), .B(new_n535), .C1(new_n536), .C2(KEYINPUT23), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(G110), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n289), .A2(G119), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n535), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT24), .B(G110), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n212), .B(new_n241), .C1(new_n538), .C2(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n208), .A2(KEYINPUT71), .A3(new_n201), .A4(new_n210), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n254), .A2(new_n212), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT72), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n540), .A2(new_n541), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(G110), .B2(new_n537), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n546), .B1(new_n545), .B2(new_n548), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n543), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT22), .B(G137), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n216), .A2(G221), .A3(G234), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n543), .B(new_n554), .C1(new_n549), .C2(new_n550), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n267), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT25), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n556), .A2(KEYINPUT25), .A3(new_n267), .A4(new_n557), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n533), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n556), .A2(new_n557), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n532), .A2(G902), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n564), .B(KEYINPUT73), .Z(new_n565));
  NOR2_X1   g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n531), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n319), .B1(new_n318), .B2(new_n467), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n468), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n569), .B(new_n329), .Z(G3));
  NAND2_X1  g384(.A1(new_n560), .A2(new_n561), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n566), .B1(new_n571), .B2(new_n532), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n522), .A2(G902), .ZN(new_n574));
  OAI22_X1  g388(.A1(new_n574), .A2(new_n469), .B1(new_n522), .B2(new_n524), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n397), .A2(new_n400), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n267), .A2(G478), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT90), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n300), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n302), .A2(new_n581), .A3(KEYINPUT33), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT33), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n300), .B(new_n301), .C1(new_n580), .C2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n579), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n303), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT91), .B1(new_n588), .B2(G478), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n587), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n266), .B2(new_n273), .ZN(new_n591));
  INV_X1    g405(.A(new_n401), .ZN(new_n592));
  AND4_X1   g406(.A1(new_n462), .A2(new_n451), .A3(new_n459), .A4(new_n460), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT88), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n464), .A2(KEYINPUT88), .A3(new_n465), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT89), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n316), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT89), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n591), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n578), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT34), .B(G104), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  INV_X1    g419(.A(KEYINPUT92), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n245), .B1(new_n247), .B2(new_n255), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n190), .ZN(new_n608));
  AOI21_X1  g422(.A(G902), .B1(new_n608), .B2(new_n256), .ZN(new_n609));
  INV_X1    g423(.A(G475), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n272), .A2(KEYINPUT92), .A3(G475), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n309), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n316), .B(KEYINPUT93), .Z(new_n618));
  NAND4_X1  g432(.A1(new_n617), .A2(new_n599), .A3(new_n601), .A4(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n578), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT35), .B(G107), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  NAND2_X1  g436(.A1(new_n551), .A2(KEYINPUT94), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n555), .A2(KEYINPUT36), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT94), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n625), .B(new_n543), .C1(new_n549), .C2(new_n550), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n624), .B1(new_n623), .B2(new_n626), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n627), .A2(new_n628), .A3(new_n565), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n562), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n575), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n468), .A2(new_n568), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT37), .B(G110), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT95), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n632), .B(new_n634), .ZN(G12));
  AND3_X1   g449(.A1(new_n595), .A2(new_n596), .A3(KEYINPUT89), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT89), .B1(new_n595), .B2(new_n596), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n397), .A2(new_n400), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n571), .A2(new_n532), .ZN(new_n640));
  OR3_X1    g454(.A1(new_n627), .A2(new_n628), .A3(new_n565), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n531), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n313), .A2(G900), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n311), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n613), .A2(new_n616), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT96), .B(G128), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G30));
  XNOR2_X1  g464(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n466), .B(new_n651), .Z(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n592), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n511), .A2(new_n487), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n267), .B1(new_n654), .B2(new_n497), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n498), .B1(new_n483), .B2(new_n487), .ZN(new_n656));
  OAI21_X1  g470(.A(G472), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n657), .A2(KEYINPUT98), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(KEYINPUT98), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n525), .A2(new_n530), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n660), .A2(new_n562), .A3(new_n629), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n308), .B1(new_n266), .B2(new_n273), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n645), .B(KEYINPUT39), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  OR3_X1    g480(.A1(new_n638), .A2(KEYINPUT99), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT99), .B1(new_n638), .B2(new_n666), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT40), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n667), .A2(KEYINPUT40), .A3(new_n668), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n664), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n225), .ZN(G45));
  AOI211_X1 g486(.A(new_n590), .B(new_n646), .C1(new_n266), .C2(new_n273), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n643), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  OAI21_X1  g489(.A(new_n267), .B1(new_n382), .B2(new_n390), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G469), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n391), .A3(new_n398), .ZN(new_n678));
  NOR4_X1   g492(.A1(new_n531), .A2(new_n562), .A3(new_n566), .A4(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n636), .A2(new_n637), .A3(new_n316), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n680), .A3(new_n591), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G15));
  INV_X1    g497(.A(new_n618), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n636), .A2(new_n637), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n679), .A2(new_n685), .A3(new_n617), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G116), .ZN(G18));
  NOR2_X1   g501(.A1(new_n636), .A2(new_n637), .ZN(new_n688));
  INV_X1    g502(.A(new_n318), .ZN(new_n689));
  INV_X1    g503(.A(new_n678), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n642), .A2(new_n688), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n636), .A2(new_n637), .A3(new_n678), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n694), .A2(KEYINPUT100), .A3(new_n689), .A4(new_n642), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  OR2_X1    g511(.A1(new_n512), .A2(new_n513), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n698), .A2(new_n498), .B1(new_n520), .B2(new_n521), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n523), .B(KEYINPUT101), .ZN(new_n700));
  OAI22_X1  g514(.A1(new_n574), .A2(new_n469), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n701), .A2(new_n562), .A3(new_n566), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n678), .A2(new_n684), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n702), .A2(new_n688), .A3(new_n663), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  NOR2_X1   g519(.A1(new_n699), .A2(new_n700), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n528), .A2(new_n267), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n706), .B1(G472), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n562), .B2(new_n629), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n694), .A3(new_n673), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT102), .B(G125), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G27));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n525), .A2(new_n530), .ZN(new_n715));
  INV_X1    g529(.A(new_n517), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n466), .A2(new_n592), .ZN(new_n718));
  INV_X1    g532(.A(new_n398), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n391), .A2(new_n392), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n396), .A2(KEYINPUT103), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n395), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n721), .A2(G469), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n719), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n572), .A2(new_n717), .A3(new_n718), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n591), .A2(new_n645), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n714), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n725), .A2(new_n718), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n673), .A2(new_n567), .A3(new_n729), .A4(KEYINPUT42), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G131), .ZN(G33));
  NAND3_X1  g546(.A1(new_n567), .A2(new_n729), .A3(new_n647), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  NAND3_X1  g548(.A1(new_n721), .A2(KEYINPUT45), .A3(new_n723), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n320), .B1(new_n396), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n738), .A2(new_n392), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n739), .A2(KEYINPUT46), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n392), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT104), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(KEYINPUT104), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n740), .A2(new_n391), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n398), .ZN(new_n745));
  INV_X1    g559(.A(new_n718), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n745), .A2(new_n666), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n575), .B1(new_n562), .B2(new_n629), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n266), .A2(new_n273), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n590), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n750), .B(new_n751), .C1(new_n755), .C2(KEYINPUT43), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n748), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT106), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n758), .A2(new_n761), .A3(new_n759), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT106), .B1(new_n757), .B2(KEYINPUT44), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n747), .B(new_n760), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G137), .ZN(G39));
  NOR4_X1   g579(.A1(new_n727), .A2(new_n717), .A3(new_n572), .A4(new_n746), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT47), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n745), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT47), .B1(new_n744), .B2(new_n398), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(KEYINPUT107), .B(G140), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n770), .B(new_n771), .ZN(G42));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n639), .B(new_n642), .C1(new_n647), .C2(new_n673), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n725), .A2(new_n645), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n661), .A2(new_n688), .A3(new_n775), .A4(new_n663), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n711), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT52), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n774), .A2(new_n711), .A3(new_n779), .A4(new_n776), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n778), .A2(KEYINPUT110), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n572), .A2(new_n717), .A3(new_n690), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n602), .B2(new_n619), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n663), .A2(new_n599), .A3(new_n601), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n572), .A2(new_n708), .A3(new_n703), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n467), .A2(new_n684), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n749), .A2(new_n751), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n266), .A2(new_n273), .A3(new_n309), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n591), .A2(KEYINPUT109), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n576), .B(new_n792), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n468), .B(new_n568), .C1(new_n631), .C2(new_n567), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n696), .A2(new_n791), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n725), .A2(new_n718), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n709), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n718), .A2(new_n397), .A3(new_n400), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n308), .B(new_n645), .C1(new_n614), .C2(new_n615), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n803), .A2(new_n804), .A3(new_n613), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n802), .A2(new_n673), .B1(new_n805), .B2(new_n642), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n731), .A2(new_n733), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n800), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n785), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n781), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n808), .A2(KEYINPUT53), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n773), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n800), .A2(new_n810), .A3(new_n807), .ZN(new_n815));
  INV_X1    g629(.A(new_n784), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT110), .B1(new_n778), .B2(new_n780), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n681), .A2(new_n686), .A3(new_n704), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n693), .B2(new_n695), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n798), .A2(new_n799), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n731), .A2(new_n733), .A3(new_n806), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n810), .B1(new_n823), .B2(new_n781), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n818), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(KEYINPUT54), .ZN(new_n826));
  OR2_X1    g640(.A1(new_n814), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n702), .A2(new_n312), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n754), .B2(new_n756), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n745), .B(new_n767), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n677), .A2(new_n391), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT108), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n400), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n718), .B(new_n829), .C1(new_n830), .C2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n678), .A2(new_n401), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n652), .B1(new_n835), .B2(KEYINPUT111), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(KEYINPUT111), .B2(new_n835), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n829), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT50), .Z(new_n839));
  NAND3_X1  g653(.A1(new_n690), .A2(new_n312), .A3(new_n718), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n754), .B2(new_n756), .ZN(new_n841));
  INV_X1    g655(.A(new_n660), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n573), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n749), .A2(new_n751), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n841), .A2(new_n710), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n834), .A2(new_n839), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n843), .A2(new_n591), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(G952), .A3(new_n216), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n829), .A2(new_n694), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(KEYINPUT112), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n841), .A2(new_n567), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT48), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OR2_X1    g670(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  AOI211_X1 g671(.A(new_n851), .B(new_n853), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n848), .A2(new_n849), .A3(new_n858), .ZN(new_n859));
  OAI22_X1  g673(.A1(new_n827), .A2(new_n859), .B1(G952), .B2(G953), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n832), .B(KEYINPUT49), .Z(new_n861));
  AND4_X1   g675(.A1(new_n572), .A2(new_n652), .A3(new_n400), .A4(new_n403), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n660), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n860), .B1(new_n752), .B2(new_n863), .ZN(G75));
  NOR2_X1   g678(.A1(new_n216), .A2(G952), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n696), .A2(new_n791), .A3(new_n798), .A4(new_n799), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n822), .A3(new_n780), .A4(new_n778), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n785), .A2(new_n815), .B1(new_n868), .B2(new_n810), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n267), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT56), .B1(new_n870), .B2(G210), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n455), .A2(new_n457), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT113), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n458), .B(KEYINPUT55), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n873), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n866), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n871), .B2(new_n875), .ZN(G51));
  INV_X1    g691(.A(KEYINPUT114), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n825), .B2(KEYINPUT54), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n869), .A2(KEYINPUT114), .A3(new_n773), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n825), .A2(KEYINPUT54), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n392), .B(KEYINPUT57), .Z(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n382), .A2(new_n390), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n738), .B(KEYINPUT115), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n870), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n865), .B1(new_n886), .B2(new_n888), .ZN(G54));
  NAND3_X1  g703(.A1(new_n870), .A2(KEYINPUT58), .A3(G475), .ZN(new_n890));
  INV_X1    g704(.A(new_n257), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n865), .ZN(G60));
  NAND2_X1  g708(.A1(G478), .A2(G902), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT59), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n814), .B2(new_n826), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n584), .A3(new_n582), .ZN(new_n898));
  INV_X1    g712(.A(new_n584), .ZN(new_n899));
  INV_X1    g713(.A(new_n582), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n882), .B(new_n896), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n898), .A2(new_n901), .A3(new_n866), .ZN(G63));
  NOR2_X1   g716(.A1(new_n627), .A2(new_n628), .ZN(new_n903));
  NAND2_X1  g717(.A1(G217), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT117), .Z(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT60), .Z(new_n906));
  NAND4_X1  g720(.A1(new_n820), .A2(KEYINPUT53), .A3(new_n822), .A4(new_n821), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n784), .B2(new_n783), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT53), .B1(new_n808), .B2(new_n812), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n903), .B(new_n906), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT118), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n825), .A2(new_n912), .A3(new_n903), .A4(new_n906), .ZN(new_n913));
  INV_X1    g727(.A(new_n906), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n563), .B1(new_n869), .B2(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n911), .A2(new_n866), .A3(new_n913), .A4(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n916), .A2(KEYINPUT116), .A3(KEYINPUT61), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT61), .B1(new_n916), .B2(KEYINPUT116), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(G66));
  INV_X1    g733(.A(G224), .ZN(new_n920));
  OAI21_X1  g734(.A(G953), .B1(new_n315), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n800), .B(KEYINPUT119), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(G953), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n873), .B1(G898), .B2(new_n216), .ZN(new_n924));
  XNOR2_X1  g738(.A(KEYINPUT120), .B(KEYINPUT121), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n923), .B(new_n926), .ZN(G69));
  AOI21_X1  g741(.A(new_n216), .B1(G227), .B2(G900), .ZN(new_n928));
  INV_X1    g742(.A(new_n764), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n774), .A2(new_n711), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT124), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n770), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n731), .A2(KEYINPUT125), .A3(new_n733), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT125), .B1(new_n731), .B2(new_n733), .ZN(new_n934));
  INV_X1    g748(.A(new_n567), .ZN(new_n935));
  NOR4_X1   g749(.A1(new_n745), .A2(new_n935), .A3(new_n666), .A4(new_n788), .ZN(new_n936));
  NOR4_X1   g750(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n930), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n764), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n931), .A2(new_n937), .A3(new_n216), .A4(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n478), .A2(new_n482), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n200), .A2(new_n205), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(G900), .A2(G953), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n671), .B2(new_n930), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n670), .A2(new_n669), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n938), .B(KEYINPUT62), .C1(new_n952), .C2(new_n664), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n796), .A2(new_n797), .ZN(new_n955));
  NOR4_X1   g769(.A1(new_n955), .A2(new_n935), .A3(new_n666), .A4(new_n803), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n830), .B2(new_n766), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n954), .A2(new_n957), .A3(new_n764), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT122), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n954), .A2(new_n957), .A3(KEYINPUT122), .A4(new_n764), .ZN(new_n961));
  AOI21_X1  g775(.A(G953), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n944), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n928), .B1(new_n949), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(KEYINPUT123), .B1(new_n941), .B2(new_n946), .ZN(new_n965));
  INV_X1    g779(.A(new_n928), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n965), .B(new_n966), .C1(new_n944), .C2(new_n962), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(G72));
  NAND4_X1  g782(.A1(new_n931), .A2(new_n937), .A3(new_n922), .A4(new_n940), .ZN(new_n969));
  XNOR2_X1  g783(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n970));
  NAND2_X1  g784(.A1(G472), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AOI211_X1 g786(.A(new_n497), .B(new_n488), .C1(new_n969), .C2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n656), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n960), .A2(new_n922), .A3(new_n961), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n972), .ZN(new_n976));
  AND2_X1   g790(.A1(new_n811), .A2(new_n813), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n499), .A2(new_n518), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n972), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n866), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n973), .A2(new_n976), .A3(new_n980), .ZN(G57));
endmodule


