

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780;

  INV_X1 U374 ( .A(G472), .ZN(n378) );
  XNOR2_X1 U375 ( .A(G113), .B(G143), .ZN(n553) );
  XNOR2_X1 U376 ( .A(G134), .B(G122), .ZN(n535) );
  XNOR2_X1 U377 ( .A(n531), .B(n530), .ZN(n426) );
  XNOR2_X2 U378 ( .A(n556), .B(n555), .ZN(n579) );
  NOR2_X2 U379 ( .A1(n688), .A2(n613), .ZN(n614) );
  AND2_X1 U380 ( .A1(n606), .A2(n620), .ZN(n607) );
  XNOR2_X2 U381 ( .A(n487), .B(n486), .ZN(n653) );
  XNOR2_X2 U382 ( .A(KEYINPUT90), .B(n654), .ZN(n752) );
  XOR2_X1 U383 ( .A(G104), .B(G107), .Z(n501) );
  XNOR2_X1 U384 ( .A(G119), .B(G116), .ZN(n522) );
  XOR2_X1 U385 ( .A(KEYINPUT11), .B(G140), .Z(n554) );
  INV_X1 U386 ( .A(G953), .ZN(n494) );
  INV_X2 U387 ( .A(KEYINPUT64), .ZN(n443) );
  BUF_X1 U388 ( .A(n436), .Z(n435) );
  BUF_X1 U389 ( .A(G110), .Z(n377) );
  NAND2_X2 U390 ( .A1(n422), .A2(n421), .ZN(n437) );
  NOR2_X2 U391 ( .A1(n433), .A2(n648), .ZN(n649) );
  NOR2_X1 U392 ( .A1(n655), .A2(n752), .ZN(n656) );
  NOR2_X1 U393 ( .A1(n668), .A2(n752), .ZN(n671) );
  AND2_X1 U394 ( .A1(n355), .A2(n488), .ZN(n354) );
  INV_X1 U395 ( .A(G134), .ZN(n499) );
  INV_X1 U396 ( .A(G119), .ZN(n367) );
  INV_X1 U397 ( .A(G110), .ZN(n368) );
  NOR2_X1 U398 ( .A1(n675), .A2(n752), .ZN(n677) );
  NAND2_X1 U399 ( .A1(n354), .A2(n353), .ZN(n352) );
  NAND2_X1 U400 ( .A1(n734), .A2(n466), .ZN(n353) );
  XNOR2_X1 U401 ( .A(n356), .B(n440), .ZN(n646) );
  NAND2_X1 U402 ( .A1(n438), .A2(n439), .ZN(n356) );
  NOR2_X1 U403 ( .A1(KEYINPUT44), .A2(n588), .ZN(n589) );
  NAND2_X1 U404 ( .A1(n461), .A2(n460), .ZN(n459) );
  NOR2_X1 U405 ( .A1(n585), .A2(KEYINPUT85), .ZN(n395) );
  NOR2_X1 U406 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U407 ( .A1(n780), .A2(n775), .ZN(n636) );
  AND2_X1 U408 ( .A1(n402), .A2(n429), .ZN(n701) );
  NOR2_X1 U409 ( .A1(n582), .A2(n565), .ZN(n567) );
  XNOR2_X1 U410 ( .A(n468), .B(n467), .ZN(n775) );
  NOR2_X1 U411 ( .A1(n739), .A2(n365), .ZN(n425) );
  XNOR2_X1 U412 ( .A(n572), .B(n449), .ZN(n699) );
  NOR2_X1 U413 ( .A1(n632), .A2(n641), .ZN(n601) );
  OR2_X1 U414 ( .A1(n698), .A2(n696), .ZN(n612) );
  NOR2_X1 U415 ( .A1(G902), .A2(n657), .ZN(n506) );
  XNOR2_X1 U416 ( .A(n410), .B(n407), .ZN(n746) );
  XNOR2_X1 U417 ( .A(n541), .B(n539), .ZN(n410) );
  INV_X1 U418 ( .A(n709), .ZN(n351) );
  NAND2_X1 U419 ( .A1(n369), .A2(n370), .ZN(n511) );
  XNOR2_X1 U420 ( .A(n409), .B(n408), .ZN(n407) );
  XNOR2_X1 U421 ( .A(n517), .B(n416), .ZN(n551) );
  NAND2_X1 U422 ( .A1(G119), .A2(n368), .ZN(n369) );
  NAND2_X1 U423 ( .A1(n367), .A2(G110), .ZN(n370) );
  XNOR2_X1 U424 ( .A(n535), .B(n533), .ZN(n408) );
  XNOR2_X1 U425 ( .A(G128), .B(KEYINPUT93), .ZN(n512) );
  XNOR2_X2 U426 ( .A(G143), .B(G128), .ZN(n481) );
  XNOR2_X2 U427 ( .A(G146), .B(G125), .ZN(n516) );
  XOR2_X2 U428 ( .A(KEYINPUT5), .B(G137), .Z(n523) );
  INV_X4 U429 ( .A(G122), .ZN(n444) );
  XOR2_X2 U430 ( .A(G137), .B(G140), .Z(n518) );
  XNOR2_X1 U431 ( .A(KEYINPUT110), .B(KEYINPUT30), .ZN(n596) );
  XNOR2_X2 U432 ( .A(n352), .B(n463), .ZN(n651) );
  NAND2_X1 U433 ( .A1(n646), .A2(n466), .ZN(n355) );
  XNOR2_X1 U434 ( .A(n361), .B(n360), .ZN(n734) );
  NAND2_X1 U435 ( .A1(n606), .A2(n718), .ZN(n597) );
  XNOR2_X2 U436 ( .A(n379), .B(n378), .ZN(n606) );
  NAND2_X1 U437 ( .A1(n599), .A2(n600), .ZN(n632) );
  XNOR2_X2 U438 ( .A(n459), .B(n458), .ZN(n414) );
  NOR2_X1 U439 ( .A1(n426), .A2(n390), .ZN(n532) );
  OR2_X2 U440 ( .A1(n390), .A2(n357), .ZN(n562) );
  NAND2_X1 U441 ( .A1(n561), .A2(n351), .ZN(n357) );
  XNOR2_X1 U442 ( .A(n442), .B(n389), .ZN(n390) );
  XNOR2_X1 U443 ( .A(n606), .B(n384), .ZN(n358) );
  XNOR2_X1 U444 ( .A(n606), .B(n384), .ZN(n619) );
  BUF_X1 U445 ( .A(n552), .Z(n359) );
  INV_X1 U446 ( .A(KEYINPUT81), .ZN(n360) );
  NAND2_X1 U447 ( .A1(n414), .A2(n388), .ZN(n361) );
  BUF_X1 U448 ( .A(n489), .Z(n362) );
  NOR2_X2 U449 ( .A1(n651), .A2(n738), .ZN(n363) );
  NOR2_X2 U450 ( .A1(n651), .A2(n738), .ZN(n364) );
  BUF_X1 U451 ( .A(n426), .Z(n365) );
  NOR2_X1 U452 ( .A1(n651), .A2(n738), .ZN(n744) );
  BUF_X1 U453 ( .A(n765), .Z(n366) );
  BUF_X1 U454 ( .A(n750), .Z(n371) );
  NAND2_X1 U455 ( .A1(n374), .A2(n372), .ZN(n588) );
  AND2_X1 U456 ( .A1(n687), .A2(n373), .ZN(n372) );
  INV_X1 U457 ( .A(n777), .ZN(n373) );
  BUF_X1 U458 ( .A(n779), .Z(n374) );
  XNOR2_X1 U459 ( .A(n567), .B(n566), .ZN(n779) );
  XNOR2_X1 U460 ( .A(n765), .B(G146), .ZN(n375) );
  XNOR2_X1 U461 ( .A(n765), .B(G146), .ZN(n529) );
  NOR2_X1 U462 ( .A1(n705), .A2(n573), .ZN(n600) );
  BUF_X1 U463 ( .A(n622), .Z(n376) );
  AND2_X1 U464 ( .A1(n621), .A2(n620), .ZN(n637) );
  NAND2_X1 U465 ( .A1(n611), .A2(n498), .ZN(n442) );
  XNOR2_X1 U466 ( .A(n441), .B(n485), .ZN(n489) );
  NOR2_X2 U467 ( .A1(n604), .A2(n709), .ZN(n473) );
  NOR2_X1 U468 ( .A1(n390), .A2(n714), .ZN(n572) );
  NOR2_X1 U469 ( .A1(n672), .A2(G902), .ZN(n379) );
  XNOR2_X1 U470 ( .A(n431), .B(n764), .ZN(n750) );
  AND2_X2 U471 ( .A1(n451), .A2(n387), .ZN(n424) );
  BUF_X1 U472 ( .A(n646), .Z(n757) );
  INV_X1 U473 ( .A(KEYINPUT71), .ZN(n462) );
  INV_X1 U474 ( .A(KEYINPUT48), .ZN(n458) );
  XNOR2_X1 U475 ( .A(n491), .B(KEYINPUT91), .ZN(n492) );
  INV_X1 U476 ( .A(KEYINPUT45), .ZN(n440) );
  INV_X1 U477 ( .A(KEYINPUT10), .ZN(n416) );
  NAND2_X2 U478 ( .A1(n424), .A2(n455), .ZN(n622) );
  INV_X1 U479 ( .A(n718), .ZN(n456) );
  XOR2_X1 U480 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n513) );
  INV_X1 U481 ( .A(KEYINPUT8), .ZN(n471) );
  INV_X1 U482 ( .A(KEYINPUT65), .ZN(n463) );
  INV_X1 U483 ( .A(KEYINPUT113), .ZN(n465) );
  INV_X1 U484 ( .A(n376), .ZN(n464) );
  OR2_X2 U485 ( .A1(n750), .A2(G902), .ZN(n406) );
  NAND2_X1 U486 ( .A1(n400), .A2(n678), .ZN(n585) );
  NAND2_X1 U487 ( .A1(n381), .A2(n401), .ZN(n400) );
  NOR2_X1 U488 ( .A1(G902), .A2(G237), .ZN(n490) );
  NOR2_X1 U489 ( .A1(G953), .A2(G237), .ZN(n546) );
  NAND2_X1 U490 ( .A1(n481), .A2(KEYINPUT4), .ZN(n421) );
  NAND2_X1 U491 ( .A1(n537), .A2(n480), .ZN(n422) );
  INV_X1 U492 ( .A(KEYINPUT4), .ZN(n480) );
  INV_X1 U493 ( .A(n776), .ZN(n434) );
  NAND2_X1 U494 ( .A1(n457), .A2(n488), .ZN(n454) );
  NAND2_X1 U495 ( .A1(n492), .A2(n453), .ZN(n452) );
  INV_X1 U496 ( .A(n488), .ZN(n453) );
  INV_X1 U497 ( .A(n608), .ZN(n573) );
  AND2_X1 U498 ( .A1(n604), .A2(n386), .ZN(n620) );
  INV_X1 U499 ( .A(n605), .ZN(n405) );
  XNOR2_X1 U500 ( .A(n534), .B(n536), .ZN(n409) );
  XNOR2_X1 U501 ( .A(n474), .B(n551), .ZN(n415) );
  XNOR2_X1 U502 ( .A(n500), .B(n501), .ZN(n503) );
  BUF_X1 U503 ( .A(n734), .Z(n769) );
  NAND2_X1 U504 ( .A1(G234), .A2(G237), .ZN(n496) );
  NAND2_X1 U505 ( .A1(n430), .A2(n429), .ZN(n714) );
  XNOR2_X1 U506 ( .A(n432), .B(n515), .ZN(n431) );
  NAND2_X1 U507 ( .A1(n540), .A2(G221), .ZN(n432) );
  XNOR2_X1 U508 ( .A(KEYINPUT42), .B(KEYINPUT112), .ZN(n467) );
  XNOR2_X1 U509 ( .A(n470), .B(n469), .ZN(n780) );
  INV_X1 U510 ( .A(KEYINPUT40), .ZN(n469) );
  XNOR2_X1 U511 ( .A(n403), .B(n624), .ZN(n402) );
  XNOR2_X1 U512 ( .A(n623), .B(KEYINPUT114), .ZN(n624) );
  INV_X1 U513 ( .A(n398), .ZN(n761) );
  AND2_X1 U514 ( .A1(n699), .A2(KEYINPUT97), .ZN(n380) );
  AND2_X1 U515 ( .A1(n446), .A2(n427), .ZN(n381) );
  XOR2_X1 U516 ( .A(KEYINPUT72), .B(G469), .Z(n382) );
  XOR2_X1 U517 ( .A(n510), .B(n509), .Z(n383) );
  XNOR2_X1 U518 ( .A(KEYINPUT6), .B(KEYINPUT106), .ZN(n384) );
  AND2_X1 U519 ( .A1(n451), .A2(n454), .ZN(n385) );
  AND2_X1 U520 ( .A1(n351), .A2(n405), .ZN(n386) );
  NOR2_X1 U521 ( .A1(n450), .A2(n456), .ZN(n387) );
  AND2_X1 U522 ( .A1(n434), .A2(n703), .ZN(n388) );
  XOR2_X1 U523 ( .A(KEYINPUT89), .B(KEYINPUT0), .Z(n389) );
  INV_X1 U524 ( .A(KEYINPUT97), .ZN(n448) );
  INV_X1 U525 ( .A(n612), .ZN(n428) );
  XNOR2_X1 U526 ( .A(G902), .B(KEYINPUT15), .ZN(n645) );
  NOR2_X1 U527 ( .A1(n577), .A2(n391), .ZN(n578) );
  XNOR2_X1 U528 ( .A(n442), .B(n389), .ZN(n575) );
  OR2_X2 U529 ( .A1(n619), .A2(n705), .ZN(n413) );
  NOR2_X2 U530 ( .A1(n413), .A2(n704), .ZN(n531) );
  INV_X1 U531 ( .A(n412), .ZN(n391) );
  XNOR2_X1 U532 ( .A(n578), .B(KEYINPUT96), .ZN(n679) );
  NAND2_X1 U533 ( .A1(n569), .A2(n412), .ZN(n687) );
  NAND2_X1 U534 ( .A1(n707), .A2(n412), .ZN(n712) );
  NAND2_X1 U535 ( .A1(n392), .A2(KEYINPUT85), .ZN(n396) );
  NAND2_X1 U536 ( .A1(n397), .A2(n393), .ZN(n392) );
  INV_X1 U537 ( .A(n585), .ZN(n393) );
  AND2_X2 U538 ( .A1(n571), .A2(n570), .ZN(n397) );
  NAND2_X1 U539 ( .A1(n396), .A2(n394), .ZN(n438) );
  NAND2_X1 U540 ( .A1(n397), .A2(n395), .ZN(n394) );
  OR2_X1 U541 ( .A1(n399), .A2(n760), .ZN(n398) );
  XNOR2_X1 U542 ( .A(n399), .B(n437), .ZN(n441) );
  XNOR2_X1 U543 ( .A(n479), .B(n478), .ZN(n399) );
  OR2_X1 U544 ( .A1(n679), .A2(n447), .ZN(n401) );
  NAND2_X1 U545 ( .A1(n404), .A2(n464), .ZN(n403) );
  XNOR2_X1 U546 ( .A(n637), .B(n465), .ZN(n404) );
  XNOR2_X2 U547 ( .A(n406), .B(n383), .ZN(n604) );
  XNOR2_X2 U548 ( .A(n411), .B(KEYINPUT69), .ZN(n543) );
  XNOR2_X2 U549 ( .A(G131), .B(KEYINPUT70), .ZN(n411) );
  XNOR2_X2 U550 ( .A(n543), .B(n499), .ZN(n423) );
  NOR2_X1 U551 ( .A1(n705), .A2(n412), .ZN(n430) );
  INV_X1 U552 ( .A(n606), .ZN(n412) );
  XNOR2_X1 U553 ( .A(n636), .B(KEYINPUT46), .ZN(n460) );
  XNOR2_X2 U554 ( .A(n622), .B(KEYINPUT19), .ZN(n611) );
  XNOR2_X2 U555 ( .A(KEYINPUT73), .B(KEYINPUT3), .ZN(n475) );
  NAND2_X1 U556 ( .A1(n414), .A2(n703), .ZN(n433) );
  NOR2_X1 U557 ( .A1(n722), .A2(n428), .ZN(n723) );
  XNOR2_X1 U558 ( .A(n417), .B(n415), .ZN(n665) );
  XNOR2_X1 U559 ( .A(n419), .B(n418), .ZN(n417) );
  XNOR2_X1 U560 ( .A(n548), .B(n547), .ZN(n418) );
  XNOR2_X1 U561 ( .A(n549), .B(n420), .ZN(n419) );
  XNOR2_X1 U562 ( .A(n359), .B(n550), .ZN(n420) );
  XNOR2_X2 U563 ( .A(n423), .B(n437), .ZN(n765) );
  NOR2_X1 U564 ( .A1(n725), .A2(n365), .ZN(n726) );
  NOR2_X1 U565 ( .A1(n380), .A2(n428), .ZN(n427) );
  INV_X1 U566 ( .A(n704), .ZN(n429) );
  XNOR2_X2 U567 ( .A(n608), .B(n507), .ZN(n704) );
  XNOR2_X2 U568 ( .A(n506), .B(n382), .ZN(n608) );
  NAND2_X1 U569 ( .A1(n436), .A2(G234), .ZN(n472) );
  XNOR2_X2 U570 ( .A(n443), .B(G953), .ZN(n436) );
  NAND2_X1 U571 ( .A1(n436), .A2(G227), .ZN(n500) );
  NAND2_X1 U572 ( .A1(n435), .A2(G224), .ZN(n483) );
  NOR2_X1 U573 ( .A1(n435), .A2(G900), .ZN(n591) );
  NOR2_X1 U574 ( .A1(n435), .A2(G952), .ZN(n654) );
  NAND2_X1 U575 ( .A1(n772), .A2(n435), .ZN(n773) );
  INV_X1 U576 ( .A(n589), .ZN(n439) );
  INV_X1 U577 ( .A(KEYINPUT2), .ZN(n466) );
  NOR2_X2 U578 ( .A1(n757), .A2(n650), .ZN(n738) );
  XNOR2_X1 U579 ( .A(n597), .B(n596), .ZN(n598) );
  XNOR2_X2 U580 ( .A(n562), .B(KEYINPUT22), .ZN(n582) );
  XNOR2_X1 U581 ( .A(n375), .B(n505), .ZN(n657) );
  XNOR2_X1 U582 ( .A(n628), .B(n462), .ZN(n461) );
  XNOR2_X2 U583 ( .A(n444), .B(G104), .ZN(n552) );
  NAND2_X1 U584 ( .A1(n445), .A2(n448), .ZN(n447) );
  INV_X1 U585 ( .A(n699), .ZN(n445) );
  NAND2_X1 U586 ( .A1(n679), .A2(KEYINPUT97), .ZN(n446) );
  INV_X1 U587 ( .A(KEYINPUT31), .ZN(n449) );
  NAND2_X1 U588 ( .A1(n455), .A2(n385), .ZN(n641) );
  INV_X1 U589 ( .A(n454), .ZN(n450) );
  OR2_X2 U590 ( .A1(n489), .A2(n452), .ZN(n451) );
  NAND2_X1 U591 ( .A1(n489), .A2(n457), .ZN(n455) );
  INV_X1 U592 ( .A(n492), .ZN(n457) );
  XNOR2_X1 U593 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U594 ( .A(n504), .B(G101), .ZN(n505) );
  NOR2_X1 U595 ( .A1(n739), .A2(n629), .ZN(n468) );
  NAND2_X1 U596 ( .A1(n643), .A2(n696), .ZN(n470) );
  XNOR2_X1 U597 ( .A(n635), .B(n634), .ZN(n643) );
  XNOR2_X2 U598 ( .A(n472), .B(n471), .ZN(n540) );
  XNOR2_X2 U599 ( .A(n473), .B(KEYINPUT67), .ZN(n705) );
  XNOR2_X1 U600 ( .A(n641), .B(KEYINPUT38), .ZN(n719) );
  BUF_X1 U601 ( .A(n364), .Z(n748) );
  XNOR2_X2 U602 ( .A(n476), .B(n475), .ZN(n525) );
  XOR2_X2 U603 ( .A(G101), .B(G113), .Z(n476) );
  XOR2_X2 U604 ( .A(G116), .B(G107), .Z(n538) );
  XOR2_X1 U605 ( .A(n554), .B(n553), .Z(n474) );
  INV_X1 U606 ( .A(KEYINPUT74), .ZN(n616) );
  XNOR2_X1 U607 ( .A(n617), .B(n616), .ZN(n627) );
  AND2_X1 U608 ( .A1(n497), .A2(n729), .ZN(n498) );
  XNOR2_X1 U609 ( .A(n484), .B(n483), .ZN(n485) );
  INV_X1 U610 ( .A(KEYINPUT36), .ZN(n623) );
  XNOR2_X1 U611 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U612 ( .A(n633), .B(KEYINPUT39), .ZN(n634) );
  INV_X1 U613 ( .A(n752), .ZN(n662) );
  BUF_X1 U614 ( .A(n586), .Z(n777) );
  XOR2_X1 U615 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n487) );
  XNOR2_X1 U616 ( .A(n538), .B(n552), .ZN(n477) );
  XNOR2_X1 U617 ( .A(n477), .B(n525), .ZN(n479) );
  XOR2_X1 U618 ( .A(n511), .B(KEYINPUT16), .Z(n478) );
  INV_X1 U619 ( .A(n481), .ZN(n537) );
  XOR2_X1 U620 ( .A(n516), .B(KEYINPUT18), .Z(n482) );
  XOR2_X1 U621 ( .A(n482), .B(KEYINPUT17), .Z(n484) );
  XNOR2_X1 U622 ( .A(n362), .B(KEYINPUT88), .ZN(n486) );
  INV_X1 U623 ( .A(n645), .ZN(n488) );
  XNOR2_X1 U624 ( .A(n490), .B(KEYINPUT75), .ZN(n493) );
  NAND2_X1 U625 ( .A1(G210), .A2(n493), .ZN(n491) );
  NAND2_X1 U626 ( .A1(G214), .A2(n493), .ZN(n718) );
  XNOR2_X1 U627 ( .A(G898), .B(KEYINPUT92), .ZN(n755) );
  NOR2_X1 U628 ( .A1(n494), .A2(n755), .ZN(n760) );
  NAND2_X1 U629 ( .A1(n760), .A2(G902), .ZN(n495) );
  NAND2_X1 U630 ( .A1(G952), .A2(n494), .ZN(n593) );
  NAND2_X1 U631 ( .A1(n495), .A2(n593), .ZN(n497) );
  XNOR2_X1 U632 ( .A(KEYINPUT14), .B(n496), .ZN(n729) );
  XOR2_X1 U633 ( .A(n518), .B(n377), .Z(n502) );
  INV_X1 U634 ( .A(KEYINPUT1), .ZN(n507) );
  XOR2_X1 U635 ( .A(KEYINPUT76), .B(KEYINPUT25), .Z(n510) );
  NAND2_X1 U636 ( .A1(G234), .A2(n645), .ZN(n508) );
  XNOR2_X1 U637 ( .A(KEYINPUT20), .B(n508), .ZN(n519) );
  NAND2_X1 U638 ( .A1(n519), .A2(G217), .ZN(n509) );
  XNOR2_X1 U639 ( .A(n511), .B(n512), .ZN(n514) );
  INV_X1 U640 ( .A(n516), .ZN(n517) );
  XNOR2_X1 U641 ( .A(n551), .B(n518), .ZN(n764) );
  XOR2_X1 U642 ( .A(KEYINPUT94), .B(KEYINPUT21), .Z(n521) );
  NAND2_X1 U643 ( .A1(n519), .A2(G221), .ZN(n520) );
  XOR2_X1 U644 ( .A(n521), .B(n520), .Z(n709) );
  XNOR2_X1 U645 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U646 ( .A(n525), .B(n524), .Z(n527) );
  NAND2_X1 U647 ( .A1(n546), .A2(G210), .ZN(n526) );
  XNOR2_X1 U648 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U649 ( .A(n529), .B(n528), .ZN(n672) );
  XNOR2_X1 U650 ( .A(KEYINPUT108), .B(KEYINPUT33), .ZN(n530) );
  XNOR2_X1 U651 ( .A(n532), .B(KEYINPUT34), .ZN(n557) );
  XOR2_X1 U652 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n534) );
  XNOR2_X1 U653 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n533) );
  XOR2_X1 U654 ( .A(KEYINPUT102), .B(KEYINPUT105), .Z(n536) );
  XOR2_X1 U655 ( .A(n538), .B(n481), .Z(n539) );
  NAND2_X1 U656 ( .A1(n540), .A2(G217), .ZN(n541) );
  NOR2_X1 U657 ( .A1(G902), .A2(n746), .ZN(n542) );
  XOR2_X1 U658 ( .A(G478), .B(n542), .Z(n580) );
  INV_X1 U659 ( .A(n580), .ZN(n560) );
  XOR2_X1 U660 ( .A(KEYINPUT13), .B(G475), .Z(n556) );
  INV_X1 U661 ( .A(n543), .ZN(n549) );
  XOR2_X1 U662 ( .A(KEYINPUT100), .B(KEYINPUT98), .Z(n545) );
  XNOR2_X1 U663 ( .A(KEYINPUT12), .B(KEYINPUT99), .ZN(n544) );
  XNOR2_X1 U664 ( .A(n545), .B(n544), .ZN(n548) );
  NAND2_X1 U665 ( .A1(G214), .A2(n546), .ZN(n547) );
  INV_X1 U666 ( .A(KEYINPUT101), .ZN(n550) );
  NOR2_X1 U667 ( .A1(G902), .A2(n665), .ZN(n555) );
  NOR2_X1 U668 ( .A1(n560), .A2(n579), .ZN(n590) );
  NAND2_X1 U669 ( .A1(n557), .A2(n590), .ZN(n558) );
  XNOR2_X1 U670 ( .A(n558), .B(KEYINPUT35), .ZN(n586) );
  NAND2_X1 U671 ( .A1(n586), .A2(KEYINPUT44), .ZN(n559) );
  XNOR2_X1 U672 ( .A(n559), .B(KEYINPUT86), .ZN(n571) );
  NAND2_X1 U673 ( .A1(n560), .A2(n579), .ZN(n721) );
  INV_X1 U674 ( .A(n721), .ZN(n561) );
  INV_X1 U675 ( .A(n358), .ZN(n581) );
  XOR2_X1 U676 ( .A(n604), .B(KEYINPUT107), .Z(n708) );
  INV_X1 U677 ( .A(n708), .ZN(n563) );
  OR2_X1 U678 ( .A1(n581), .A2(n563), .ZN(n564) );
  OR2_X1 U679 ( .A1(n704), .A2(n564), .ZN(n565) );
  XNOR2_X1 U680 ( .A(KEYINPUT32), .B(KEYINPUT77), .ZN(n566) );
  NAND2_X1 U681 ( .A1(n604), .A2(n704), .ZN(n568) );
  NOR2_X1 U682 ( .A1(n582), .A2(n568), .ZN(n569) );
  NAND2_X1 U683 ( .A1(n779), .A2(n687), .ZN(n587) );
  NAND2_X1 U684 ( .A1(n587), .A2(KEYINPUT44), .ZN(n570) );
  INV_X1 U685 ( .A(n600), .ZN(n574) );
  NOR2_X1 U686 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U687 ( .A(n576), .B(KEYINPUT95), .ZN(n577) );
  NOR2_X1 U688 ( .A1(n579), .A2(n580), .ZN(n618) );
  BUF_X1 U689 ( .A(n618), .Z(n696) );
  NAND2_X1 U690 ( .A1(n580), .A2(n579), .ZN(n689) );
  INV_X1 U691 ( .A(n689), .ZN(n698) );
  NOR2_X1 U692 ( .A1(n582), .A2(n581), .ZN(n584) );
  NOR2_X1 U693 ( .A1(n429), .A2(n708), .ZN(n583) );
  NAND2_X1 U694 ( .A1(n584), .A2(n583), .ZN(n678) );
  INV_X1 U695 ( .A(n590), .ZN(n603) );
  NAND2_X1 U696 ( .A1(G902), .A2(n591), .ZN(n592) );
  NAND2_X1 U697 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U698 ( .A1(n594), .A2(n729), .ZN(n595) );
  XNOR2_X1 U699 ( .A(KEYINPUT78), .B(n595), .ZN(n605) );
  NOR2_X1 U700 ( .A1(n605), .A2(n598), .ZN(n599) );
  XNOR2_X1 U701 ( .A(n601), .B(KEYINPUT111), .ZN(n602) );
  NOR2_X1 U702 ( .A1(n603), .A2(n602), .ZN(n692) );
  XNOR2_X1 U703 ( .A(n607), .B(KEYINPUT28), .ZN(n609) );
  NAND2_X1 U704 ( .A1(n609), .A2(n608), .ZN(n629) );
  INV_X1 U705 ( .A(n629), .ZN(n610) );
  NAND2_X1 U706 ( .A1(n611), .A2(n610), .ZN(n688) );
  NAND2_X1 U707 ( .A1(KEYINPUT68), .A2(n612), .ZN(n613) );
  XOR2_X1 U708 ( .A(KEYINPUT47), .B(n614), .Z(n615) );
  NOR2_X1 U709 ( .A1(n692), .A2(n615), .ZN(n617) );
  INV_X1 U710 ( .A(n618), .ZN(n693) );
  NOR2_X1 U711 ( .A1(n358), .A2(n693), .ZN(n621) );
  INV_X1 U712 ( .A(KEYINPUT83), .ZN(n625) );
  XNOR2_X1 U713 ( .A(n701), .B(n625), .ZN(n626) );
  NAND2_X1 U714 ( .A1(n719), .A2(n718), .ZN(n722) );
  NOR2_X1 U715 ( .A1(n722), .A2(n721), .ZN(n630) );
  XNOR2_X1 U716 ( .A(n630), .B(KEYINPUT41), .ZN(n739) );
  INV_X1 U717 ( .A(n719), .ZN(n631) );
  NOR2_X1 U718 ( .A1(n632), .A2(n631), .ZN(n635) );
  INV_X1 U719 ( .A(KEYINPUT84), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n637), .A2(n718), .ZN(n638) );
  XNOR2_X1 U721 ( .A(n638), .B(KEYINPUT109), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n639), .A2(n704), .ZN(n640) );
  XNOR2_X1 U723 ( .A(n640), .B(KEYINPUT43), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n703) );
  NAND2_X1 U725 ( .A1(n643), .A2(n698), .ZN(n644) );
  XNOR2_X1 U726 ( .A(KEYINPUT115), .B(n644), .ZN(n776) );
  OR2_X1 U727 ( .A1(n466), .A2(n776), .ZN(n647) );
  XOR2_X1 U728 ( .A(KEYINPUT79), .B(n647), .Z(n648) );
  XOR2_X1 U729 ( .A(KEYINPUT82), .B(n649), .Z(n650) );
  NAND2_X1 U730 ( .A1(n363), .A2(G210), .ZN(n652) );
  XNOR2_X1 U731 ( .A(n652), .B(n653), .ZN(n655) );
  XNOR2_X1 U732 ( .A(n656), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U733 ( .A1(n363), .A2(G469), .ZN(n661) );
  XNOR2_X1 U734 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n657), .B(KEYINPUT57), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n661), .B(n660), .ZN(n663) );
  NAND2_X1 U738 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U739 ( .A(n664), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U740 ( .A1(n744), .A2(G475), .ZN(n667) );
  XOR2_X1 U741 ( .A(n665), .B(KEYINPUT59), .Z(n666) );
  XNOR2_X1 U742 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U743 ( .A(KEYINPUT66), .B(KEYINPUT122), .ZN(n669) );
  XNOR2_X1 U744 ( .A(n669), .B(KEYINPUT60), .ZN(n670) );
  XNOR2_X1 U745 ( .A(n671), .B(n670), .ZN(G60) );
  XNOR2_X1 U746 ( .A(n672), .B(KEYINPUT62), .ZN(n674) );
  NAND2_X1 U747 ( .A1(n364), .A2(G472), .ZN(n673) );
  XNOR2_X1 U748 ( .A(n673), .B(n674), .ZN(n675) );
  XNOR2_X1 U749 ( .A(KEYINPUT63), .B(KEYINPUT87), .ZN(n676) );
  XNOR2_X1 U750 ( .A(n677), .B(n676), .ZN(G57) );
  XNOR2_X1 U751 ( .A(G101), .B(n678), .ZN(G3) );
  XNOR2_X1 U752 ( .A(G104), .B(KEYINPUT116), .ZN(n681) );
  BUF_X1 U753 ( .A(n679), .Z(n682) );
  NAND2_X1 U754 ( .A1(n696), .A2(n682), .ZN(n680) );
  XNOR2_X1 U755 ( .A(n681), .B(n680), .ZN(G6) );
  XOR2_X1 U756 ( .A(KEYINPUT26), .B(KEYINPUT117), .Z(n684) );
  NAND2_X1 U757 ( .A1(n698), .A2(n682), .ZN(n683) );
  XNOR2_X1 U758 ( .A(n684), .B(n683), .ZN(n686) );
  XOR2_X1 U759 ( .A(G107), .B(KEYINPUT27), .Z(n685) );
  XNOR2_X1 U760 ( .A(n686), .B(n685), .ZN(G9) );
  XNOR2_X1 U761 ( .A(n377), .B(n687), .ZN(G12) );
  NOR2_X1 U762 ( .A1(n689), .A2(n688), .ZN(n691) );
  XNOR2_X1 U763 ( .A(G128), .B(KEYINPUT29), .ZN(n690) );
  XNOR2_X1 U764 ( .A(n691), .B(n690), .ZN(G30) );
  XOR2_X1 U765 ( .A(n692), .B(G143), .Z(G45) );
  NOR2_X1 U766 ( .A1(n693), .A2(n688), .ZN(n694) );
  XOR2_X1 U767 ( .A(KEYINPUT118), .B(n694), .Z(n695) );
  XNOR2_X1 U768 ( .A(G146), .B(n695), .ZN(G48) );
  NAND2_X1 U769 ( .A1(n699), .A2(n696), .ZN(n697) );
  XNOR2_X1 U770 ( .A(n697), .B(G113), .ZN(G15) );
  NAND2_X1 U771 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U772 ( .A(n700), .B(G116), .ZN(G18) );
  XNOR2_X1 U773 ( .A(G125), .B(n701), .ZN(n702) );
  XNOR2_X1 U774 ( .A(n702), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U775 ( .A(G140), .B(n703), .ZN(G42) );
  NAND2_X1 U776 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U777 ( .A(n706), .B(KEYINPUT50), .ZN(n707) );
  NAND2_X1 U778 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U779 ( .A(KEYINPUT49), .B(n710), .ZN(n711) );
  NOR2_X1 U780 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U781 ( .A(n713), .B(KEYINPUT119), .ZN(n715) );
  NAND2_X1 U782 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U783 ( .A(KEYINPUT51), .B(n716), .ZN(n717) );
  NOR2_X1 U784 ( .A1(n739), .A2(n717), .ZN(n727) );
  NOR2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U786 ( .A1(n721), .A2(n720), .ZN(n724) );
  NOR2_X1 U787 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U788 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U789 ( .A(KEYINPUT52), .B(n728), .ZN(n731) );
  NAND2_X1 U790 ( .A1(G952), .A2(n729), .ZN(n730) );
  NOR2_X1 U791 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U792 ( .A1(G953), .A2(n732), .ZN(n742) );
  NAND2_X1 U793 ( .A1(n757), .A2(n466), .ZN(n733) );
  XNOR2_X1 U794 ( .A(n733), .B(KEYINPUT80), .ZN(n736) );
  NAND2_X1 U795 ( .A1(n769), .A2(n466), .ZN(n735) );
  NAND2_X1 U796 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U797 ( .A1(n738), .A2(n737), .ZN(n740) );
  NOR2_X1 U798 ( .A1(n740), .A2(n425), .ZN(n741) );
  NAND2_X1 U799 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U800 ( .A(KEYINPUT53), .B(n743), .Z(G75) );
  NAND2_X1 U801 ( .A1(G478), .A2(n748), .ZN(n745) );
  XNOR2_X1 U802 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U803 ( .A1(n752), .A2(n747), .ZN(G63) );
  NAND2_X1 U804 ( .A1(G217), .A2(n748), .ZN(n749) );
  XNOR2_X1 U805 ( .A(n371), .B(n749), .ZN(n751) );
  NOR2_X1 U806 ( .A1(n752), .A2(n751), .ZN(G66) );
  XOR2_X1 U807 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n754) );
  NAND2_X1 U808 ( .A1(G224), .A2(G953), .ZN(n753) );
  XNOR2_X1 U809 ( .A(n754), .B(n753), .ZN(n756) );
  NAND2_X1 U810 ( .A1(n756), .A2(n755), .ZN(n759) );
  OR2_X1 U811 ( .A1(n757), .A2(G953), .ZN(n758) );
  NAND2_X1 U812 ( .A1(n759), .A2(n758), .ZN(n763) );
  XNOR2_X1 U813 ( .A(n761), .B(KEYINPUT124), .ZN(n762) );
  XNOR2_X1 U814 ( .A(n763), .B(n762), .ZN(G69) );
  XOR2_X1 U815 ( .A(n366), .B(n764), .Z(n770) );
  XOR2_X1 U816 ( .A(G227), .B(n770), .Z(n766) );
  NAND2_X1 U817 ( .A1(n766), .A2(G900), .ZN(n767) );
  NAND2_X1 U818 ( .A1(G953), .A2(n767), .ZN(n768) );
  XNOR2_X1 U819 ( .A(n768), .B(KEYINPUT126), .ZN(n774) );
  XNOR2_X1 U820 ( .A(n769), .B(KEYINPUT125), .ZN(n771) );
  XNOR2_X1 U821 ( .A(n771), .B(n770), .ZN(n772) );
  NAND2_X1 U822 ( .A1(n774), .A2(n773), .ZN(G72) );
  XOR2_X1 U823 ( .A(G137), .B(n775), .Z(G39) );
  XOR2_X1 U824 ( .A(G134), .B(n776), .Z(G36) );
  XNOR2_X1 U825 ( .A(n777), .B(G122), .ZN(n778) );
  XNOR2_X1 U826 ( .A(n778), .B(KEYINPUT127), .ZN(G24) );
  XNOR2_X1 U827 ( .A(G119), .B(n374), .ZN(G21) );
  XOR2_X1 U828 ( .A(n780), .B(G131), .Z(G33) );
endmodule

