//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n190), .B(KEYINPUT76), .Z(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n193), .A2(new_n195), .A3(KEYINPUT16), .ZN(new_n196));
  OR3_X1    g010(.A1(new_n194), .A2(KEYINPUT16), .A3(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n197), .A3(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G128), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n205), .B(new_n207), .C1(G119), .C2(new_n206), .ZN(new_n208));
  XNOR2_X1  g022(.A(G119), .B(G128), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT24), .B(G110), .Z(new_n210));
  AOI22_X1  g024(.A1(new_n208), .A2(G110), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n202), .A2(new_n211), .ZN(new_n212));
  OAI22_X1  g026(.A1(new_n208), .A2(G110), .B1(new_n209), .B2(new_n210), .ZN(new_n213));
  XNOR2_X1  g027(.A(G125), .B(G140), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n199), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n213), .A2(new_n201), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n212), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n191), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n212), .A2(new_n216), .A3(new_n190), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT25), .ZN(new_n220));
  AOI21_X1  g034(.A(G902), .B1(new_n220), .B2(KEYINPUT77), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n220), .A2(KEYINPUT77), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n223), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n218), .A2(new_n225), .A3(new_n219), .A4(new_n221), .ZN(new_n226));
  INV_X1    g040(.A(G217), .ZN(new_n227));
  INV_X1    g041(.A(G902), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(G234), .B2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n224), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n218), .A2(new_n219), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n229), .A2(G902), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n234), .B(KEYINPUT78), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G472), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT74), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT11), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(G137), .ZN(new_n241));
  INV_X1    g055(.A(G137), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT11), .A3(G134), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(G137), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G131), .ZN(new_n246));
  INV_X1    g060(.A(G131), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n241), .A2(new_n243), .A3(new_n247), .A4(new_n244), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n199), .A2(G143), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G146), .ZN(new_n252));
  AND2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT66), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n250), .A2(new_n252), .A3(new_n253), .A4(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT64), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n259), .B1(new_n251), .B2(G146), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n199), .A2(KEYINPUT64), .A3(G143), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n250), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT0), .B(G128), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT65), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n251), .A2(G146), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT64), .B1(new_n199), .B2(G143), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n259), .A2(new_n251), .A3(G146), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n269), .A2(new_n270), .A3(new_n263), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n249), .B(new_n258), .C1(new_n265), .C2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n273), .A2(new_n250), .A3(new_n252), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n206), .B1(new_n250), .B2(KEYINPUT1), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n262), .B2(new_n276), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n240), .A2(G137), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n242), .A2(G134), .ZN(new_n279));
  OAI21_X1  g093(.A(G131), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n248), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT67), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n248), .A2(new_n280), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n273), .A2(new_n250), .A3(new_n252), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n269), .B2(new_n275), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n272), .A2(new_n282), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT30), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n291));
  INV_X1    g105(.A(G116), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n292), .B2(G119), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n204), .A2(KEYINPUT68), .A3(G116), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(G119), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT2), .B(G113), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT69), .A4(new_n295), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n296), .A2(new_n299), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n283), .A2(new_n285), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT70), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT70), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n283), .A2(new_n285), .A3(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n272), .A2(new_n305), .A3(KEYINPUT30), .A4(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n290), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n272), .A2(new_n305), .A3(new_n307), .ZN(new_n310));
  INV_X1    g124(.A(new_n303), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G237), .A2(G953), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G210), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT27), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT26), .B(G101), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n238), .B1(new_n313), .B2(new_n319), .ZN(new_n320));
  AOI211_X1 g134(.A(KEYINPUT74), .B(new_n318), .C1(new_n309), .C2(new_n312), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n288), .A2(new_n303), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT71), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n326), .A2(new_n327), .B1(new_n310), .B2(new_n311), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n288), .A2(KEYINPUT71), .A3(new_n303), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n311), .A2(new_n272), .A3(new_n304), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n325), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n318), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n324), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n333), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n288), .A2(KEYINPUT71), .A3(new_n303), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT71), .B1(new_n288), .B2(new_n303), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n272), .A2(new_n305), .A3(new_n307), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(new_n303), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n336), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(KEYINPUT73), .B(new_n335), .C1(new_n340), .C2(new_n325), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n322), .A2(new_n323), .A3(new_n334), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(new_n303), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n312), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT28), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n333), .A2(new_n323), .ZN(new_n346));
  AOI21_X1  g160(.A(G902), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n237), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n332), .B1(new_n340), .B2(new_n325), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n309), .A2(new_n312), .A3(new_n318), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT31), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n309), .A2(KEYINPUT31), .A3(new_n312), .A4(new_n318), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n350), .A2(new_n319), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(G472), .A2(G902), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT72), .ZN(new_n357));
  OAI21_X1  g171(.A(KEYINPUT32), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n332), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n319), .B1(new_n330), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n354), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT32), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n348), .A2(new_n349), .B1(new_n358), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n313), .A2(new_n319), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT74), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n313), .A2(new_n238), .A3(new_n319), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n341), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n326), .A2(new_n327), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(new_n329), .A3(new_n312), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n333), .B1(new_n371), .B2(KEYINPUT28), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n323), .B1(new_n372), .B2(KEYINPUT73), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n347), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G472), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT75), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n236), .B1(new_n365), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G210), .B1(G237), .B2(G902), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT90), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT89), .ZN(new_n381));
  INV_X1    g195(.A(G104), .ZN(new_n382));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(new_n382), .B2(G107), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G104), .ZN(new_n386));
  INV_X1    g200(.A(G101), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(G107), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n383), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n382), .A2(G107), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n385), .A2(G104), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n389), .B(new_n392), .C1(new_n296), .C2(new_n299), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT5), .A4(new_n295), .ZN(new_n394));
  INV_X1    g208(.A(G113), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n292), .A2(G119), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT88), .B1(new_n393), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n389), .A2(new_n392), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT88), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n394), .A2(new_n398), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n401), .A2(new_n302), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n389), .A2(new_n392), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n397), .B1(new_n298), .B2(new_n300), .ZN(new_n407));
  INV_X1    g221(.A(new_n398), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n302), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n405), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G122), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT8), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n381), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n409), .A2(new_n406), .ZN(new_n415));
  OAI211_X1 g229(.A(KEYINPUT89), .B(new_n412), .C1(new_n415), .C2(new_n405), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n262), .A2(KEYINPUT65), .A3(new_n264), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n270), .B1(new_n269), .B2(new_n263), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n418), .A2(new_n419), .B1(new_n255), .B2(new_n257), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT86), .B1(new_n420), .B2(new_n194), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n258), .B1(new_n265), .B2(new_n271), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT86), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(G125), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n194), .B(new_n284), .C1(new_n269), .C2(new_n275), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT87), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n421), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G224), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT7), .B1(new_n428), .B2(G953), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n383), .A2(new_n386), .A3(new_n388), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT4), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(G101), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n432), .B1(new_n431), .B2(G101), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT79), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n436), .A2(new_n437), .A3(new_n389), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n437), .B1(new_n436), .B2(new_n389), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n435), .B(new_n303), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n406), .A2(KEYINPUT81), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT81), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n389), .A2(new_n392), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n444), .B(new_n302), .C1(new_n407), .C2(new_n408), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n440), .A2(new_n445), .A3(new_n411), .ZN(new_n446));
  INV_X1    g260(.A(new_n429), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n421), .A2(new_n424), .A3(new_n426), .A4(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n430), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n380), .B(new_n228), .C1(new_n417), .C2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n428), .A2(G953), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n427), .B(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n440), .A2(new_n445), .ZN(new_n453));
  INV_X1    g267(.A(new_n411), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(KEYINPUT6), .A3(new_n446), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n453), .A2(new_n457), .A3(new_n454), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n450), .A2(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n446), .A2(new_n448), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n461), .A2(new_n430), .A3(new_n414), .A4(new_n416), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n380), .B1(new_n462), .B2(new_n228), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n379), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n228), .B1(new_n417), .B2(new_n449), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT90), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n466), .A2(new_n378), .A3(new_n459), .A4(new_n450), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G214), .B1(G237), .B2(G902), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT9), .B(G234), .ZN(new_n471));
  OAI21_X1  g285(.A(G221), .B1(new_n471), .B2(G902), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n401), .A2(new_n285), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT83), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n474), .A2(new_n475), .B1(new_n246), .B2(new_n248), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT1), .B1(new_n251), .B2(G146), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n477), .A2(G128), .B1(new_n250), .B2(new_n252), .ZN(new_n478));
  OAI211_X1 g292(.A(new_n389), .B(new_n392), .C1(new_n478), .C2(new_n274), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n479), .B(KEYINPUT83), .C1(new_n285), .C2(new_n401), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT12), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n277), .A2(new_n475), .A3(new_n406), .ZN(new_n482));
  AND4_X1   g296(.A1(KEYINPUT12), .A2(new_n480), .A3(new_n249), .A4(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT84), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n435), .B(new_n420), .C1(new_n438), .C2(new_n439), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n479), .A2(KEYINPUT10), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n277), .B1(new_n441), .B2(new_n443), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT10), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n249), .B(KEYINPUT82), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n485), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G110), .B(G140), .ZN(new_n492));
  INV_X1    g306(.A(G227), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(G953), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n492), .B(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT12), .ZN(new_n497));
  INV_X1    g311(.A(new_n480), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n482), .A2(new_n249), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n476), .A2(KEYINPUT12), .A3(new_n480), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT84), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n484), .A2(new_n491), .A3(new_n496), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT85), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n491), .A2(new_n496), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT85), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n506), .A2(new_n507), .A3(new_n484), .A4(new_n503), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n485), .A2(new_n489), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n249), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n491), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n495), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n505), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G469), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n513), .A2(new_n514), .A3(new_n228), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n514), .A2(new_n228), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n491), .B1(new_n483), .B2(new_n481), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n495), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n510), .A2(new_n491), .A3(new_n496), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n516), .B1(new_n521), .B2(G469), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n473), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n471), .A2(new_n227), .A3(G953), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT95), .B1(new_n206), .B2(G143), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(new_n251), .A3(G128), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n251), .A2(G128), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n240), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(G122), .ZN(new_n534));
  INV_X1    g348(.A(G122), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n535), .A2(KEYINPUT94), .ZN(new_n536));
  OAI21_X1  g350(.A(G116), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n535), .A2(G116), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n385), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n535), .A2(KEYINPUT94), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n533), .A2(G122), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n292), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n543), .A2(G107), .A3(new_n538), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n532), .B1(new_n540), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT13), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n530), .B1(new_n529), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n526), .A2(new_n528), .A3(KEYINPUT13), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n240), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n537), .A2(new_n385), .A3(new_n539), .ZN(new_n550));
  AOI211_X1 g364(.A(G134), .B(new_n530), .C1(new_n528), .C2(new_n526), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n240), .B1(new_n529), .B2(new_n531), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT14), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n292), .A3(G122), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n538), .A2(new_n554), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n543), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n385), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  OAI22_X1  g374(.A1(new_n545), .A2(new_n549), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT97), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n551), .A2(new_n552), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n537), .B1(new_n554), .B2(new_n538), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n555), .B(KEYINPUT96), .ZN(new_n566));
  OAI21_X1  g380(.A(G107), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n564), .A2(new_n567), .A3(new_n550), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n547), .A2(new_n548), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G134), .ZN(new_n570));
  OAI21_X1  g384(.A(G107), .B1(new_n543), .B2(new_n538), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n551), .B1(new_n571), .B2(new_n550), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n568), .A2(new_n573), .A3(KEYINPUT97), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n525), .B1(new_n563), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n525), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n561), .B2(new_n562), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n228), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G478), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n578), .A2(new_n580), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n188), .A2(G952), .ZN(new_n584));
  INV_X1    g398(.A(G234), .ZN(new_n585));
  INV_X1    g399(.A(G237), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI211_X1 g402(.A(new_n228), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT21), .B(G898), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G475), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n214), .B(new_n199), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT18), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(KEYINPUT91), .ZN(new_n596));
  AND4_X1   g410(.A1(G143), .A2(new_n586), .A3(new_n188), .A4(G214), .ZN(new_n597));
  AOI21_X1  g411(.A(G143), .B1(new_n314), .B2(G214), .ZN(new_n598));
  OAI211_X1 g412(.A(G131), .B(new_n596), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n586), .A2(new_n188), .A3(G214), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n251), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(G131), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n314), .A2(G143), .A3(G214), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n594), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n597), .A2(new_n598), .A3(G131), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n247), .B1(new_n601), .B2(new_n603), .ZN(new_n607));
  NOR3_X1   g421(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT17), .ZN(new_n608));
  OAI211_X1 g422(.A(KEYINPUT17), .B(G131), .C1(new_n597), .C2(new_n598), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n200), .A2(new_n201), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n605), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(G113), .B(G122), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(new_n382), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n613), .B(new_n605), .C1(new_n608), .C2(new_n610), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n593), .B1(new_n617), .B2(new_n228), .ZN(new_n618));
  NOR2_X1   g432(.A1(G475), .A2(G902), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT92), .B1(new_n606), .B2(new_n607), .ZN(new_n620));
  OAI21_X1  g434(.A(G131), .B1(new_n597), .B2(new_n598), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT92), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n601), .A2(new_n247), .A3(new_n603), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT93), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n625), .A2(KEYINPUT19), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(KEYINPUT19), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n214), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n628), .B(new_n199), .C1(new_n214), .C2(new_n627), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n620), .A2(new_n201), .A3(new_n624), .A4(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n613), .B1(new_n630), .B2(new_n605), .ZN(new_n631));
  INV_X1    g445(.A(new_n616), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n619), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(KEYINPUT20), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT20), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n635), .B(new_n619), .C1(new_n631), .C2(new_n632), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n618), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n583), .A2(new_n592), .A3(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n470), .A2(new_n524), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n377), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G101), .ZN(G3));
  INV_X1    g455(.A(new_n469), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n464), .B2(new_n467), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n561), .A2(KEYINPUT98), .A3(new_n525), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n525), .A2(KEYINPUT98), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n568), .B2(new_n573), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT33), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n579), .A2(G902), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n563), .A2(new_n574), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n577), .B1(new_n649), .B2(new_n576), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n647), .B(new_n648), .C1(new_n650), .C2(KEYINPUT33), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n578), .A2(new_n579), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n637), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n643), .A2(new_n592), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n360), .A2(new_n361), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n228), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n362), .B1(new_n656), .B2(G472), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n523), .A2(new_n657), .A3(new_n235), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT34), .B(G104), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  OAI211_X1 g475(.A(new_n592), .B(new_n637), .C1(new_n581), .C2(new_n582), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n643), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n658), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT35), .B(G107), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  OR2_X1    g482(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n669), .A2(new_n217), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n217), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n232), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n230), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(KEYINPUT100), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n676), .B(new_n230), .C1(new_n672), .C2(new_n673), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n638), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n643), .A2(new_n523), .A3(new_n679), .A4(new_n657), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n374), .A2(new_n349), .A3(G472), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n364), .A2(new_n358), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n348), .A2(new_n349), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(G900), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n589), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n587), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n637), .B(new_n691), .C1(new_n581), .C2(new_n582), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n678), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n643), .A2(new_n523), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n683), .B1(new_n688), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n365), .A2(new_n376), .ZN(new_n696));
  INV_X1    g510(.A(new_n694), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(KEYINPUT101), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G128), .ZN(G30));
  XNOR2_X1  g514(.A(new_n691), .B(KEYINPUT39), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n523), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT40), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n468), .B(KEYINPUT38), .Z(new_n704));
  INV_X1    g518(.A(new_n344), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n351), .B1(new_n705), .B2(new_n318), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n237), .B1(new_n706), .B2(new_n228), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n685), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n674), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n583), .A2(new_n637), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n469), .ZN(new_n713));
  NOR4_X1   g527(.A1(new_n703), .A2(new_n704), .A3(new_n711), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n251), .ZN(G45));
  INV_X1    g529(.A(new_n653), .ZN(new_n716));
  INV_X1    g530(.A(new_n691), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n468), .A2(new_n469), .A3(new_n718), .ZN(new_n719));
  AOI211_X1 g533(.A(new_n473), .B(new_n678), .C1(new_n515), .C2(new_n522), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n719), .B(new_n720), .C1(new_n686), .C2(new_n687), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G146), .ZN(G48));
  INV_X1    g536(.A(new_n654), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n513), .A2(new_n228), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n472), .A3(new_n515), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n377), .A2(new_n723), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT102), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NOR2_X1   g546(.A1(new_n665), .A2(new_n726), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n377), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G116), .ZN(G18));
  OAI21_X1  g549(.A(KEYINPUT103), .B1(new_n470), .B2(new_n726), .ZN(new_n736));
  INV_X1    g550(.A(new_n515), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n514), .B1(new_n513), .B2(new_n228), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT103), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n643), .A3(new_n740), .A4(new_n472), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n679), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(new_n365), .B2(new_n376), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  NAND3_X1  g560(.A1(new_n468), .A2(new_n712), .A3(new_n469), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n725), .A2(new_n472), .A3(new_n515), .A4(new_n592), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n318), .B1(new_n345), .B2(new_n332), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n353), .B2(new_n354), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n357), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n753));
  AOI21_X1  g567(.A(G902), .B1(new_n360), .B2(new_n361), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n753), .B1(new_n754), .B2(new_n237), .ZN(new_n755));
  OAI211_X1 g569(.A(KEYINPUT104), .B(G472), .C1(new_n355), .C2(G902), .ZN(new_n756));
  AOI211_X1 g570(.A(new_n234), .B(new_n752), .C1(new_n755), .C2(new_n756), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n749), .A2(KEYINPUT105), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT105), .B1(new_n749), .B2(new_n757), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n535), .ZN(G24));
  NAND2_X1  g575(.A1(new_n755), .A2(new_n756), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n651), .A2(new_n652), .ZN(new_n764));
  INV_X1    g578(.A(new_n637), .ZN(new_n765));
  AND4_X1   g579(.A1(new_n763), .A2(new_n764), .A3(new_n765), .A4(new_n691), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n763), .B1(new_n653), .B2(new_n691), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n752), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n762), .A2(new_n674), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n770), .B1(new_n736), .B2(new_n741), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n194), .ZN(G27));
  OAI21_X1  g586(.A(KEYINPUT108), .B1(new_n468), .B2(new_n642), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n464), .A2(new_n467), .A3(new_n774), .A4(new_n469), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT107), .B1(new_n517), .B2(new_n495), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n776), .B1(new_n520), .B2(KEYINPUT107), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n516), .B1(new_n777), .B2(G469), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n473), .B1(new_n778), .B2(new_n515), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n773), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT42), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n781), .A2(new_n377), .A3(new_n782), .A4(new_n768), .ZN(new_n783));
  INV_X1    g597(.A(new_n234), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n784), .B(new_n768), .C1(new_n686), .C2(new_n687), .ZN(new_n785));
  OAI21_X1  g599(.A(KEYINPUT42), .B1(new_n785), .B2(new_n780), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n247), .ZN(G33));
  NOR2_X1   g602(.A1(new_n583), .A2(new_n765), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n781), .A2(new_n377), .A3(new_n789), .A4(new_n691), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  AOI21_X1  g605(.A(new_n765), .B1(new_n652), .B2(new_n651), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT43), .Z(new_n793));
  NOR3_X1   g607(.A1(new_n793), .A2(new_n657), .A3(new_n710), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT44), .ZN(new_n795));
  OAI21_X1  g609(.A(G469), .B1(new_n521), .B2(KEYINPUT45), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(KEYINPUT45), .B2(new_n777), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n516), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(KEYINPUT46), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n515), .B1(new_n798), .B2(KEYINPUT46), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n472), .B(new_n701), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n773), .A2(new_n775), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n795), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT109), .B(G137), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(G39));
  OAI21_X1  g620(.A(new_n472), .B1(new_n799), .B2(new_n800), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n807), .A2(KEYINPUT110), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(KEYINPUT110), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT111), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(KEYINPUT111), .A3(new_n810), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n810), .A2(KEYINPUT111), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n808), .A2(new_n814), .A3(new_n809), .A4(new_n811), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n236), .A2(new_n802), .A3(new_n688), .A4(new_n718), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  INV_X1    g633(.A(new_n739), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT112), .Z(new_n822));
  NAND4_X1  g636(.A1(new_n792), .A2(new_n784), .A3(new_n472), .A4(new_n469), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n823), .B(new_n709), .C1(KEYINPUT49), .C2(new_n820), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n704), .A3(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n803), .A2(new_n587), .A3(new_n726), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n709), .A2(new_n236), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n828), .A2(new_n765), .A3(new_n764), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n762), .A2(new_n784), .A3(new_n769), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n832), .A2(new_n793), .A3(new_n587), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n833), .A2(new_n642), .A3(new_n704), .A4(new_n727), .ZN(new_n834));
  NAND2_X1  g648(.A1(KEYINPUT119), .A2(KEYINPUT50), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n834), .B(new_n835), .Z(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(KEYINPUT119), .B2(KEYINPUT50), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n762), .A2(new_n674), .A3(new_n769), .ZN(new_n838));
  INV_X1    g652(.A(new_n793), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n826), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n831), .B(new_n837), .C1(new_n838), .C2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT51), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n813), .A2(new_n815), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n739), .A2(new_n473), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT121), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n844), .A2(new_n848), .A3(new_n845), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n833), .A2(new_n802), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n847), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n843), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g666(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n853));
  AND2_X1   g667(.A1(new_n846), .A2(new_n850), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(new_n841), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n696), .A2(new_n784), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n840), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT48), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n833), .A2(new_n742), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n584), .B(new_n859), .C1(new_n828), .C2(new_n716), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n852), .A2(new_n855), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n468), .A2(new_n469), .A3(new_n592), .A4(new_n789), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n680), .B1(new_n658), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n745), .A2(new_n640), .A3(new_n734), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n654), .A2(KEYINPUT113), .ZN(new_n868));
  INV_X1    g682(.A(new_n658), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT113), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n643), .A2(new_n870), .A3(new_n592), .A4(new_n653), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n758), .B2(new_n759), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n783), .A2(new_n790), .A3(new_n786), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n780), .A2(new_n770), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n581), .A2(new_n765), .A3(new_n582), .A4(new_n717), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n773), .A2(new_n775), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT114), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n696), .A2(new_n720), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n874), .A2(new_n730), .A3(new_n875), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n771), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n674), .B1(new_n685), .B2(new_n708), .ZN(new_n884));
  AOI211_X1 g698(.A(new_n473), .B(new_n717), .C1(new_n778), .C2(new_n515), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n884), .A2(new_n643), .A3(new_n712), .A4(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n721), .A2(new_n886), .ZN(new_n887));
  AND4_X1   g701(.A1(KEYINPUT52), .A2(new_n699), .A3(new_n883), .A4(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n771), .B1(new_n695), .B2(new_n698), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT52), .B1(new_n889), .B2(new_n887), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT116), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n889), .A2(new_n887), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT52), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT116), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n889), .A2(KEYINPUT52), .A3(new_n887), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n863), .B(new_n882), .C1(new_n891), .C2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT115), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n888), .B2(new_n890), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n894), .A2(KEYINPUT115), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n882), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT53), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT54), .B1(new_n898), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n902), .A2(KEYINPUT53), .A3(new_n903), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT54), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n882), .B1(new_n897), .B2(new_n891), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n906), .B(new_n907), .C1(KEYINPUT53), .C2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n905), .A2(KEYINPUT117), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n911), .B(KEYINPUT54), .C1(new_n898), .C2(new_n904), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n862), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n825), .B1(new_n913), .B2(new_n914), .ZN(G75));
  OAI21_X1  g729(.A(new_n906), .B1(KEYINPUT53), .B2(new_n908), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n916), .A2(G902), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(G210), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n456), .A2(new_n458), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n452), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT55), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n918), .A2(new_n919), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n922), .B1(new_n918), .B2(new_n919), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n188), .A2(G952), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(G51));
  XOR2_X1   g740(.A(new_n513), .B(KEYINPUT122), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n916), .B(new_n907), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n516), .B(KEYINPUT57), .Z(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n917), .A2(new_n797), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n925), .B1(new_n930), .B2(new_n931), .ZN(G54));
  NAND3_X1  g746(.A1(new_n917), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n631), .A2(new_n632), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n935), .A2(new_n936), .A3(new_n925), .ZN(G60));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT59), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n910), .A2(new_n912), .A3(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n650), .A2(KEYINPUT33), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n942), .A2(new_n647), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n940), .A2(new_n941), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n941), .B1(new_n940), .B2(new_n944), .ZN(new_n946));
  INV_X1    g760(.A(new_n925), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n939), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n928), .B2(new_n948), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(G63));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT60), .Z(new_n952));
  AND2_X1   g766(.A1(new_n916), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n947), .B1(new_n953), .B2(new_n231), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n916), .A2(new_n952), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(new_n672), .ZN(new_n957));
  INV_X1    g771(.A(new_n672), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n953), .A2(KEYINPUT124), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n954), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n953), .B2(new_n231), .ZN(new_n962));
  INV_X1    g776(.A(new_n231), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n956), .A2(KEYINPUT125), .A3(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n962), .A2(KEYINPUT61), .A3(new_n947), .A4(new_n964), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n959), .A2(new_n957), .ZN(new_n966));
  OAI22_X1  g780(.A1(new_n960), .A2(KEYINPUT61), .B1(new_n965), .B2(new_n966), .ZN(G66));
  OAI21_X1  g781(.A(G953), .B1(new_n590), .B2(new_n428), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n874), .A2(new_n730), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n968), .B1(new_n970), .B2(G953), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n920), .B1(G898), .B2(new_n188), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n971), .B(new_n972), .ZN(G69));
  NAND2_X1  g787(.A1(new_n290), .A2(new_n308), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n628), .B1(new_n214), .B2(new_n627), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n804), .B1(new_n816), .B2(new_n817), .ZN(new_n977));
  INV_X1    g791(.A(new_n377), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n789), .A2(new_n653), .ZN(new_n979));
  OR3_X1    g793(.A1(new_n803), .A2(new_n702), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n977), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n889), .A2(new_n721), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(new_n714), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n188), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n981), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n976), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n493), .A2(G900), .A3(G953), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n875), .B(KEYINPUT126), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n801), .A2(new_n747), .A3(new_n856), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n982), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n977), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n989), .B1(new_n994), .B2(G953), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n988), .B1(new_n976), .B2(new_n995), .ZN(G72));
  OR2_X1    g810(.A1(new_n898), .A2(new_n904), .ZN(new_n997));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  NAND2_X1  g813(.A1(new_n322), .A2(new_n351), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n984), .A2(new_n970), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n999), .B1(new_n981), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n313), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n999), .B1(new_n993), .B2(new_n969), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n319), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  AOI211_X1 g821(.A(new_n925), .B(new_n1001), .C1(new_n1007), .C2(new_n366), .ZN(G57));
endmodule


