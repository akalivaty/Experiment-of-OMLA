

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(KEYINPUT71), .B(n618), .ZN(n948) );
  XNOR2_X1 U552 ( .A(n521), .B(n520), .ZN(n524) );
  INV_X1 U553 ( .A(KEYINPUT23), .ZN(n520) );
  NOR2_X1 U554 ( .A1(n588), .A2(n589), .ZN(G164) );
  NOR2_X1 U555 ( .A1(n727), .A2(n725), .ZN(n517) );
  INV_X1 U556 ( .A(KEYINPUT30), .ZN(n649) );
  XNOR2_X1 U557 ( .A(n650), .B(n649), .ZN(n651) );
  INV_X1 U558 ( .A(n595), .ZN(n634) );
  NOR2_X1 U559 ( .A1(G1966), .A2(n727), .ZN(n646) );
  INV_X1 U560 ( .A(KEYINPUT32), .ZN(n671) );
  XNOR2_X1 U561 ( .A(n594), .B(KEYINPUT64), .ZN(n595) );
  NOR2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  XNOR2_X1 U563 ( .A(n519), .B(KEYINPUT65), .ZN(n568) );
  NOR2_X1 U564 ( .A1(G651), .A2(n535), .ZN(n785) );
  BUF_X1 U565 ( .A(n568), .Z(n881) );
  INV_X1 U566 ( .A(G2105), .ZN(n518) );
  NAND2_X1 U567 ( .A1(n518), .A2(G2104), .ZN(n519) );
  NAND2_X1 U568 ( .A1(n568), .A2(G101), .ZN(n521) );
  INV_X1 U569 ( .A(G2105), .ZN(n522) );
  NOR2_X1 U570 ( .A1(G2104), .A2(n522), .ZN(n571) );
  BUF_X1 U571 ( .A(n571), .Z(n877) );
  NAND2_X1 U572 ( .A1(n877), .A2(G125), .ZN(n523) );
  NAND2_X1 U573 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U574 ( .A(n525), .B(KEYINPUT66), .ZN(n531) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n878) );
  NAND2_X1 U576 ( .A1(n878), .A2(G113), .ZN(n529) );
  XOR2_X1 U577 ( .A(KEYINPUT17), .B(n526), .Z(n527) );
  BUF_X2 U578 ( .A(n527), .Z(n882) );
  NAND2_X1 U579 ( .A1(n882), .A2(G137), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X4 U581 ( .A1(n531), .A2(n530), .ZN(G160) );
  INV_X1 U582 ( .A(G651), .ZN(n536) );
  NOR2_X1 U583 ( .A1(G543), .A2(n536), .ZN(n532) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n532), .Z(n787) );
  NAND2_X1 U585 ( .A1(G64), .A2(n787), .ZN(n534) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n535) );
  NAND2_X1 U587 ( .A1(G52), .A2(n785), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n542) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n790) );
  NAND2_X1 U590 ( .A1(G90), .A2(n790), .ZN(n539) );
  OR2_X1 U591 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X2 U592 ( .A(KEYINPUT67), .B(n537), .ZN(n791) );
  NAND2_X1 U593 ( .A1(G77), .A2(n791), .ZN(n538) );
  NAND2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U595 ( .A(KEYINPUT9), .B(n540), .Z(n541) );
  NOR2_X1 U596 ( .A1(n542), .A2(n541), .ZN(G171) );
  NAND2_X1 U597 ( .A1(n790), .A2(G89), .ZN(n543) );
  XNOR2_X1 U598 ( .A(n543), .B(KEYINPUT4), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G76), .A2(n791), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U601 ( .A(n546), .B(KEYINPUT5), .ZN(n551) );
  NAND2_X1 U602 ( .A1(G63), .A2(n787), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G51), .A2(n785), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U605 ( .A(KEYINPUT6), .B(n549), .Z(n550) );
  NAND2_X1 U606 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U607 ( .A(n552), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U608 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U609 ( .A1(G50), .A2(n785), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G75), .A2(n791), .ZN(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U612 ( .A1(G62), .A2(n787), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G88), .A2(n790), .ZN(n555) );
  NAND2_X1 U614 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U615 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U616 ( .A(n559), .B(KEYINPUT78), .ZN(G166) );
  INV_X1 U617 ( .A(G166), .ZN(G303) );
  NAND2_X1 U618 ( .A1(n787), .A2(G61), .ZN(n566) );
  NAND2_X1 U619 ( .A1(G48), .A2(n785), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G86), .A2(n790), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n791), .A2(G73), .ZN(n562) );
  XOR2_X1 U623 ( .A(KEYINPUT2), .B(n562), .Z(n563) );
  NOR2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U626 ( .A(KEYINPUT77), .B(n567), .Z(G305) );
  NAND2_X1 U627 ( .A1(G102), .A2(n881), .ZN(n570) );
  NAND2_X1 U628 ( .A1(G138), .A2(n882), .ZN(n569) );
  NAND2_X1 U629 ( .A1(n570), .A2(n569), .ZN(n588) );
  NAND2_X1 U630 ( .A1(n571), .A2(G126), .ZN(n572) );
  XNOR2_X1 U631 ( .A(n572), .B(KEYINPUT80), .ZN(n574) );
  NAND2_X1 U632 ( .A1(G114), .A2(n878), .ZN(n573) );
  NAND2_X1 U633 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U634 ( .A(KEYINPUT81), .B(n575), .Z(n589) );
  NAND2_X1 U635 ( .A1(G60), .A2(n787), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G47), .A2(n785), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U638 ( .A(KEYINPUT68), .B(n578), .Z(n582) );
  NAND2_X1 U639 ( .A1(G85), .A2(n790), .ZN(n580) );
  NAND2_X1 U640 ( .A1(G72), .A2(n791), .ZN(n579) );
  AND2_X1 U641 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n582), .A2(n581), .ZN(G290) );
  NAND2_X1 U643 ( .A1(G49), .A2(n785), .ZN(n584) );
  NAND2_X1 U644 ( .A1(G74), .A2(G651), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U646 ( .A1(n787), .A2(n585), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n535), .A2(G87), .ZN(n586) );
  NAND2_X1 U648 ( .A1(n587), .A2(n586), .ZN(G288) );
  NOR2_X1 U649 ( .A1(n589), .A2(n588), .ZN(n592) );
  INV_X1 U650 ( .A(G40), .ZN(n590) );
  OR2_X1 U651 ( .A1(n590), .A2(G1384), .ZN(n591) );
  NOR2_X1 U652 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U653 ( .A1(G160), .A2(n593), .ZN(n594) );
  NAND2_X1 U654 ( .A1(n595), .A2(G8), .ZN(n727) );
  INV_X1 U655 ( .A(n634), .ZN(n663) );
  AND2_X1 U656 ( .A1(n663), .A2(G1961), .ZN(n597) );
  XNOR2_X1 U657 ( .A(G2078), .B(KEYINPUT25), .ZN(n1003) );
  NOR2_X1 U658 ( .A1(n663), .A2(n1003), .ZN(n596) );
  NOR2_X1 U659 ( .A1(n597), .A2(n596), .ZN(n652) );
  NAND2_X1 U660 ( .A1(n652), .A2(G171), .ZN(n645) );
  NAND2_X1 U661 ( .A1(G56), .A2(n787), .ZN(n598) );
  XOR2_X1 U662 ( .A(KEYINPUT14), .B(n598), .Z(n604) );
  NAND2_X1 U663 ( .A1(n790), .A2(G81), .ZN(n599) );
  XNOR2_X1 U664 ( .A(n599), .B(KEYINPUT12), .ZN(n601) );
  NAND2_X1 U665 ( .A1(G68), .A2(n791), .ZN(n600) );
  NAND2_X1 U666 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U667 ( .A(KEYINPUT13), .B(n602), .Z(n603) );
  NOR2_X1 U668 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U669 ( .A1(n785), .A2(G43), .ZN(n605) );
  NAND2_X1 U670 ( .A1(n606), .A2(n605), .ZN(n958) );
  NAND2_X1 U671 ( .A1(G1996), .A2(n634), .ZN(n607) );
  XOR2_X1 U672 ( .A(KEYINPUT26), .B(n607), .Z(n608) );
  NOR2_X1 U673 ( .A1(n958), .A2(n608), .ZN(n610) );
  NAND2_X1 U674 ( .A1(n663), .A2(G1341), .ZN(n609) );
  NAND2_X1 U675 ( .A1(n610), .A2(n609), .ZN(n624) );
  NAND2_X1 U676 ( .A1(G66), .A2(n787), .ZN(n612) );
  NAND2_X1 U677 ( .A1(G92), .A2(n790), .ZN(n611) );
  NAND2_X1 U678 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U679 ( .A1(G54), .A2(n785), .ZN(n614) );
  NAND2_X1 U680 ( .A1(G79), .A2(n791), .ZN(n613) );
  NAND2_X1 U681 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U682 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U683 ( .A(KEYINPUT15), .B(n617), .Z(n618) );
  NOR2_X2 U684 ( .A1(n624), .A2(n948), .ZN(n619) );
  XOR2_X1 U685 ( .A(n619), .B(KEYINPUT86), .Z(n623) );
  NOR2_X1 U686 ( .A1(G2067), .A2(n663), .ZN(n621) );
  NOR2_X1 U687 ( .A1(G1348), .A2(n634), .ZN(n620) );
  NOR2_X1 U688 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U689 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U690 ( .A1(n624), .A2(n948), .ZN(n625) );
  NAND2_X1 U691 ( .A1(n626), .A2(n625), .ZN(n638) );
  NAND2_X1 U692 ( .A1(G65), .A2(n787), .ZN(n628) );
  NAND2_X1 U693 ( .A1(G53), .A2(n785), .ZN(n627) );
  NAND2_X1 U694 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U695 ( .A1(G91), .A2(n790), .ZN(n630) );
  NAND2_X1 U696 ( .A1(G78), .A2(n791), .ZN(n629) );
  NAND2_X1 U697 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U698 ( .A1(n632), .A2(n631), .ZN(n951) );
  NAND2_X1 U699 ( .A1(G2072), .A2(n634), .ZN(n633) );
  XNOR2_X1 U700 ( .A(n633), .B(KEYINPUT27), .ZN(n636) );
  INV_X1 U701 ( .A(G1956), .ZN(n984) );
  NOR2_X1 U702 ( .A1(n634), .A2(n984), .ZN(n635) );
  NOR2_X1 U703 ( .A1(n636), .A2(n635), .ZN(n639) );
  NAND2_X1 U704 ( .A1(n951), .A2(n639), .ZN(n637) );
  NAND2_X1 U705 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U706 ( .A1(n951), .A2(n639), .ZN(n640) );
  XOR2_X1 U707 ( .A(n640), .B(KEYINPUT28), .Z(n641) );
  NAND2_X1 U708 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U709 ( .A(KEYINPUT29), .B(n643), .Z(n644) );
  NAND2_X1 U710 ( .A1(n645), .A2(n644), .ZN(n659) );
  XOR2_X1 U711 ( .A(KEYINPUT85), .B(n646), .Z(n676) );
  NOR2_X1 U712 ( .A1(n663), .A2(G2084), .ZN(n673) );
  NOR2_X1 U713 ( .A1(n676), .A2(n673), .ZN(n647) );
  NAND2_X1 U714 ( .A1(G8), .A2(n647), .ZN(n648) );
  XNOR2_X1 U715 ( .A(n648), .B(KEYINPUT87), .ZN(n650) );
  NOR2_X1 U716 ( .A1(G168), .A2(n651), .ZN(n654) );
  NOR2_X1 U717 ( .A1(G171), .A2(n652), .ZN(n653) );
  NOR2_X1 U718 ( .A1(n654), .A2(n653), .ZN(n657) );
  XNOR2_X1 U719 ( .A(KEYINPUT88), .B(KEYINPUT89), .ZN(n655) );
  XNOR2_X1 U720 ( .A(n655), .B(KEYINPUT31), .ZN(n656) );
  XNOR2_X1 U721 ( .A(n657), .B(n656), .ZN(n658) );
  NAND2_X1 U722 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U723 ( .A(n660), .B(KEYINPUT90), .ZN(n674) );
  AND2_X1 U724 ( .A1(G286), .A2(G8), .ZN(n661) );
  NAND2_X1 U725 ( .A1(n674), .A2(n661), .ZN(n670) );
  INV_X1 U726 ( .A(G8), .ZN(n668) );
  NOR2_X1 U727 ( .A1(G1971), .A2(n727), .ZN(n662) );
  XNOR2_X1 U728 ( .A(KEYINPUT91), .B(n662), .ZN(n666) );
  NOR2_X1 U729 ( .A1(n663), .A2(G2090), .ZN(n664) );
  NOR2_X1 U730 ( .A1(G166), .A2(n664), .ZN(n665) );
  NAND2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n667) );
  OR2_X1 U732 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U733 ( .A1(n670), .A2(n669), .ZN(n672) );
  XNOR2_X1 U734 ( .A(n672), .B(n671), .ZN(n680) );
  NAND2_X1 U735 ( .A1(G8), .A2(n673), .ZN(n678) );
  INV_X1 U736 ( .A(n674), .ZN(n675) );
  NOR2_X1 U737 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U739 ( .A1(n680), .A2(n679), .ZN(n722) );
  NOR2_X1 U740 ( .A1(G2090), .A2(G303), .ZN(n681) );
  NAND2_X1 U741 ( .A1(G8), .A2(n681), .ZN(n682) );
  NAND2_X1 U742 ( .A1(n722), .A2(n682), .ZN(n683) );
  NAND2_X1 U743 ( .A1(n727), .A2(n683), .ZN(n684) );
  XNOR2_X1 U744 ( .A(n684), .B(KEYINPUT94), .ZN(n688) );
  NOR2_X1 U745 ( .A1(G1981), .A2(G305), .ZN(n685) );
  XOR2_X1 U746 ( .A(n685), .B(KEYINPUT24), .Z(n686) );
  OR2_X1 U747 ( .A1(n727), .A2(n686), .ZN(n687) );
  NAND2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n720) );
  NOR2_X1 U749 ( .A1(G164), .A2(G1384), .ZN(n690) );
  NAND2_X1 U750 ( .A1(G160), .A2(G40), .ZN(n689) );
  NOR2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n753) );
  NAND2_X1 U752 ( .A1(G104), .A2(n881), .ZN(n692) );
  NAND2_X1 U753 ( .A1(G140), .A2(n882), .ZN(n691) );
  NAND2_X1 U754 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U755 ( .A(KEYINPUT34), .B(n693), .ZN(n699) );
  NAND2_X1 U756 ( .A1(n877), .A2(G128), .ZN(n694) );
  XNOR2_X1 U757 ( .A(n694), .B(KEYINPUT82), .ZN(n696) );
  NAND2_X1 U758 ( .A1(G116), .A2(n878), .ZN(n695) );
  NAND2_X1 U759 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U760 ( .A(KEYINPUT35), .B(n697), .Z(n698) );
  NOR2_X1 U761 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U762 ( .A(KEYINPUT36), .B(n700), .ZN(n896) );
  XNOR2_X1 U763 ( .A(KEYINPUT37), .B(G2067), .ZN(n750) );
  NOR2_X1 U764 ( .A1(n896), .A2(n750), .ZN(n930) );
  NAND2_X1 U765 ( .A1(n753), .A2(n930), .ZN(n748) );
  NAND2_X1 U766 ( .A1(G119), .A2(n877), .ZN(n702) );
  NAND2_X1 U767 ( .A1(G131), .A2(n882), .ZN(n701) );
  NAND2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U769 ( .A1(G95), .A2(n881), .ZN(n704) );
  NAND2_X1 U770 ( .A1(G107), .A2(n878), .ZN(n703) );
  NAND2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n891) );
  INV_X1 U773 ( .A(G1991), .ZN(n741) );
  NOR2_X1 U774 ( .A1(n891), .A2(n741), .ZN(n717) );
  NAND2_X1 U775 ( .A1(G129), .A2(n877), .ZN(n708) );
  NAND2_X1 U776 ( .A1(G117), .A2(n878), .ZN(n707) );
  NAND2_X1 U777 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U778 ( .A1(n881), .A2(G105), .ZN(n709) );
  XOR2_X1 U779 ( .A(KEYINPUT38), .B(n709), .Z(n710) );
  NOR2_X1 U780 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U781 ( .A(KEYINPUT83), .B(n712), .ZN(n715) );
  NAND2_X1 U782 ( .A1(n882), .A2(G141), .ZN(n713) );
  XOR2_X1 U783 ( .A(KEYINPUT84), .B(n713), .Z(n714) );
  OR2_X1 U784 ( .A1(n715), .A2(n714), .ZN(n895) );
  AND2_X1 U785 ( .A1(G1996), .A2(n895), .ZN(n716) );
  NOR2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n928) );
  XOR2_X1 U787 ( .A(G1986), .B(G290), .Z(n950) );
  NAND2_X1 U788 ( .A1(n928), .A2(n950), .ZN(n718) );
  NAND2_X1 U789 ( .A1(n753), .A2(n718), .ZN(n719) );
  AND2_X1 U790 ( .A1(n748), .A2(n719), .ZN(n729) );
  NAND2_X1 U791 ( .A1(n720), .A2(n729), .ZN(n739) );
  NOR2_X1 U792 ( .A1(G1976), .A2(G288), .ZN(n726) );
  NOR2_X1 U793 ( .A1(G303), .A2(G1971), .ZN(n721) );
  NOR2_X1 U794 ( .A1(n726), .A2(n721), .ZN(n955) );
  NAND2_X1 U795 ( .A1(n722), .A2(n955), .ZN(n723) );
  XNOR2_X1 U796 ( .A(n723), .B(KEYINPUT92), .ZN(n732) );
  NAND2_X1 U797 ( .A1(G288), .A2(G1976), .ZN(n724) );
  XOR2_X1 U798 ( .A(KEYINPUT93), .B(n724), .Z(n954) );
  INV_X1 U799 ( .A(n954), .ZN(n725) );
  NAND2_X1 U800 ( .A1(n726), .A2(KEYINPUT33), .ZN(n728) );
  OR2_X1 U801 ( .A1(n728), .A2(n727), .ZN(n733) );
  AND2_X1 U802 ( .A1(n517), .A2(n733), .ZN(n730) );
  XOR2_X1 U803 ( .A(G1981), .B(G305), .Z(n966) );
  AND2_X1 U804 ( .A1(n966), .A2(n729), .ZN(n735) );
  AND2_X1 U805 ( .A1(n730), .A2(n735), .ZN(n731) );
  NAND2_X1 U806 ( .A1(n732), .A2(n731), .ZN(n737) );
  AND2_X1 U807 ( .A1(n733), .A2(KEYINPUT33), .ZN(n734) );
  NAND2_X1 U808 ( .A1(n735), .A2(n734), .ZN(n736) );
  AND2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U810 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U811 ( .A(n740), .B(KEYINPUT95), .ZN(n755) );
  NOR2_X1 U812 ( .A1(G1996), .A2(n895), .ZN(n938) );
  INV_X1 U813 ( .A(n928), .ZN(n745) );
  AND2_X1 U814 ( .A1(n741), .A2(n891), .ZN(n742) );
  XNOR2_X1 U815 ( .A(KEYINPUT96), .B(n742), .ZN(n922) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n743) );
  NOR2_X1 U817 ( .A1(n922), .A2(n743), .ZN(n744) );
  NOR2_X1 U818 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U819 ( .A1(n938), .A2(n746), .ZN(n747) );
  XNOR2_X1 U820 ( .A(KEYINPUT39), .B(n747), .ZN(n749) );
  NAND2_X1 U821 ( .A1(n749), .A2(n748), .ZN(n751) );
  NAND2_X1 U822 ( .A1(n896), .A2(n750), .ZN(n927) );
  NAND2_X1 U823 ( .A1(n751), .A2(n927), .ZN(n752) );
  NAND2_X1 U824 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U825 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U826 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U827 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U828 ( .A(G57), .ZN(G237) );
  INV_X1 U829 ( .A(G132), .ZN(G219) );
  INV_X1 U830 ( .A(G82), .ZN(G220) );
  NAND2_X1 U831 ( .A1(G7), .A2(G661), .ZN(n757) );
  XNOR2_X1 U832 ( .A(n757), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U833 ( .A(G223), .ZN(n831) );
  NAND2_X1 U834 ( .A1(n831), .A2(G567), .ZN(n758) );
  XNOR2_X1 U835 ( .A(n758), .B(KEYINPUT69), .ZN(n759) );
  XNOR2_X1 U836 ( .A(KEYINPUT11), .B(n759), .ZN(G234) );
  INV_X1 U837 ( .A(G860), .ZN(n784) );
  OR2_X1 U838 ( .A1(n958), .A2(n784), .ZN(G153) );
  XOR2_X1 U839 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  INV_X1 U840 ( .A(G868), .ZN(n806) );
  NAND2_X1 U841 ( .A1(n948), .A2(n806), .ZN(n760) );
  XNOR2_X1 U842 ( .A(n760), .B(KEYINPUT72), .ZN(n762) );
  NAND2_X1 U843 ( .A1(G301), .A2(G868), .ZN(n761) );
  NAND2_X1 U844 ( .A1(n762), .A2(n761), .ZN(G284) );
  INV_X1 U845 ( .A(n951), .ZN(G299) );
  NOR2_X1 U846 ( .A1(G286), .A2(n806), .ZN(n763) );
  XOR2_X1 U847 ( .A(KEYINPUT73), .B(n763), .Z(n765) );
  NOR2_X1 U848 ( .A1(G868), .A2(G299), .ZN(n764) );
  NOR2_X1 U849 ( .A1(n765), .A2(n764), .ZN(G297) );
  NAND2_X1 U850 ( .A1(n784), .A2(G559), .ZN(n766) );
  INV_X1 U851 ( .A(n948), .ZN(n782) );
  NAND2_X1 U852 ( .A1(n766), .A2(n782), .ZN(n767) );
  XNOR2_X1 U853 ( .A(n767), .B(KEYINPUT16), .ZN(n768) );
  XNOR2_X1 U854 ( .A(KEYINPUT74), .B(n768), .ZN(G148) );
  NOR2_X1 U855 ( .A1(G868), .A2(n958), .ZN(n771) );
  NAND2_X1 U856 ( .A1(n782), .A2(G868), .ZN(n769) );
  NOR2_X1 U857 ( .A1(G559), .A2(n769), .ZN(n770) );
  NOR2_X1 U858 ( .A1(n771), .A2(n770), .ZN(G282) );
  NAND2_X1 U859 ( .A1(G123), .A2(n877), .ZN(n772) );
  XNOR2_X1 U860 ( .A(n772), .B(KEYINPUT18), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G135), .A2(n882), .ZN(n773) );
  XOR2_X1 U862 ( .A(KEYINPUT75), .B(n773), .Z(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n779) );
  NAND2_X1 U864 ( .A1(G99), .A2(n881), .ZN(n777) );
  NAND2_X1 U865 ( .A1(G111), .A2(n878), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n921) );
  XNOR2_X1 U868 ( .A(n921), .B(G2096), .ZN(n781) );
  INV_X1 U869 ( .A(G2100), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(G156) );
  NAND2_X1 U871 ( .A1(G559), .A2(n782), .ZN(n783) );
  XOR2_X1 U872 ( .A(n958), .B(n783), .Z(n802) );
  NAND2_X1 U873 ( .A1(n784), .A2(n802), .ZN(n796) );
  NAND2_X1 U874 ( .A1(G55), .A2(n785), .ZN(n786) );
  XNOR2_X1 U875 ( .A(n786), .B(KEYINPUT76), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n787), .A2(G67), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n795) );
  NAND2_X1 U878 ( .A1(G93), .A2(n790), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G80), .A2(n791), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U881 ( .A1(n795), .A2(n794), .ZN(n805) );
  XOR2_X1 U882 ( .A(n796), .B(n805), .Z(G145) );
  XNOR2_X1 U883 ( .A(n951), .B(n805), .ZN(n799) );
  XNOR2_X1 U884 ( .A(KEYINPUT19), .B(G290), .ZN(n797) );
  XNOR2_X1 U885 ( .A(n797), .B(G288), .ZN(n798) );
  XNOR2_X1 U886 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U887 ( .A(G303), .B(n800), .ZN(n801) );
  XNOR2_X1 U888 ( .A(n801), .B(G305), .ZN(n907) );
  XOR2_X1 U889 ( .A(n802), .B(n907), .Z(n803) );
  XNOR2_X1 U890 ( .A(KEYINPUT79), .B(n803), .ZN(n804) );
  NOR2_X1 U891 ( .A1(n806), .A2(n804), .ZN(n808) );
  AND2_X1 U892 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U893 ( .A1(n808), .A2(n807), .ZN(G295) );
  NAND2_X1 U894 ( .A1(G2084), .A2(G2078), .ZN(n809) );
  XOR2_X1 U895 ( .A(KEYINPUT20), .B(n809), .Z(n810) );
  NAND2_X1 U896 ( .A1(G2090), .A2(n810), .ZN(n811) );
  XNOR2_X1 U897 ( .A(KEYINPUT21), .B(n811), .ZN(n812) );
  NAND2_X1 U898 ( .A1(n812), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U899 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U900 ( .A1(G220), .A2(G219), .ZN(n813) );
  XOR2_X1 U901 ( .A(KEYINPUT22), .B(n813), .Z(n814) );
  NOR2_X1 U902 ( .A1(G218), .A2(n814), .ZN(n815) );
  NAND2_X1 U903 ( .A1(G96), .A2(n815), .ZN(n919) );
  NAND2_X1 U904 ( .A1(n919), .A2(G2106), .ZN(n819) );
  NAND2_X1 U905 ( .A1(G69), .A2(G120), .ZN(n816) );
  NOR2_X1 U906 ( .A1(G237), .A2(n816), .ZN(n817) );
  NAND2_X1 U907 ( .A1(G108), .A2(n817), .ZN(n920) );
  NAND2_X1 U908 ( .A1(n920), .A2(G567), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n835) );
  NAND2_X1 U910 ( .A1(G483), .A2(G661), .ZN(n820) );
  NOR2_X1 U911 ( .A1(n835), .A2(n820), .ZN(n834) );
  NAND2_X1 U912 ( .A1(n834), .A2(G36), .ZN(G176) );
  XOR2_X1 U913 ( .A(KEYINPUT97), .B(G2446), .Z(n822) );
  XNOR2_X1 U914 ( .A(G2435), .B(G2438), .ZN(n821) );
  XNOR2_X1 U915 ( .A(n822), .B(n821), .ZN(n829) );
  XOR2_X1 U916 ( .A(G2451), .B(G2430), .Z(n824) );
  XNOR2_X1 U917 ( .A(G2454), .B(G2427), .ZN(n823) );
  XNOR2_X1 U918 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U919 ( .A(n825), .B(G2443), .Z(n827) );
  XNOR2_X1 U920 ( .A(G1341), .B(G1348), .ZN(n826) );
  XNOR2_X1 U921 ( .A(n827), .B(n826), .ZN(n828) );
  XNOR2_X1 U922 ( .A(n829), .B(n828), .ZN(n830) );
  NAND2_X1 U923 ( .A1(n830), .A2(G14), .ZN(n911) );
  XOR2_X1 U924 ( .A(KEYINPUT98), .B(n911), .Z(G401) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U927 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U929 ( .A1(n834), .A2(n833), .ZN(G188) );
  INV_X1 U930 ( .A(n835), .ZN(G319) );
  XOR2_X1 U931 ( .A(KEYINPUT42), .B(G2090), .Z(n837) );
  XNOR2_X1 U932 ( .A(G2084), .B(G2078), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U934 ( .A(n838), .B(G2100), .Z(n840) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2072), .ZN(n839) );
  XNOR2_X1 U936 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U937 ( .A(G2096), .B(KEYINPUT43), .Z(n842) );
  XNOR2_X1 U938 ( .A(KEYINPUT99), .B(G2678), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U940 ( .A(n844), .B(n843), .Z(G227) );
  XOR2_X1 U941 ( .A(G1966), .B(G1971), .Z(n846) );
  XNOR2_X1 U942 ( .A(G1981), .B(G1976), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n856) );
  XOR2_X1 U944 ( .A(KEYINPUT41), .B(KEYINPUT101), .Z(n848) );
  XNOR2_X1 U945 ( .A(G1996), .B(KEYINPUT100), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U947 ( .A(G1956), .B(G1961), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1991), .B(G1986), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U951 ( .A(G2474), .B(KEYINPUT102), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U954 ( .A1(G100), .A2(n881), .ZN(n858) );
  NAND2_X1 U955 ( .A1(G112), .A2(n878), .ZN(n857) );
  NAND2_X1 U956 ( .A1(n858), .A2(n857), .ZN(n864) );
  NAND2_X1 U957 ( .A1(n877), .A2(G124), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U959 ( .A1(G136), .A2(n882), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U961 ( .A(KEYINPUT103), .B(n862), .Z(n863) );
  NOR2_X1 U962 ( .A1(n864), .A2(n863), .ZN(G162) );
  XNOR2_X1 U963 ( .A(G164), .B(G162), .ZN(n900) );
  NAND2_X1 U964 ( .A1(G103), .A2(n881), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G139), .A2(n882), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G127), .A2(n877), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G115), .A2(n878), .ZN(n867) );
  NAND2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U970 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n933) );
  XOR2_X1 U972 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT46), .B(KEYINPUT105), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U975 ( .A(n874), .B(KEYINPUT109), .Z(n876) );
  XNOR2_X1 U976 ( .A(KEYINPUT48), .B(KEYINPUT106), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(n890) );
  NAND2_X1 U978 ( .A1(G130), .A2(n877), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G118), .A2(n878), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n888) );
  NAND2_X1 U981 ( .A1(G106), .A2(n881), .ZN(n884) );
  NAND2_X1 U982 ( .A1(G142), .A2(n882), .ZN(n883) );
  NAND2_X1 U983 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n885), .Z(n886) );
  XNOR2_X1 U985 ( .A(KEYINPUT104), .B(n886), .ZN(n887) );
  NOR2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U987 ( .A(n890), .B(n889), .Z(n893) );
  XNOR2_X1 U988 ( .A(n891), .B(n921), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n933), .B(n894), .ZN(n898) );
  XOR2_X1 U991 ( .A(n896), .B(n895), .Z(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U993 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n901), .B(G160), .ZN(n902) );
  NOR2_X1 U995 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U996 ( .A(G171), .B(G286), .Z(n903) );
  XNOR2_X1 U997 ( .A(n958), .B(n903), .ZN(n909) );
  XNOR2_X1 U998 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n905) );
  XNOR2_X1 U999 ( .A(n948), .B(KEYINPUT110), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1001 ( .A(n907), .B(n906), .Z(n908) );
  XNOR2_X1 U1002 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n910), .ZN(G397) );
  NAND2_X1 U1004 ( .A1(G319), .A2(n911), .ZN(n915) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n912) );
  XOR2_X1 U1006 ( .A(KEYINPUT113), .B(n912), .Z(n913) );
  XNOR2_X1 U1007 ( .A(n913), .B(KEYINPUT49), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1009 ( .A(KEYINPUT114), .B(n916), .ZN(n918) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1011 ( .A1(n918), .A2(n917), .ZN(G225) );
  XNOR2_X1 U1012 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G120), .ZN(G236) );
  INV_X1 U1015 ( .A(G96), .ZN(G221) );
  INV_X1 U1016 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(G325) );
  INV_X1 U1018 ( .A(G325), .ZN(G261) );
  INV_X1 U1019 ( .A(G108), .ZN(G238) );
  NOR2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(n923), .B(KEYINPUT117), .ZN(n926) );
  XOR2_X1 U1022 ( .A(G2084), .B(G160), .Z(n924) );
  XNOR2_X1 U1023 ( .A(KEYINPUT116), .B(n924), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n932) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n943) );
  XOR2_X1 U1028 ( .A(G2072), .B(n933), .Z(n935) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(KEYINPUT50), .B(n936), .ZN(n941) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1034 ( .A(KEYINPUT51), .B(n939), .Z(n940) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n944), .ZN(n946) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n947), .A2(G29), .ZN(n1028) );
  XNOR2_X1 U1041 ( .A(G16), .B(KEYINPUT56), .ZN(n973) );
  XOR2_X1 U1042 ( .A(G1348), .B(n948), .Z(n949) );
  NAND2_X1 U1043 ( .A1(n950), .A2(n949), .ZN(n964) );
  XNOR2_X1 U1044 ( .A(G1956), .B(n951), .ZN(n953) );
  NAND2_X1 U1045 ( .A1(G1971), .A2(G303), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n957) );
  NAND2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n962) );
  XOR2_X1 U1049 ( .A(G171), .B(G1961), .Z(n960) );
  XNOR2_X1 U1050 ( .A(n958), .B(G1341), .ZN(n959) );
  NOR2_X1 U1051 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1052 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1053 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1054 ( .A(KEYINPUT123), .B(n965), .Z(n971) );
  XNOR2_X1 U1055 ( .A(G1966), .B(G168), .ZN(n967) );
  NAND2_X1 U1056 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1057 ( .A(n968), .B(KEYINPUT122), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(KEYINPUT57), .B(n969), .ZN(n970) );
  NAND2_X1 U1059 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1060 ( .A1(n973), .A2(n972), .ZN(n1001) );
  INV_X1 U1061 ( .A(G16), .ZN(n999) );
  XNOR2_X1 U1062 ( .A(G1986), .B(G24), .ZN(n978) );
  XNOR2_X1 U1063 ( .A(G1976), .B(G23), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(G1971), .B(G22), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(KEYINPUT125), .B(n976), .ZN(n977) );
  NOR2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1068 ( .A(KEYINPUT58), .B(n979), .ZN(n983) );
  XNOR2_X1 U1069 ( .A(G1966), .B(G21), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G1961), .B(G5), .ZN(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n995) );
  XNOR2_X1 U1073 ( .A(G20), .B(n984), .ZN(n988) );
  XNOR2_X1 U1074 ( .A(G1981), .B(G6), .ZN(n986) );
  XNOR2_X1 U1075 ( .A(G1341), .B(G19), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n991) );
  XOR2_X1 U1078 ( .A(KEYINPUT59), .B(G1348), .Z(n989) );
  XNOR2_X1 U1079 ( .A(G4), .B(n989), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1081 ( .A(KEYINPUT60), .B(n992), .Z(n993) );
  XNOR2_X1 U1082 ( .A(KEYINPUT124), .B(n993), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1084 ( .A(n996), .B(KEYINPUT126), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(n997), .B(KEYINPUT61), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1026) );
  XOR2_X1 U1088 ( .A(G2084), .B(G34), .Z(n1002) );
  XNOR2_X1 U1089 ( .A(KEYINPUT54), .B(n1002), .ZN(n1018) );
  XNOR2_X1 U1090 ( .A(G2090), .B(G35), .ZN(n1016) );
  XNOR2_X1 U1091 ( .A(G27), .B(n1003), .ZN(n1007) );
  XNOR2_X1 U1092 ( .A(G2067), .B(G26), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G33), .B(G2072), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G32), .B(G1996), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1098 ( .A(KEYINPUT118), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(G28), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G25), .B(G1991), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT53), .B(n1014), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(n1019), .B(KEYINPUT119), .ZN(n1020) );
  XOR2_X1 U1106 ( .A(KEYINPUT55), .B(n1020), .Z(n1021) );
  NOR2_X1 U1107 ( .A1(G29), .A2(n1021), .ZN(n1022) );
  XOR2_X1 U1108 ( .A(KEYINPUT120), .B(n1022), .Z(n1023) );
  NAND2_X1 U1109 ( .A1(n1023), .A2(G11), .ZN(n1024) );
  XOR2_X1 U1110 ( .A(KEYINPUT121), .B(n1024), .Z(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(n1029), .B(KEYINPUT62), .ZN(n1030) );
  XNOR2_X1 U1114 ( .A(KEYINPUT127), .B(n1030), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

