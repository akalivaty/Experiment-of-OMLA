//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  XOR2_X1   g000(.A(KEYINPUT73), .B(G217), .Z(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G128), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT24), .B(G110), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(KEYINPUT23), .A3(G119), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n190), .A2(G128), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n197), .B(new_n191), .C1(new_n198), .C2(KEYINPUT23), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n196), .B1(new_n199), .B2(G110), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G125), .ZN(new_n203));
  XOR2_X1   g017(.A(G125), .B(G140), .Z(new_n204));
  OAI211_X1 g018(.A(G146), .B(new_n203), .C1(new_n204), .C2(new_n201), .ZN(new_n205));
  XNOR2_X1  g019(.A(G125), .B(G140), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n200), .A2(new_n205), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT75), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n209), .B(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n203), .B1(new_n204), .B2(new_n201), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n207), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(new_n205), .ZN(new_n214));
  INV_X1    g028(.A(G110), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n215), .B1(new_n199), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n216), .B2(new_n199), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n214), .B(new_n218), .C1(new_n194), .C2(new_n195), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n211), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G953), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G221), .A3(G234), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n222), .B(KEYINPUT76), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT22), .B(G137), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n223), .B(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n220), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n211), .A2(new_n219), .A3(new_n225), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT25), .B1(new_n229), .B2(new_n188), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n231));
  AOI211_X1 g045(.A(new_n231), .B(G902), .C1(new_n227), .C2(new_n228), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n189), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n189), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n188), .ZN(new_n236));
  XOR2_X1   g050(.A(new_n236), .B(KEYINPUT77), .Z(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(new_n227), .B2(new_n228), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(G472), .A2(G902), .ZN(new_n241));
  INV_X1    g055(.A(G143), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(G146), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n244), .B1(new_n207), .B2(G143), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n242), .A2(KEYINPUT65), .A3(G146), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n243), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n248), .A2(G128), .ZN(new_n249));
  OAI21_X1  g063(.A(G128), .B1(new_n248), .B2(new_n243), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n207), .A2(KEYINPUT64), .A3(G143), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT64), .B1(new_n207), .B2(G143), .ZN(new_n252));
  OAI22_X1  g066(.A1(new_n251), .A2(new_n252), .B1(G143), .B2(new_n207), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n247), .A2(new_n249), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G137), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G134), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G134), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(G137), .ZN(new_n261));
  AND2_X1   g075(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G131), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(G137), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n259), .A2(new_n263), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n257), .A2(new_n265), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G131), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n254), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT11), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n262), .B1(new_n261), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n265), .B1(new_n257), .B2(new_n255), .ZN(new_n275));
  OAI21_X1  g089(.A(G131), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n266), .ZN(new_n277));
  AND2_X1   g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  NOR2_X1   g092(.A1(KEYINPUT0), .A2(G128), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n253), .A2(new_n280), .B1(new_n247), .B2(new_n278), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT67), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n277), .A2(new_n284), .A3(new_n281), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n270), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT69), .B1(new_n286), .B2(KEYINPUT30), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n190), .A2(G116), .ZN(new_n288));
  INV_X1    g102(.A(G116), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G119), .ZN(new_n290));
  INV_X1    g104(.A(G113), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n291), .A2(KEYINPUT2), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n291), .A2(KEYINPUT2), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n288), .B(new_n290), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n292), .A2(new_n293), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n288), .A2(new_n290), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n296), .B(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n249), .A2(new_n247), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n250), .A2(new_n253), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n266), .A3(new_n268), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n282), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT30), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n277), .A2(new_n284), .A3(new_n281), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n284), .B1(new_n277), .B2(new_n281), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n304), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n287), .A2(new_n300), .A3(new_n307), .A4(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n305), .A2(new_n300), .ZN(new_n315));
  NOR2_X1   g129(.A1(G237), .A2(G953), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G210), .ZN(new_n317));
  XOR2_X1   g131(.A(new_n317), .B(KEYINPUT27), .Z(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT26), .B(G101), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n318), .B(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n314), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT31), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(KEYINPUT71), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n322), .A2(new_n325), .A3(KEYINPUT31), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT31), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n314), .A2(new_n328), .A3(new_n321), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT28), .ZN(new_n330));
  INV_X1    g144(.A(new_n300), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(new_n306), .B2(new_n331), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n305), .A2(KEYINPUT28), .A3(new_n300), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n286), .A2(new_n331), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n320), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT72), .B1(new_n327), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n325), .B1(new_n322), .B2(KEYINPUT31), .ZN(new_n339));
  AOI211_X1 g153(.A(KEYINPUT71), .B(new_n328), .C1(new_n314), .C2(new_n321), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n337), .B(KEYINPUT72), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n241), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT32), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT72), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n341), .ZN(new_n349));
  INV_X1    g163(.A(new_n241), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n350), .A2(new_n344), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n306), .A2(new_n331), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n352), .A2(new_n320), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n314), .A2(new_n353), .ZN(new_n354));
  NOR3_X1   g168(.A1(new_n334), .A2(KEYINPUT29), .A3(new_n335), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n355), .A2(new_n320), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n305), .A2(new_n300), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n357), .B1(new_n332), .B2(new_n333), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n358), .A2(KEYINPUT29), .ZN(new_n359));
  OAI221_X1 g173(.A(new_n188), .B1(KEYINPUT29), .B2(new_n354), .C1(new_n356), .C2(new_n359), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n349), .A2(new_n351), .B1(G472), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n240), .B1(new_n345), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n221), .A3(G214), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n242), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n316), .A2(G143), .A3(G214), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n264), .A3(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT88), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G131), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT17), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n365), .A2(KEYINPUT88), .A3(new_n264), .A4(new_n366), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n369), .A2(new_n371), .A3(new_n372), .A4(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n370), .A2(KEYINPUT17), .A3(G131), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n374), .A2(new_n205), .A3(new_n213), .A4(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G113), .B(G122), .ZN(new_n377));
  XOR2_X1   g191(.A(new_n377), .B(G104), .Z(new_n378));
  NAND4_X1  g192(.A1(new_n370), .A2(KEYINPUT87), .A3(KEYINPUT18), .A4(G131), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n204), .A2(G146), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n208), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT87), .A2(KEYINPUT18), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n365), .B(new_n366), .C1(new_n264), .C2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n376), .A2(new_n378), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n369), .A2(new_n371), .A3(new_n373), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n206), .A2(KEYINPUT19), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n206), .A2(KEYINPUT19), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n207), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n205), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n378), .B1(new_n391), .B2(new_n384), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT89), .B1(new_n386), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(G475), .A2(G902), .ZN(new_n394));
  INV_X1    g208(.A(new_n392), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT89), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n396), .A3(new_n385), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT20), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n385), .ZN(new_n400));
  NOR3_X1   g214(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT90), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT90), .ZN(new_n403));
  INV_X1    g217(.A(new_n401), .ZN(new_n404));
  AOI211_X1 g218(.A(new_n403), .B(new_n404), .C1(new_n395), .C2(new_n385), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G475), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n378), .B1(new_n376), .B2(new_n384), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(KEYINPUT91), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n385), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n409), .B2(KEYINPUT91), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT92), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n407), .A2(KEYINPUT92), .A3(new_n414), .ZN(new_n418));
  INV_X1    g232(.A(G107), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n289), .A2(G122), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT93), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n289), .A2(G122), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n420), .B2(new_n421), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n419), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n192), .A2(G143), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n242), .A2(G128), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(new_n260), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n420), .A2(new_n424), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n419), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n426), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT94), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n431), .B(new_n419), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n429), .A2(new_n260), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n427), .A2(KEYINPUT13), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n427), .A2(KEYINPUT13), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n438), .A2(new_n439), .A3(new_n428), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n436), .B(new_n437), .C1(new_n260), .C2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT9), .B(G234), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n187), .A2(G953), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n434), .A2(new_n435), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n441), .B(new_n443), .C1(new_n426), .C2(new_n433), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(KEYINPUT94), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n441), .B1(new_n426), .B2(new_n433), .ZN(new_n447));
  INV_X1    g261(.A(new_n443), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n188), .ZN(new_n451));
  INV_X1    g265(.A(G478), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(KEYINPUT15), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n451), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n417), .A2(new_n418), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(G952), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(G953), .ZN(new_n458));
  NAND2_X1  g272(.A1(G234), .A2(G237), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(G902), .A3(G953), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT21), .B(G898), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G214), .B1(G237), .B2(G902), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n467), .B(KEYINPUT84), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n281), .A2(G125), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n469), .B1(G125), .B2(new_n254), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n221), .A2(G224), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT7), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n470), .B(new_n472), .Z(new_n473));
  XNOR2_X1  g287(.A(G110), .B(G122), .ZN(new_n474));
  XOR2_X1   g288(.A(new_n474), .B(KEYINPUT8), .Z(new_n475));
  NAND2_X1  g289(.A1(KEYINPUT78), .A2(G104), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(KEYINPUT78), .A2(G104), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n419), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT3), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT3), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n419), .A3(G104), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT79), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT79), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n484), .A2(new_n481), .A3(new_n419), .A4(G104), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G101), .ZN(new_n487));
  OR2_X1    g301(.A1(KEYINPUT78), .A2(G104), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(G107), .A3(new_n476), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n480), .A2(new_n486), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(G107), .B1(new_n488), .B2(new_n476), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n419), .A2(G104), .ZN(new_n492));
  OAI21_X1  g306(.A(G101), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n288), .A2(new_n290), .A3(KEYINPUT5), .ZN(new_n495));
  OAI21_X1  g309(.A(G113), .B1(new_n288), .B2(KEYINPUT5), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n294), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n497), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n475), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n473), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n489), .B1(new_n491), .B2(new_n481), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n483), .A2(new_n485), .ZN(new_n503));
  OAI21_X1  g317(.A(G101), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(KEYINPUT4), .A3(new_n490), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT4), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n506), .B(G101), .C1(new_n502), .C2(new_n503), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(new_n300), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n474), .A3(new_n498), .ZN(new_n509));
  AOI21_X1  g323(.A(G902), .B1(new_n501), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n498), .ZN(new_n511));
  INV_X1    g325(.A(new_n474), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT6), .A3(new_n509), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n471), .B(KEYINPUT85), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n470), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT6), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n511), .A2(new_n517), .A3(new_n512), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n510), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(G210), .B1(G237), .B2(G902), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(KEYINPUT86), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n522), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n524), .B1(new_n510), .B2(new_n519), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n466), .B(new_n468), .C1(new_n523), .C2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n456), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(G221), .B1(new_n442), .B2(G902), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n494), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(new_n303), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n245), .A2(new_n246), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n207), .A2(G143), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n192), .B1(new_n533), .B2(KEYINPUT1), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(KEYINPUT81), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT81), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n538), .B1(new_n247), .B2(new_n535), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n301), .A3(new_n539), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n540), .A2(new_n490), .A3(new_n493), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n277), .B1(new_n531), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT12), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(KEYINPUT12), .B(new_n277), .C1(new_n531), .C2(new_n541), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n505), .A2(new_n281), .A3(new_n507), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT80), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n505), .A2(KEYINPUT80), .A3(new_n281), .A4(new_n507), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n277), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n530), .A2(KEYINPUT82), .A3(KEYINPUT10), .A4(new_n303), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT82), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n303), .A2(KEYINPUT10), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(new_n494), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n530), .A2(new_n540), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT10), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n553), .A2(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n551), .A2(new_n552), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n546), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(G110), .B(G140), .ZN(new_n562));
  INV_X1    g376(.A(G227), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(G953), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n562), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n551), .A2(new_n559), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n277), .ZN(new_n568));
  INV_X1    g382(.A(new_n565), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n560), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT83), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n566), .A2(new_n570), .A3(KEYINPUT83), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(G469), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G469), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(new_n188), .ZN(new_n577));
  INV_X1    g391(.A(new_n560), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n552), .B1(new_n551), .B2(new_n559), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n565), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n546), .A2(new_n560), .A3(new_n569), .ZN(new_n581));
  AOI21_X1  g395(.A(G902), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n577), .B1(new_n582), .B2(new_n576), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n529), .B1(new_n575), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n527), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n362), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  AOI21_X1  g401(.A(new_n350), .B1(new_n348), .B2(new_n341), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n349), .A2(new_n188), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n589), .B2(G472), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n584), .A2(new_n239), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n590), .A2(KEYINPUT95), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n348), .B2(new_n341), .ZN(new_n595));
  INV_X1    g409(.A(G472), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n343), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n594), .B1(new_n597), .B2(new_n591), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n417), .A2(new_n418), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n450), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n449), .A2(KEYINPUT33), .A3(new_n445), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n604), .A2(G478), .A3(new_n188), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n451), .A2(new_n452), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n520), .A2(new_n521), .ZN(new_n609));
  INV_X1    g423(.A(new_n521), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n510), .A2(new_n610), .A3(new_n519), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n467), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n466), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n599), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT96), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT34), .B(G104), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  NAND2_X1  g433(.A1(new_n393), .A2(new_n397), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n399), .B1(new_n620), .B2(new_n404), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n454), .A2(new_n621), .A3(new_n414), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n599), .A2(new_n466), .A3(new_n613), .A4(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NOR2_X1   g440(.A1(new_n225), .A2(KEYINPUT36), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n220), .B(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n237), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n233), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n527), .A2(new_n584), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n590), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  NAND2_X1  g449(.A1(new_n575), .A2(new_n583), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n631), .A2(new_n609), .A3(new_n467), .A4(new_n611), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(G900), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n461), .B1(new_n463), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n622), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n636), .A2(new_n638), .A3(new_n528), .A4(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n349), .A2(new_n351), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n360), .A2(G472), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n588), .A2(KEYINPUT32), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT97), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n345), .A2(new_n361), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n651), .A3(new_n643), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  NAND2_X1  g468(.A1(new_n353), .A2(new_n357), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n188), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n320), .B1(new_n314), .B2(new_n352), .ZN(new_n657));
  OAI21_X1  g471(.A(G472), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n644), .B(new_n658), .C1(KEYINPUT32), .C2(new_n588), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT98), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n640), .B(KEYINPUT39), .Z(new_n661));
  NAND2_X1  g475(.A1(new_n584), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(KEYINPUT40), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n523), .A2(new_n525), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT38), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT92), .B1(new_n407), .B2(new_n414), .ZN(new_n667));
  AOI211_X1 g481(.A(new_n416), .B(new_n413), .C1(new_n399), .C2(new_n406), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n631), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n454), .A3(new_n467), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n666), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n660), .A2(new_n663), .A3(new_n664), .A4(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT99), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G143), .ZN(G45));
  INV_X1    g489(.A(new_n640), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n607), .B(new_n676), .C1(new_n667), .C2(new_n668), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n678), .A2(new_n584), .A3(new_n638), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n650), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n207), .ZN(G48));
  AOI21_X1  g495(.A(new_n569), .B1(new_n568), .B2(new_n560), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n546), .A2(new_n560), .A3(new_n569), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n188), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G469), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n576), .B(new_n188), .C1(new_n682), .C2(new_n683), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n528), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n362), .A2(new_n615), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NOR2_X1   g505(.A1(new_n614), .A2(new_n687), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n362), .A2(new_n623), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G116), .ZN(G18));
  NOR2_X1   g508(.A1(new_n687), .A2(new_n637), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n456), .A2(new_n465), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n650), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  INV_X1    g512(.A(KEYINPUT100), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n358), .A2(new_n320), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n323), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n701), .A2(new_n329), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n323), .A2(new_n700), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT100), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n241), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n706), .B1(new_n595), .B2(new_n596), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n669), .A2(new_n455), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n239), .A3(new_n692), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NAND2_X1  g525(.A1(new_n695), .A2(new_n678), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT101), .B1(new_n707), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n589), .A2(G472), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT101), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n677), .A2(new_n687), .A3(new_n637), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n714), .A2(new_n715), .A3(new_n706), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n720));
  INV_X1    g534(.A(new_n467), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n523), .A2(new_n525), .A3(new_n721), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n560), .A2(new_n569), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n723), .A2(new_n568), .B1(new_n561), .B2(new_n565), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n577), .B1(new_n724), .B2(G469), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n529), .B1(new_n725), .B2(new_n686), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT102), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n722), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI211_X1 g542(.A(KEYINPUT102), .B(new_n529), .C1(new_n725), .C2(new_n686), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n728), .A2(new_n677), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n362), .A2(KEYINPUT42), .A3(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT42), .B1(new_n362), .B2(new_n730), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n720), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n650), .A2(new_n239), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n728), .A2(new_n729), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n678), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n731), .A3(KEYINPUT103), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G131), .ZN(G33));
  INV_X1    g556(.A(new_n641), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n728), .A2(new_n743), .A3(new_n729), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n362), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  AOI21_X1  g560(.A(KEYINPUT45), .B1(new_n573), .B2(new_n574), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n576), .B(new_n747), .C1(KEYINPUT45), .C2(new_n724), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n577), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  OR3_X1    g564(.A1(new_n749), .A2(new_n750), .A3(KEYINPUT46), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n750), .B1(new_n749), .B2(KEYINPUT46), .ZN(new_n752));
  INV_X1    g566(.A(new_n686), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n753), .B1(new_n749), .B2(KEYINPUT46), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n528), .A3(new_n661), .ZN(new_n756));
  INV_X1    g570(.A(new_n722), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n669), .A2(new_n607), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n758), .B(KEYINPUT43), .Z(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n597), .A3(new_n631), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n756), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(new_n256), .ZN(G39));
  NAND2_X1  g579(.A1(new_n755), .A2(new_n528), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(KEYINPUT47), .ZN(new_n767));
  INV_X1    g581(.A(new_n650), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n240), .A3(new_n678), .A4(new_n722), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n202), .ZN(G42));
  NAND2_X1  g585(.A1(new_n759), .A2(new_n461), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n772), .B(KEYINPUT109), .Z(new_n773));
  NOR2_X1   g587(.A1(new_n757), .A2(new_n687), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n362), .A3(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT48), .Z(new_n776));
  INV_X1    g590(.A(new_n660), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n239), .A3(new_n461), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n708), .A2(new_n239), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n773), .A2(new_n688), .A3(new_n780), .ZN(new_n781));
  OAI221_X1 g595(.A(new_n458), .B1(new_n608), .B2(new_n778), .C1(new_n781), .C2(new_n612), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n776), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n773), .A2(new_n631), .A3(new_n708), .A4(new_n774), .ZN(new_n784));
  OR3_X1    g598(.A1(new_n778), .A2(new_n600), .A3(new_n607), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n666), .A2(new_n721), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n786), .B1(new_n781), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n784), .B(new_n785), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g606(.A(KEYINPUT108), .B(KEYINPUT51), .Z(new_n793));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n685), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(new_n753), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n529), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n767), .A2(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n773), .A2(new_n780), .A3(new_n722), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n795), .B1(new_n801), .B2(KEYINPUT51), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n783), .B1(new_n792), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n767), .A2(KEYINPUT110), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n798), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n767), .A2(KEYINPUT110), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n800), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n794), .B1(new_n790), .B2(new_n791), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n793), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT106), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n726), .A2(new_n670), .A3(new_n676), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n600), .A2(new_n613), .A3(new_n454), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n650), .A2(new_n679), .B1(new_n659), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g630(.A(KEYINPUT97), .B(new_n642), .C1(new_n345), .C2(new_n361), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n651), .B1(new_n650), .B2(new_n643), .ZN(new_n818));
  OAI211_X1 g632(.A(new_n816), .B(new_n718), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n653), .A2(KEYINPUT52), .A3(new_n718), .A4(new_n816), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(KEYINPUT105), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT105), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n819), .A2(new_n824), .A3(new_n820), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n456), .B1(new_n669), .B2(new_n607), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n526), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n593), .A2(new_n598), .A3(new_n828), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n362), .A2(new_n585), .B1(new_n632), .B2(new_n590), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n454), .A2(new_n413), .A3(new_n640), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n831), .A2(new_n621), .A3(new_n631), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n832), .A2(new_n584), .A3(new_n722), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n362), .A2(new_n744), .B1(new_n650), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n730), .A2(new_n708), .A3(new_n631), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n829), .A2(new_n830), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n689), .A2(new_n693), .A3(new_n697), .A4(new_n710), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n734), .A3(new_n740), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n812), .B1(new_n826), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n838), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n821), .A2(new_n822), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n840), .A2(KEYINPUT53), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n811), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n842), .A2(new_n811), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT54), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n821), .A2(new_n822), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n812), .B1(new_n846), .B2(new_n838), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT107), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n829), .A2(new_n830), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n834), .A2(new_n835), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n650), .A2(new_n833), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n745), .A2(new_n835), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT107), .A3(new_n829), .A4(new_n830), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n812), .B1(new_n739), .B2(new_n731), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n856), .A2(new_n837), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n855), .A2(new_n823), .A3(new_n825), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n847), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n845), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g675(.A1(new_n810), .A2(new_n861), .B1(new_n457), .B2(new_n221), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n666), .A2(new_n239), .A3(new_n528), .A4(new_n468), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT49), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n797), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n796), .A2(new_n753), .A3(KEYINPUT49), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n865), .A2(new_n758), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n660), .A2(new_n863), .A3(new_n867), .ZN(new_n868));
  OR2_X1    g682(.A1(new_n862), .A2(new_n868), .ZN(G75));
  NOR2_X1   g683(.A1(new_n221), .A2(G952), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT116), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n188), .B1(new_n847), .B2(new_n858), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(G210), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT114), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n514), .A2(new_n518), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n516), .ZN(new_n879));
  XNOR2_X1  g693(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n879), .B(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT56), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT114), .B1(new_n881), .B2(KEYINPUT115), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n875), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n872), .B1(new_n882), .B2(new_n885), .ZN(G51));
  NAND2_X1  g700(.A1(new_n847), .A2(new_n858), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT54), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n860), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n577), .B(KEYINPUT57), .Z(new_n891));
  OAI22_X1  g705(.A1(new_n890), .A2(new_n891), .B1(new_n682), .B2(new_n683), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n874), .A2(new_n748), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n870), .B1(new_n892), .B2(new_n893), .ZN(G54));
  NAND3_X1  g708(.A1(new_n874), .A2(KEYINPUT58), .A3(G475), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n870), .B1(new_n895), .B2(new_n620), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n896), .B1(new_n620), .B2(new_n895), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT117), .Z(G60));
  INV_X1    g712(.A(new_n604), .ZN(new_n899));
  XNOR2_X1  g713(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n900));
  NAND2_X1  g714(.A1(G478), .A2(G902), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n900), .B(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n847), .A2(new_n859), .A3(new_n858), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n859), .B1(new_n847), .B2(new_n858), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT119), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n908), .B(new_n903), .C1(new_n904), .C2(new_n905), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n872), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n902), .B1(new_n845), .B2(new_n860), .ZN(new_n911));
  OAI22_X1  g725(.A1(new_n910), .A2(KEYINPUT120), .B1(new_n604), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n913), .B(new_n872), .C1(new_n907), .C2(new_n909), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT121), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n908), .B1(new_n889), .B2(new_n903), .ZN(new_n916));
  INV_X1    g730(.A(new_n909), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n871), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n913), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n910), .A2(KEYINPUT120), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n899), .B1(new_n861), .B2(new_n902), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n915), .A2(new_n923), .ZN(G63));
  NAND2_X1  g738(.A1(G217), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT60), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n847), .B2(new_n858), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n628), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n872), .B1(KEYINPUT122), .B2(new_n929), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n928), .B(new_n930), .C1(new_n229), .C2(new_n927), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n929), .A2(KEYINPUT122), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n931), .B(new_n932), .Z(G66));
  NAND3_X1  g747(.A1(new_n837), .A2(new_n829), .A3(new_n830), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n221), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT123), .Z(new_n936));
  INV_X1    g750(.A(G224), .ZN(new_n937));
  OAI21_X1  g751(.A(G953), .B1(new_n464), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n878), .B1(G898), .B2(new_n221), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G69));
  NOR4_X1   g755(.A1(new_n736), .A2(new_n662), .A3(new_n757), .A4(new_n827), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n770), .A2(new_n764), .A3(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n653), .ZN(new_n944));
  INV_X1    g758(.A(new_n718), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n944), .A2(new_n680), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n674), .A2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(KEYINPUT62), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n943), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n221), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n287), .A2(new_n307), .A3(new_n313), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n388), .A2(new_n389), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT124), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(G900), .A2(G953), .ZN(new_n957));
  INV_X1    g771(.A(new_n770), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n756), .A2(new_n814), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n362), .B1(new_n959), .B2(new_n744), .ZN(new_n960));
  INV_X1    g774(.A(new_n946), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n764), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n958), .A2(new_n741), .A3(new_n960), .A4(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n957), .B(new_n954), .C1(new_n963), .C2(G953), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n956), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(G953), .B1(new_n563), .B2(new_n639), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT126), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n965), .A2(new_n969), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n971), .ZN(G72));
  XNOR2_X1  g786(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n596), .A2(new_n188), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n973), .B(new_n974), .Z(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n950), .B2(new_n934), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n657), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n976), .B1(new_n963), .B2(new_n934), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n314), .A2(new_n353), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n870), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n843), .A2(new_n844), .ZN(new_n983));
  NOR3_X1   g797(.A1(new_n980), .A2(new_n657), .A3(new_n975), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(G57));
endmodule


