

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742;

  OR2_X1 U370 ( .A1(n549), .A2(n675), .ZN(n559) );
  AND2_X2 U371 ( .A1(n556), .A2(n352), .ZN(n670) );
  NOR2_X2 U372 ( .A1(n698), .A2(n520), .ZN(n460) );
  XNOR2_X2 U373 ( .A(n434), .B(n435), .ZN(n698) );
  XNOR2_X2 U374 ( .A(n489), .B(n488), .ZN(n523) );
  NOR2_X1 U375 ( .A1(n688), .A2(n597), .ZN(n598) );
  INV_X1 U376 ( .A(n559), .ZN(n678) );
  XNOR2_X1 U377 ( .A(n406), .B(KEYINPUT25), .ZN(n549) );
  XNOR2_X1 U378 ( .A(KEYINPUT4), .B(G146), .ZN(n380) );
  AND2_X1 U379 ( .A1(n620), .A2(n542), .ZN(n610) );
  AND2_X1 U380 ( .A1(n533), .A2(n532), .ZN(n540) );
  AND2_X1 U381 ( .A1(n507), .A2(n506), .ZN(n513) );
  XNOR2_X1 U382 ( .A(n460), .B(KEYINPUT34), .ZN(n351) );
  NOR2_X1 U383 ( .A1(n603), .A2(n553), .ZN(n554) );
  BUF_X1 U384 ( .A(n567), .Z(n607) );
  XNOR2_X1 U385 ( .A(n363), .B(G472), .ZN(n573) );
  OR2_X1 U386 ( .A1(n630), .A2(G902), .ZN(n421) );
  XNOR2_X1 U387 ( .A(n380), .B(KEYINPUT64), .ZN(n379) );
  XNOR2_X1 U388 ( .A(G143), .B(G131), .ZN(n476) );
  XNOR2_X1 U389 ( .A(G104), .B(G122), .ZN(n475) );
  INV_X1 U390 ( .A(n495), .ZN(n534) );
  XNOR2_X2 U391 ( .A(n350), .B(n349), .ZN(n495) );
  INV_X1 U392 ( .A(n494), .ZN(n349) );
  NAND2_X1 U393 ( .A1(n351), .A2(n492), .ZN(n350) );
  INV_X1 U394 ( .A(n555), .ZN(n352) );
  XNOR2_X1 U395 ( .A(n577), .B(n422), .ZN(n499) );
  XNOR2_X1 U396 ( .A(n353), .B(KEYINPUT110), .ZN(n592) );
  AND2_X1 U397 ( .A1(n524), .A2(n525), .ZN(n353) );
  XNOR2_X1 U398 ( .A(G137), .B(KEYINPUT23), .ZN(n391) );
  INV_X1 U399 ( .A(KEYINPUT46), .ZN(n376) );
  NOR2_X1 U400 ( .A1(n587), .A2(n378), .ZN(n377) );
  NOR2_X1 U401 ( .A1(n592), .A2(n609), .ZN(n694) );
  XNOR2_X1 U402 ( .A(n449), .B(n448), .ZN(n567) );
  INV_X1 U403 ( .A(n573), .ZN(n681) );
  XNOR2_X1 U404 ( .A(G113), .B(G119), .ZN(n423) );
  XOR2_X1 U405 ( .A(KEYINPUT74), .B(KEYINPUT3), .Z(n424) );
  NAND2_X2 U406 ( .A1(n620), .A2(n384), .ZN(n361) );
  XNOR2_X1 U407 ( .A(n619), .B(KEYINPUT91), .ZN(n384) );
  XNOR2_X1 U408 ( .A(G116), .B(KEYINPUT105), .ZN(n426) );
  XOR2_X1 U409 ( .A(KEYINPUT5), .B(KEYINPUT77), .Z(n427) );
  XNOR2_X1 U410 ( .A(KEYINPUT71), .B(KEYINPUT10), .ZN(n398) );
  XNOR2_X1 U411 ( .A(G113), .B(KEYINPUT12), .ZN(n479) );
  XOR2_X1 U412 ( .A(KEYINPUT106), .B(KEYINPUT11), .Z(n480) );
  XNOR2_X1 U413 ( .A(G131), .B(G134), .ZN(n414) );
  XNOR2_X1 U414 ( .A(n364), .B(KEYINPUT72), .ZN(n415) );
  INV_X1 U415 ( .A(G137), .ZN(n364) );
  OR2_X1 U416 ( .A1(n577), .A2(n558), .ZN(n560) );
  XOR2_X1 U417 ( .A(G116), .B(G122), .Z(n462) );
  INV_X1 U418 ( .A(G119), .ZN(n399) );
  XNOR2_X1 U419 ( .A(G128), .B(G110), .ZN(n389) );
  AND2_X1 U420 ( .A1(n361), .A2(G475), .ZN(n370) );
  XNOR2_X1 U421 ( .A(n446), .B(n445), .ZN(n623) );
  INV_X1 U422 ( .A(KEYINPUT48), .ZN(n373) );
  NAND2_X1 U423 ( .A1(n377), .A2(n375), .ZN(n374) );
  XNOR2_X1 U424 ( .A(n599), .B(n376), .ZN(n375) );
  XNOR2_X1 U425 ( .A(n591), .B(n590), .ZN(n608) );
  INV_X1 U426 ( .A(KEYINPUT39), .ZN(n590) );
  NAND2_X1 U427 ( .A1(n645), .A2(n472), .ZN(n363) );
  XNOR2_X1 U428 ( .A(n592), .B(KEYINPUT116), .ZN(n654) );
  XNOR2_X1 U429 ( .A(n573), .B(n362), .ZN(n551) );
  INV_X1 U430 ( .A(KEYINPUT6), .ZN(n362) );
  AND2_X1 U431 ( .A1(n361), .A2(G472), .ZN(n371) );
  AND2_X1 U432 ( .A1(n361), .A2(G469), .ZN(n369) );
  AND2_X1 U433 ( .A1(n361), .A2(G210), .ZN(n368) );
  NOR2_X1 U434 ( .A1(n736), .A2(G952), .ZN(n714) );
  XOR2_X1 U435 ( .A(KEYINPUT42), .B(n598), .Z(n741) );
  NAND2_X1 U436 ( .A1(n367), .A2(n366), .ZN(n706) );
  NOR2_X1 U437 ( .A1(n705), .A2(n355), .ZN(n366) );
  NOR2_X1 U438 ( .A1(n681), .A2(n517), .ZN(n354) );
  OR2_X1 U439 ( .A1(G953), .A2(n674), .ZN(n355) );
  XOR2_X1 U440 ( .A(G125), .B(G140), .Z(n356) );
  XNOR2_X1 U441 ( .A(KEYINPUT76), .B(n602), .ZN(n357) );
  OR2_X1 U442 ( .A1(n704), .A2(KEYINPUT2), .ZN(n358) );
  NOR2_X1 U443 ( .A1(n613), .A2(n611), .ZN(n359) );
  NOR2_X1 U444 ( .A1(n359), .A2(n615), .ZN(n360) );
  AND2_X1 U445 ( .A1(n385), .A2(n361), .ZN(n372) );
  NAND2_X1 U446 ( .A1(n358), .A2(n361), .ZN(n367) );
  XNOR2_X2 U447 ( .A(n365), .B(n413), .ZN(n446) );
  XNOR2_X1 U448 ( .A(n432), .B(n365), .ZN(n645) );
  XNOR2_X2 U449 ( .A(n728), .B(n411), .ZN(n365) );
  NOR2_X1 U450 ( .A1(n648), .A2(n714), .ZN(n651) );
  NAND2_X1 U451 ( .A1(n371), .A2(n385), .ZN(n647) );
  XNOR2_X2 U452 ( .A(n461), .B(n379), .ZN(n728) );
  NAND2_X1 U453 ( .A1(n368), .A2(n385), .ZN(n625) );
  NAND2_X1 U454 ( .A1(n369), .A2(n385), .ZN(n632) );
  NAND2_X1 U455 ( .A1(n370), .A2(n385), .ZN(n637) );
  NAND2_X1 U456 ( .A1(n372), .A2(G478), .ZN(n709) );
  NAND2_X1 U457 ( .A1(n372), .A2(G217), .ZN(n712) );
  XNOR2_X2 U458 ( .A(n374), .B(n373), .ZN(n618) );
  NAND2_X1 U459 ( .A1(n357), .A2(n588), .ZN(n378) );
  XNOR2_X2 U460 ( .A(n382), .B(n381), .ZN(n461) );
  XNOR2_X2 U461 ( .A(KEYINPUT65), .B(KEYINPUT84), .ZN(n381) );
  XNOR2_X2 U462 ( .A(G143), .B(G128), .ZN(n382) );
  NAND2_X2 U463 ( .A1(n383), .A2(n360), .ZN(n385) );
  NAND2_X1 U464 ( .A1(n610), .A2(n734), .ZN(n383) );
  XOR2_X1 U465 ( .A(n606), .B(KEYINPUT43), .Z(n386) );
  XOR2_X1 U466 ( .A(n636), .B(n635), .Z(n387) );
  XNOR2_X1 U467 ( .A(KEYINPUT89), .B(n694), .ZN(n388) );
  INV_X1 U468 ( .A(KEYINPUT87), .ZN(n585) );
  INV_X1 U469 ( .A(n675), .ZN(n410) );
  XNOR2_X1 U470 ( .A(n486), .B(n399), .ZN(n400) );
  XNOR2_X1 U471 ( .A(n401), .B(n400), .ZN(n711) );
  XOR2_X1 U472 ( .A(n523), .B(KEYINPUT107), .Z(n525) );
  XOR2_X1 U473 ( .A(KEYINPUT114), .B(KEYINPUT33), .Z(n435) );
  XOR2_X1 U474 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n390) );
  XNOR2_X1 U475 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U476 ( .A(KEYINPUT79), .B(KEYINPUT24), .Z(n392) );
  XNOR2_X1 U477 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U478 ( .A(n394), .B(n393), .Z(n397) );
  INV_X2 U479 ( .A(G953), .ZN(n736) );
  NAND2_X1 U480 ( .A1(G234), .A2(n736), .ZN(n395) );
  XOR2_X1 U481 ( .A(KEYINPUT8), .B(n395), .Z(n468) );
  NAND2_X1 U482 ( .A1(n468), .A2(G221), .ZN(n396) );
  XNOR2_X1 U483 ( .A(n397), .B(n396), .ZN(n401) );
  XNOR2_X1 U484 ( .A(n356), .B(n398), .ZN(n727) );
  XNOR2_X1 U485 ( .A(n727), .B(G146), .ZN(n486) );
  NOR2_X1 U486 ( .A1(G902), .A2(n711), .ZN(n405) );
  XNOR2_X1 U487 ( .A(G902), .B(KEYINPUT98), .ZN(n402) );
  XNOR2_X1 U488 ( .A(n402), .B(KEYINPUT15), .ZN(n613) );
  NAND2_X1 U489 ( .A1(n613), .A2(G234), .ZN(n403) );
  XNOR2_X1 U490 ( .A(n403), .B(KEYINPUT20), .ZN(n407) );
  AND2_X1 U491 ( .A1(G217), .A2(n407), .ZN(n404) );
  XNOR2_X1 U492 ( .A(n405), .B(n404), .ZN(n406) );
  AND2_X1 U493 ( .A1(n407), .A2(G221), .ZN(n409) );
  INV_X1 U494 ( .A(KEYINPUT21), .ZN(n408) );
  XNOR2_X1 U495 ( .A(n409), .B(n408), .ZN(n675) );
  XNOR2_X1 U496 ( .A(KEYINPUT69), .B(G101), .ZN(n411) );
  XNOR2_X1 U497 ( .A(G110), .B(G107), .ZN(n412) );
  XNOR2_X1 U498 ( .A(n412), .B(G104), .ZN(n715) );
  XNOR2_X1 U499 ( .A(n715), .B(KEYINPUT75), .ZN(n413) );
  XNOR2_X1 U500 ( .A(n415), .B(n414), .ZN(n429) );
  XOR2_X1 U501 ( .A(n429), .B(KEYINPUT101), .Z(n730) );
  XOR2_X1 U502 ( .A(G140), .B(KEYINPUT80), .Z(n417) );
  NAND2_X1 U503 ( .A1(G227), .A2(n736), .ZN(n416) );
  XNOR2_X1 U504 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U505 ( .A(n730), .B(n418), .ZN(n419) );
  XNOR2_X1 U506 ( .A(n446), .B(n419), .ZN(n630) );
  INV_X1 U507 ( .A(G469), .ZN(n420) );
  XNOR2_X2 U508 ( .A(n421), .B(n420), .ZN(n577) );
  INV_X1 U509 ( .A(KEYINPUT1), .ZN(n422) );
  NAND2_X1 U510 ( .A1(n678), .A2(n499), .ZN(n517) );
  INV_X1 U511 ( .A(n517), .ZN(n433) );
  XNOR2_X1 U512 ( .A(n424), .B(n423), .ZN(n436) );
  NOR2_X1 U513 ( .A1(G953), .A2(G237), .ZN(n483) );
  AND2_X1 U514 ( .A1(n483), .A2(G210), .ZN(n425) );
  XNOR2_X1 U515 ( .A(n436), .B(n425), .ZN(n431) );
  XNOR2_X1 U516 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U517 ( .A(n429), .B(n428), .Z(n430) );
  XNOR2_X1 U518 ( .A(n431), .B(n430), .ZN(n432) );
  INV_X1 U519 ( .A(G902), .ZN(n472) );
  NAND2_X1 U520 ( .A1(n433), .A2(n551), .ZN(n434) );
  XNOR2_X1 U521 ( .A(n462), .B(KEYINPUT16), .ZN(n437) );
  XNOR2_X1 U522 ( .A(n437), .B(n436), .ZN(n716) );
  XOR2_X1 U523 ( .A(G125), .B(KEYINPUT96), .Z(n439) );
  XOR2_X1 U524 ( .A(KEYINPUT18), .B(KEYINPUT99), .Z(n438) );
  XNOR2_X1 U525 ( .A(n439), .B(n438), .ZN(n443) );
  XNOR2_X1 U526 ( .A(KEYINPUT81), .B(KEYINPUT17), .ZN(n441) );
  NAND2_X1 U527 ( .A1(G224), .A2(n736), .ZN(n440) );
  XNOR2_X1 U528 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U529 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U530 ( .A(n716), .B(n444), .ZN(n445) );
  NAND2_X1 U531 ( .A1(n623), .A2(n613), .ZN(n449) );
  INV_X1 U532 ( .A(G237), .ZN(n447) );
  NAND2_X1 U533 ( .A1(n472), .A2(n447), .ZN(n450) );
  NAND2_X1 U534 ( .A1(n450), .A2(G210), .ZN(n448) );
  INV_X1 U535 ( .A(n567), .ZN(n451) );
  NAND2_X1 U536 ( .A1(n450), .A2(G214), .ZN(n689) );
  NAND2_X1 U537 ( .A1(n451), .A2(n689), .ZN(n553) );
  XNOR2_X1 U538 ( .A(KEYINPUT67), .B(KEYINPUT19), .ZN(n452) );
  XNOR2_X1 U539 ( .A(n553), .B(n452), .ZN(n580) );
  NAND2_X1 U540 ( .A1(G234), .A2(G237), .ZN(n453) );
  XNOR2_X1 U541 ( .A(KEYINPUT14), .B(n453), .ZN(n455) );
  NAND2_X1 U542 ( .A1(G952), .A2(n455), .ZN(n703) );
  NOR2_X1 U543 ( .A1(G953), .A2(n703), .ZN(n454) );
  XNOR2_X1 U544 ( .A(n454), .B(KEYINPUT100), .ZN(n547) );
  NOR2_X1 U545 ( .A1(G898), .A2(n736), .ZN(n718) );
  INV_X1 U546 ( .A(n718), .ZN(n456) );
  NAND2_X1 U547 ( .A1(G902), .A2(n455), .ZN(n543) );
  NOR2_X1 U548 ( .A1(n456), .A2(n543), .ZN(n457) );
  NOR2_X1 U549 ( .A1(n547), .A2(n457), .ZN(n458) );
  NOR2_X2 U550 ( .A1(n580), .A2(n458), .ZN(n459) );
  XNOR2_X2 U551 ( .A(n459), .B(KEYINPUT0), .ZN(n516) );
  INV_X1 U552 ( .A(n516), .ZN(n520) );
  XNOR2_X1 U553 ( .A(KEYINPUT109), .B(KEYINPUT108), .ZN(n463) );
  XNOR2_X1 U554 ( .A(n463), .B(n462), .ZN(n467) );
  XOR2_X1 U555 ( .A(G107), .B(KEYINPUT9), .Z(n465) );
  XNOR2_X1 U556 ( .A(G134), .B(KEYINPUT7), .ZN(n464) );
  XNOR2_X1 U557 ( .A(n465), .B(n464), .ZN(n466) );
  XOR2_X1 U558 ( .A(n467), .B(n466), .Z(n470) );
  NAND2_X1 U559 ( .A1(G217), .A2(n468), .ZN(n469) );
  XNOR2_X1 U560 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U561 ( .A(n461), .B(n471), .ZN(n707) );
  NAND2_X1 U562 ( .A1(n707), .A2(n472), .ZN(n474) );
  INV_X1 U563 ( .A(G478), .ZN(n473) );
  XNOR2_X1 U564 ( .A(n474), .B(n473), .ZN(n524) );
  INV_X1 U565 ( .A(n524), .ZN(n490) );
  INV_X1 U566 ( .A(n475), .ZN(n477) );
  XNOR2_X1 U567 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U568 ( .A(n478), .ZN(n482) );
  XNOR2_X1 U569 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U570 ( .A(n482), .B(n481), .ZN(n485) );
  NAND2_X1 U571 ( .A1(G214), .A2(n483), .ZN(n484) );
  XNOR2_X1 U572 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U573 ( .A(n487), .B(n486), .ZN(n636) );
  NOR2_X1 U574 ( .A1(n636), .A2(G902), .ZN(n489) );
  XNOR2_X1 U575 ( .A(KEYINPUT13), .B(G475), .ZN(n488) );
  NAND2_X1 U576 ( .A1(n490), .A2(n523), .ZN(n491) );
  XOR2_X1 U577 ( .A(KEYINPUT115), .B(n491), .Z(n566) );
  INV_X1 U578 ( .A(n566), .ZN(n492) );
  INV_X1 U579 ( .A(KEYINPUT82), .ZN(n493) );
  XNOR2_X1 U580 ( .A(n493), .B(KEYINPUT35), .ZN(n494) );
  NAND2_X1 U581 ( .A1(n495), .A2(KEYINPUT94), .ZN(n507) );
  INV_X1 U582 ( .A(n523), .ZN(n496) );
  AND2_X1 U583 ( .A1(n496), .A2(n524), .ZN(n595) );
  AND2_X1 U584 ( .A1(n595), .A2(n410), .ZN(n497) );
  NAND2_X1 U585 ( .A1(n516), .A2(n497), .ZN(n498) );
  XNOR2_X1 U586 ( .A(n498), .B(KEYINPUT22), .ZN(n530) );
  INV_X1 U587 ( .A(n499), .ZN(n555) );
  INV_X1 U588 ( .A(KEYINPUT112), .ZN(n500) );
  XNOR2_X1 U589 ( .A(n549), .B(n500), .ZN(n527) );
  OR2_X1 U590 ( .A1(n551), .A2(n527), .ZN(n501) );
  NOR2_X1 U591 ( .A1(n555), .A2(n501), .ZN(n502) );
  XNOR2_X1 U592 ( .A(n502), .B(KEYINPUT83), .ZN(n503) );
  OR2_X1 U593 ( .A1(n530), .A2(n503), .ZN(n505) );
  INV_X1 U594 ( .A(KEYINPUT32), .ZN(n504) );
  XNOR2_X2 U595 ( .A(n505), .B(n504), .ZN(n740) );
  INV_X1 U596 ( .A(n740), .ZN(n506) );
  AND2_X1 U597 ( .A1(n681), .A2(n549), .ZN(n508) );
  NAND2_X1 U598 ( .A1(n555), .A2(n508), .ZN(n509) );
  OR2_X1 U599 ( .A1(n530), .A2(n509), .ZN(n511) );
  INV_X1 U600 ( .A(KEYINPUT113), .ZN(n510) );
  XNOR2_X2 U601 ( .A(n511), .B(n510), .ZN(n644) );
  AND2_X1 U602 ( .A1(n644), .A2(KEYINPUT44), .ZN(n512) );
  NAND2_X1 U603 ( .A1(n513), .A2(n512), .ZN(n515) );
  INV_X1 U604 ( .A(KEYINPUT44), .ZN(n535) );
  NAND2_X1 U605 ( .A1(n535), .A2(KEYINPUT94), .ZN(n514) );
  NAND2_X1 U606 ( .A1(n515), .A2(n514), .ZN(n533) );
  NAND2_X1 U607 ( .A1(n516), .A2(n354), .ZN(n518) );
  XNOR2_X1 U608 ( .A(n518), .B(KEYINPUT31), .ZN(n668) );
  OR2_X1 U609 ( .A1(n577), .A2(n559), .ZN(n519) );
  NOR2_X1 U610 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U611 ( .A(KEYINPUT104), .B(n521), .Z(n522) );
  NOR2_X1 U612 ( .A1(n573), .A2(n522), .ZN(n656) );
  OR2_X1 U613 ( .A1(n668), .A2(n656), .ZN(n526) );
  NOR2_X1 U614 ( .A1(n525), .A2(n524), .ZN(n667) );
  XOR2_X1 U615 ( .A(KEYINPUT111), .B(n667), .Z(n609) );
  NAND2_X1 U616 ( .A1(n526), .A2(n388), .ZN(n531) );
  INV_X1 U617 ( .A(n527), .ZN(n676) );
  NOR2_X1 U618 ( .A1(n551), .A2(n676), .ZN(n528) );
  NAND2_X1 U619 ( .A1(n555), .A2(n528), .ZN(n529) );
  OR2_X1 U620 ( .A1(n530), .A2(n529), .ZN(n652) );
  AND2_X1 U621 ( .A1(n531), .A2(n652), .ZN(n532) );
  NAND2_X1 U622 ( .A1(n644), .A2(n535), .ZN(n536) );
  OR2_X1 U623 ( .A1(n536), .A2(n740), .ZN(n537) );
  NAND2_X1 U624 ( .A1(n537), .A2(KEYINPUT94), .ZN(n538) );
  NAND2_X1 U625 ( .A1(n534), .A2(n538), .ZN(n539) );
  NAND2_X1 U626 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X2 U627 ( .A(n541), .B(KEYINPUT45), .ZN(n620) );
  INV_X1 U628 ( .A(n613), .ZN(n542) );
  NOR2_X1 U629 ( .A1(G900), .A2(n543), .ZN(n544) );
  NAND2_X1 U630 ( .A1(G953), .A2(n544), .ZN(n545) );
  XNOR2_X1 U631 ( .A(KEYINPUT117), .B(n545), .ZN(n546) );
  NOR2_X1 U632 ( .A1(n547), .A2(n546), .ZN(n558) );
  NOR2_X1 U633 ( .A1(n675), .A2(n558), .ZN(n548) );
  NAND2_X1 U634 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U635 ( .A(KEYINPUT73), .B(n550), .ZN(n574) );
  AND2_X1 U636 ( .A1(n551), .A2(n574), .ZN(n552) );
  NAND2_X1 U637 ( .A1(n552), .A2(n654), .ZN(n603) );
  XNOR2_X1 U638 ( .A(n554), .B(KEYINPUT36), .ZN(n556) );
  XNOR2_X1 U639 ( .A(KEYINPUT93), .B(n670), .ZN(n588) );
  NAND2_X1 U640 ( .A1(n694), .A2(KEYINPUT47), .ZN(n557) );
  XNOR2_X1 U641 ( .A(KEYINPUT88), .B(n557), .ZN(n571) );
  NOR2_X1 U642 ( .A1(n560), .A2(n559), .ZN(n564) );
  XOR2_X1 U643 ( .A(KEYINPUT118), .B(KEYINPUT30), .Z(n562) );
  NAND2_X1 U644 ( .A1(n573), .A2(n689), .ZN(n561) );
  XNOR2_X1 U645 ( .A(n562), .B(n561), .ZN(n563) );
  NAND2_X1 U646 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U647 ( .A(n565), .B(KEYINPUT78), .ZN(n589) );
  NOR2_X1 U648 ( .A1(n589), .A2(n566), .ZN(n569) );
  INV_X1 U649 ( .A(n607), .ZN(n568) );
  NAND2_X1 U650 ( .A1(n569), .A2(n568), .ZN(n642) );
  XNOR2_X1 U651 ( .A(n642), .B(KEYINPUT90), .ZN(n570) );
  NAND2_X1 U652 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U653 ( .A(n572), .B(KEYINPUT85), .ZN(n584) );
  XOR2_X1 U654 ( .A(KEYINPUT28), .B(KEYINPUT119), .Z(n576) );
  NAND2_X1 U655 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U656 ( .A(n576), .B(n575), .Z(n579) );
  INV_X1 U657 ( .A(n577), .ZN(n578) );
  NAND2_X1 U658 ( .A1(n579), .A2(n578), .ZN(n597) );
  INV_X1 U659 ( .A(n597), .ZN(n582) );
  INV_X1 U660 ( .A(n580), .ZN(n581) );
  NAND2_X1 U661 ( .A1(n582), .A2(n581), .ZN(n660) );
  NAND2_X1 U662 ( .A1(n660), .A2(KEYINPUT47), .ZN(n583) );
  NAND2_X1 U663 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U664 ( .A(n586), .B(n585), .ZN(n587) );
  XOR2_X1 U665 ( .A(KEYINPUT38), .B(n607), .Z(n594) );
  NOR2_X1 U666 ( .A1(n589), .A2(n594), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n608), .A2(n592), .ZN(n593) );
  XNOR2_X1 U668 ( .A(n593), .B(KEYINPUT40), .ZN(n742) );
  INV_X1 U669 ( .A(n594), .ZN(n690) );
  NAND2_X1 U670 ( .A1(n690), .A2(n689), .ZN(n693) );
  INV_X1 U671 ( .A(n595), .ZN(n692) );
  NOR2_X1 U672 ( .A1(n693), .A2(n692), .ZN(n596) );
  XNOR2_X1 U673 ( .A(n596), .B(KEYINPUT41), .ZN(n688) );
  NAND2_X1 U674 ( .A1(n742), .A2(n741), .ZN(n599) );
  XNOR2_X1 U675 ( .A(KEYINPUT70), .B(KEYINPUT47), .ZN(n600) );
  NOR2_X1 U676 ( .A1(n660), .A2(n600), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n601), .A2(n388), .ZN(n602) );
  INV_X1 U678 ( .A(n603), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n604), .A2(n689), .ZN(n605) );
  NOR2_X1 U680 ( .A1(n352), .A2(n605), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n386), .A2(n607), .ZN(n643) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n673) );
  AND2_X1 U683 ( .A1(n643), .A2(n673), .ZN(n616) );
  AND2_X1 U684 ( .A1(n618), .A2(n616), .ZN(n734) );
  NAND2_X1 U685 ( .A1(KEYINPUT2), .A2(KEYINPUT66), .ZN(n611) );
  INV_X1 U686 ( .A(KEYINPUT2), .ZN(n612) );
  NOR2_X1 U687 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U688 ( .A1(n614), .A2(KEYINPUT66), .ZN(n615) );
  AND2_X1 U689 ( .A1(n616), .A2(KEYINPUT2), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U691 ( .A(KEYINPUT86), .B(KEYINPUT55), .Z(n621) );
  XOR2_X1 U692 ( .A(n621), .B(KEYINPUT54), .Z(n622) );
  XNOR2_X1 U693 ( .A(n623), .B(n622), .ZN(n624) );
  XNOR2_X1 U694 ( .A(n625), .B(n624), .ZN(n626) );
  NOR2_X1 U695 ( .A1(n626), .A2(n714), .ZN(n628) );
  XNOR2_X1 U696 ( .A(KEYINPUT92), .B(KEYINPUT56), .ZN(n627) );
  XNOR2_X1 U697 ( .A(n628), .B(n627), .ZN(G51) );
  XOR2_X1 U698 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n629) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(n631) );
  XNOR2_X1 U700 ( .A(n632), .B(n631), .ZN(n633) );
  NOR2_X1 U701 ( .A1(n633), .A2(n714), .ZN(n634) );
  XNOR2_X1 U702 ( .A(n634), .B(KEYINPUT122), .ZN(G54) );
  XOR2_X1 U703 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n635) );
  XNOR2_X1 U704 ( .A(n637), .B(n387), .ZN(n638) );
  NOR2_X1 U705 ( .A1(n638), .A2(n714), .ZN(n641) );
  XNOR2_X1 U706 ( .A(KEYINPUT68), .B(KEYINPUT124), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n639), .B(KEYINPUT60), .ZN(n640) );
  XNOR2_X1 U708 ( .A(n641), .B(n640), .ZN(G60) );
  XNOR2_X1 U709 ( .A(n642), .B(G143), .ZN(G45) );
  XNOR2_X1 U710 ( .A(n643), .B(G140), .ZN(G42) );
  XNOR2_X1 U711 ( .A(n644), .B(G110), .ZN(G12) );
  XOR2_X1 U712 ( .A(n645), .B(KEYINPUT62), .Z(n646) );
  XNOR2_X1 U713 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U714 ( .A(KEYINPUT97), .B(KEYINPUT63), .ZN(n649) );
  XOR2_X1 U715 ( .A(n649), .B(KEYINPUT95), .Z(n650) );
  XNOR2_X1 U716 ( .A(n651), .B(n650), .ZN(G57) );
  INV_X1 U717 ( .A(n652), .ZN(n653) );
  XOR2_X1 U718 ( .A(G101), .B(n653), .Z(G3) );
  BUF_X1 U719 ( .A(n654), .Z(n665) );
  NAND2_X1 U720 ( .A1(n665), .A2(n656), .ZN(n655) );
  XNOR2_X1 U721 ( .A(n655), .B(G104), .ZN(G6) );
  XOR2_X1 U722 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n658) );
  NAND2_X1 U723 ( .A1(n656), .A2(n667), .ZN(n657) );
  XNOR2_X1 U724 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U725 ( .A(G107), .B(n659), .ZN(G9) );
  XOR2_X1 U726 ( .A(G128), .B(KEYINPUT29), .Z(n662) );
  INV_X1 U727 ( .A(n660), .ZN(n663) );
  NAND2_X1 U728 ( .A1(n663), .A2(n667), .ZN(n661) );
  XNOR2_X1 U729 ( .A(n662), .B(n661), .ZN(G30) );
  NAND2_X1 U730 ( .A1(n663), .A2(n665), .ZN(n664) );
  XNOR2_X1 U731 ( .A(n664), .B(G146), .ZN(G48) );
  NAND2_X1 U732 ( .A1(n665), .A2(n668), .ZN(n666) );
  XNOR2_X1 U733 ( .A(n666), .B(G113), .ZN(G15) );
  NAND2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U735 ( .A(n669), .B(G116), .ZN(G18) );
  XNOR2_X1 U736 ( .A(n670), .B(KEYINPUT37), .ZN(n671) );
  XNOR2_X1 U737 ( .A(n671), .B(KEYINPUT120), .ZN(n672) );
  XNOR2_X1 U738 ( .A(G125), .B(n672), .ZN(G27) );
  XNOR2_X1 U739 ( .A(G134), .B(n673), .ZN(G36) );
  NOR2_X1 U740 ( .A1(n698), .A2(n688), .ZN(n674) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U742 ( .A(n677), .B(KEYINPUT49), .ZN(n683) );
  NOR2_X1 U743 ( .A1(n678), .A2(n499), .ZN(n679) );
  XOR2_X1 U744 ( .A(KEYINPUT50), .B(n679), .Z(n680) );
  NAND2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U746 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U747 ( .A1(n354), .A2(n684), .ZN(n685) );
  XNOR2_X1 U748 ( .A(n685), .B(KEYINPUT51), .ZN(n686) );
  XNOR2_X1 U749 ( .A(KEYINPUT121), .B(n686), .ZN(n687) );
  NOR2_X1 U750 ( .A1(n688), .A2(n687), .ZN(n700) );
  NOR2_X1 U751 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U752 ( .A1(n692), .A2(n691), .ZN(n696) );
  NOR2_X1 U753 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U754 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U755 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U756 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U757 ( .A(n701), .B(KEYINPUT52), .ZN(n702) );
  NOR2_X1 U758 ( .A1(n703), .A2(n702), .ZN(n705) );
  AND2_X1 U759 ( .A1(n620), .A2(n734), .ZN(n704) );
  XOR2_X1 U760 ( .A(KEYINPUT53), .B(n706), .Z(G75) );
  XNOR2_X1 U761 ( .A(n707), .B(KEYINPUT125), .ZN(n708) );
  XNOR2_X1 U762 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U763 ( .A1(n714), .A2(n710), .ZN(G63) );
  XNOR2_X1 U764 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(G66) );
  XNOR2_X1 U766 ( .A(G101), .B(n715), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n717), .B(n716), .ZN(n719) );
  NOR2_X1 U768 ( .A1(n719), .A2(n718), .ZN(n726) );
  NAND2_X1 U769 ( .A1(n620), .A2(n736), .ZN(n723) );
  NAND2_X1 U770 ( .A1(G953), .A2(G224), .ZN(n720) );
  XNOR2_X1 U771 ( .A(KEYINPUT61), .B(n720), .ZN(n721) );
  NAND2_X1 U772 ( .A1(n721), .A2(G898), .ZN(n722) );
  NAND2_X1 U773 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U774 ( .A(n724), .B(KEYINPUT126), .ZN(n725) );
  XNOR2_X1 U775 ( .A(n726), .B(n725), .ZN(G69) );
  XNOR2_X1 U776 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U777 ( .A(n730), .B(n729), .ZN(n735) );
  XNOR2_X1 U778 ( .A(n735), .B(KEYINPUT127), .ZN(n731) );
  XNOR2_X1 U779 ( .A(G227), .B(n731), .ZN(n732) );
  NAND2_X1 U780 ( .A1(G900), .A2(n732), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n733), .A2(G953), .ZN(n739) );
  XNOR2_X1 U782 ( .A(n735), .B(n734), .ZN(n737) );
  NAND2_X1 U783 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U784 ( .A1(n739), .A2(n738), .ZN(G72) );
  XNOR2_X1 U785 ( .A(G122), .B(n534), .ZN(G24) );
  XOR2_X1 U786 ( .A(n740), .B(G119), .Z(G21) );
  XNOR2_X1 U787 ( .A(G137), .B(n741), .ZN(G39) );
  XNOR2_X1 U788 ( .A(G131), .B(n742), .ZN(G33) );
endmodule

