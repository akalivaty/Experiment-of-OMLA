//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  INV_X1    g000(.A(G131), .ZN(new_n187));
  INV_X1    g001(.A(G137), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G134), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G137), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n187), .B1(new_n189), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G128), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n199), .B1(G143), .B2(new_n193), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n197), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(new_n199), .A3(G128), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n192), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n205), .B1(new_n190), .B2(G137), .ZN(new_n206));
  AOI21_X1  g020(.A(G131), .B1(new_n190), .B2(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n188), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n211));
  NAND4_X1  g025(.A1(new_n206), .A2(new_n207), .A3(new_n211), .A4(new_n208), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n204), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G116), .B(G119), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT2), .B(G113), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XOR2_X1   g032(.A(KEYINPUT2), .B(G113), .Z(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n215), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n206), .A2(new_n208), .A3(new_n191), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n210), .A2(new_n212), .B1(G131), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  OR2_X1    g039(.A1(KEYINPUT0), .A2(G128), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n197), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n202), .A2(KEYINPUT0), .A3(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n214), .B(new_n222), .C1(new_n224), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(G131), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n213), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n227), .A2(new_n228), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(KEYINPUT65), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n224), .B2(new_n229), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n204), .A2(new_n213), .A3(KEYINPUT67), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT67), .B1(new_n204), .B2(new_n213), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT30), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n232), .A2(new_n233), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n214), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT30), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n221), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n230), .B1(new_n241), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n247));
  XOR2_X1   g061(.A(KEYINPUT26), .B(G101), .Z(new_n248));
  NOR2_X1   g062(.A1(G237), .A2(G953), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G210), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n248), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n246), .A2(new_n247), .A3(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n247), .B1(new_n246), .B2(new_n253), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n230), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n242), .A2(KEYINPUT28), .A3(new_n222), .A4(new_n214), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT65), .B1(new_n232), .B2(new_n233), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n224), .A2(new_n235), .A3(new_n229), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n239), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n204), .A2(new_n213), .A3(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n221), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n253), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n259), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT29), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n254), .A2(new_n255), .A3(new_n270), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n257), .A2(KEYINPUT70), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n243), .A2(new_n221), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n256), .B1(new_n273), .B2(new_n230), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n257), .A2(KEYINPUT70), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n272), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(KEYINPUT29), .A3(new_n267), .ZN(new_n277));
  INV_X1    g091(.A(G902), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(G472), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT71), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n267), .B1(new_n259), .B2(new_n266), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n267), .B(new_n230), .C1(new_n241), .C2(new_n245), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT31), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n284), .A2(new_n285), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n283), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  NOR2_X1   g103(.A1(G472), .A2(G902), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n244), .B1(new_n262), .B2(new_n265), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n242), .A2(new_n214), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n222), .B1(new_n293), .B2(KEYINPUT30), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n295), .A2(KEYINPUT31), .A3(new_n267), .A4(new_n230), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n284), .A2(new_n285), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n282), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n290), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT32), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n291), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT71), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n302), .B(G472), .C1(new_n271), .C2(new_n279), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n281), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G128), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT88), .B1(new_n305), .B2(G143), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT88), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(new_n195), .A3(G128), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT89), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n310), .B1(new_n198), .B2(G143), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n305), .A2(KEYINPUT66), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G128), .ZN(new_n314));
  AND4_X1   g128(.A1(new_n310), .A2(new_n312), .A3(new_n314), .A4(G143), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n309), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT90), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n312), .A2(new_n314), .A3(G143), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT89), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n198), .A2(new_n310), .A3(G143), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT90), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(new_n309), .ZN(new_n323));
  AOI21_X1  g137(.A(G134), .B1(new_n317), .B2(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n311), .A2(new_n315), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT13), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n309), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT13), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(G134), .B1(new_n325), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G116), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G122), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n331), .A2(G122), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OR2_X1    g149(.A1(KEYINPUT76), .A2(G107), .ZN(new_n336));
  NAND2_X1  g150(.A1(KEYINPUT76), .A2(G107), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n335), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n330), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT91), .B1(new_n324), .B2(new_n340), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n321), .A2(new_n322), .A3(new_n309), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n322), .B1(new_n321), .B2(new_n309), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n190), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT91), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n333), .A2(new_n334), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(new_n338), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n321), .A2(new_n327), .A3(new_n328), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n348), .B2(G134), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n344), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n341), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g165(.A(KEYINPUT9), .B(G234), .Z(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT75), .ZN(new_n353));
  INV_X1    g167(.A(G953), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(G217), .A3(new_n354), .ZN(new_n355));
  XOR2_X1   g169(.A(new_n355), .B(KEYINPUT93), .Z(new_n356));
  NOR2_X1   g170(.A1(new_n335), .A2(new_n338), .ZN(new_n357));
  INV_X1    g171(.A(G107), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT92), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT14), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n359), .B1(new_n333), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n332), .B1(new_n334), .B2(KEYINPUT14), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n358), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n362), .A2(KEYINPUT92), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n357), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n342), .A2(new_n343), .A3(new_n190), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n365), .B1(new_n366), .B2(new_n324), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n351), .A2(new_n356), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n356), .B1(new_n351), .B2(new_n367), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n278), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G478), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT94), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(KEYINPUT15), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(KEYINPUT15), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n376), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n278), .B(new_n378), .C1(new_n368), .C2(new_n369), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G475), .ZN(new_n382));
  XNOR2_X1  g196(.A(G125), .B(G140), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n193), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT74), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT74), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n386), .A3(new_n193), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G140), .ZN(new_n389));
  INV_X1    g203(.A(G125), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n389), .B1(new_n390), .B2(KEYINPUT73), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT73), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(G125), .A3(G140), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT84), .B1(new_n394), .B2(new_n193), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n193), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n388), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G237), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n354), .A3(G214), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n195), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n249), .A2(G143), .A3(G214), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT18), .A2(G131), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n399), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n402), .A2(new_n404), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G131), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n402), .A2(new_n187), .A3(new_n404), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(KEYINPUT17), .A3(G131), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT16), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n390), .B2(G140), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n193), .B(new_n416), .C1(new_n394), .C2(new_n415), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n416), .B1(new_n394), .B2(new_n415), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G146), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n413), .A2(new_n414), .A3(new_n417), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n408), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G113), .B(G122), .ZN(new_n422));
  INV_X1    g236(.A(G104), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n408), .A2(new_n424), .A3(new_n420), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n382), .B1(new_n428), .B2(new_n278), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT86), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n410), .A2(new_n412), .B1(new_n418), .B2(G146), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT19), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n383), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n434), .B(new_n193), .C1(new_n433), .C2(new_n394), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n399), .A2(new_n407), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n431), .B1(new_n436), .B2(new_n424), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n385), .A2(new_n387), .B1(new_n396), .B2(new_n397), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n405), .A2(new_n406), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n405), .A2(new_n406), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n438), .A2(new_n395), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n410), .A2(new_n412), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n442), .A2(new_n419), .A3(new_n435), .ZN(new_n443));
  OAI211_X1 g257(.A(KEYINPUT86), .B(new_n425), .C1(new_n441), .C2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n437), .A2(new_n427), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n382), .A2(new_n278), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT87), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n446), .B1(new_n445), .B2(new_n448), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n430), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G952), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(G953), .ZN(new_n454));
  NAND2_X1  g268(.A1(G234), .A2(G237), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT95), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(G902), .ZN(new_n458));
  INV_X1    g272(.A(G898), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n354), .B1(KEYINPUT21), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(KEYINPUT21), .B2(new_n459), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n457), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n452), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n381), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G221), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n466), .B1(new_n353), .B2(new_n278), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT77), .B(G469), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n197), .B1(new_n200), .B2(new_n305), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n203), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n423), .A2(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n336), .A3(new_n337), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT3), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n358), .B1(new_n473), .B2(G104), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(G104), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G101), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n472), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(G104), .B2(G107), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n479), .B1(new_n338), .B2(G104), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n470), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT10), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT4), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n471), .A2(new_n336), .A3(new_n337), .ZN(new_n485));
  AOI21_X1  g299(.A(G107), .B1(new_n423), .B2(KEYINPUT3), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(new_n471), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n484), .B(G101), .C1(new_n485), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n478), .A2(KEYINPUT4), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n477), .B1(new_n472), .B2(new_n476), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n233), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n201), .A2(new_n203), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(KEYINPUT10), .A3(new_n478), .A4(new_n480), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n483), .A2(new_n491), .A3(new_n224), .A4(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G110), .B(G140), .ZN(new_n495));
  INV_X1    g309(.A(G227), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(G953), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n495), .B(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n478), .A2(new_n480), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n481), .B1(new_n501), .B2(new_n492), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n502), .A2(KEYINPUT12), .A3(new_n232), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT12), .B1(new_n502), .B2(new_n232), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n494), .B(new_n499), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n483), .A2(new_n491), .A3(new_n493), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n232), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n499), .B1(new_n507), .B2(new_n494), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT78), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI211_X1 g324(.A(KEYINPUT78), .B(new_n499), .C1(new_n507), .C2(new_n494), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n278), .B(new_n468), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n494), .B1(new_n503), .B2(new_n504), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n494), .A2(new_n499), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n513), .A2(new_n498), .B1(new_n514), .B2(new_n507), .ZN(new_n515));
  OAI21_X1  g329(.A(G469), .B1(new_n515), .B2(G902), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n467), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G214), .B1(G237), .B2(G902), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n519));
  INV_X1    g333(.A(G113), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n331), .A2(G119), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT79), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT79), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT5), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n215), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n523), .A2(new_n529), .B1(new_n215), .B2(new_n219), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n501), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n221), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(G110), .B(G122), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n519), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT80), .ZN(new_n537));
  OAI21_X1  g351(.A(G101), .B1(new_n485), .B2(new_n487), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT4), .A3(new_n478), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n490), .A2(new_n484), .B1(new_n218), .B2(new_n220), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n539), .A2(new_n540), .B1(new_n501), .B2(new_n530), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n541), .B2(new_n534), .ZN(new_n542));
  AND4_X1   g356(.A1(new_n537), .A2(new_n531), .A3(new_n532), .A4(new_n534), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n536), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n541), .A2(KEYINPUT6), .A3(new_n534), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n229), .A2(G125), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n201), .A2(new_n390), .A3(new_n203), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n354), .A2(G224), .ZN(new_n550));
  XOR2_X1   g364(.A(new_n550), .B(KEYINPUT81), .Z(new_n551));
  XNOR2_X1  g365(.A(new_n549), .B(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n544), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT7), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n547), .A2(new_n555), .A3(new_n548), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n523), .B1(new_n524), .B2(new_n216), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n501), .A2(new_n220), .A3(new_n560), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n501), .A2(new_n530), .A3(KEYINPUT83), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT83), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n523), .A2(new_n529), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n220), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n563), .B1(new_n565), .B2(new_n500), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n561), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n534), .B(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n559), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT80), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n541), .A2(new_n537), .A3(new_n534), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(G902), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n553), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(G210), .B1(G237), .B2(G902), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n553), .A2(new_n575), .A3(new_n577), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n517), .A2(new_n518), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n465), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G217), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(G234), .B2(new_n278), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT25), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT22), .B(G137), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n354), .A2(G221), .A3(G234), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n312), .A2(new_n314), .A3(G119), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT72), .ZN(new_n593));
  INV_X1    g407(.A(G119), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G128), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n593), .B1(new_n592), .B2(new_n595), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT24), .B(G110), .Z(new_n598));
  NOR3_X1   g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT23), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n594), .B2(G128), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n595), .B(new_n601), .C1(new_n592), .C2(new_n600), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(G110), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n419), .B(new_n388), .C1(new_n599), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n419), .A2(new_n417), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n598), .B1(new_n596), .B2(new_n597), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n602), .A2(G110), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n591), .B1(new_n604), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n604), .A2(new_n608), .A3(new_n591), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n587), .B1(new_n612), .B2(G902), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n604), .A2(new_n608), .A3(new_n591), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n609), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(KEYINPUT25), .A3(new_n278), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n586), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n585), .A2(G902), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n304), .A2(new_n583), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G101), .ZN(G3));
  OAI21_X1  g436(.A(G472), .B1(new_n298), .B2(G902), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n298), .A2(new_n299), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT96), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT96), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n626), .A2(new_n620), .A3(new_n517), .A4(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n579), .A2(new_n630), .A3(new_n580), .ZN(new_n631));
  INV_X1    g445(.A(new_n518), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n577), .B1(new_n553), .B2(new_n575), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(KEYINPUT97), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n445), .A2(new_n448), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT20), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n429), .B1(new_n637), .B2(new_n449), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT33), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(new_n368), .B2(new_n369), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n324), .A2(new_n340), .A3(KEYINPUT91), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n345), .B1(new_n344), .B2(new_n349), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n367), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n356), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n351), .A2(new_n356), .A3(new_n367), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n645), .A2(KEYINPUT33), .A3(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n371), .A2(G902), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n640), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n370), .A2(new_n371), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n638), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n462), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n629), .A2(new_n635), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(KEYINPUT34), .B(G104), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  NAND4_X1  g469(.A1(new_n464), .A2(new_n380), .A3(new_n631), .A4(new_n634), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n629), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT35), .B(G107), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  NOR3_X1   g473(.A1(new_n612), .A2(new_n587), .A3(G902), .ZN(new_n660));
  AOI21_X1  g474(.A(KEYINPUT25), .B1(new_n615), .B2(new_n278), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n585), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n604), .A2(new_n608), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n590), .A2(KEYINPUT36), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n618), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n381), .A2(new_n464), .A3(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n582), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n626), .A3(new_n628), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT37), .B(G110), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G12));
  NAND4_X1  g486(.A1(new_n517), .A2(new_n631), .A3(new_n667), .A4(new_n634), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n354), .A2(G900), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(G902), .A3(new_n455), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT98), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n457), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT99), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n380), .A2(new_n638), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n673), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n304), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  INV_X1    g497(.A(new_n666), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n617), .A2(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n380), .A2(new_n685), .A3(new_n518), .A4(new_n452), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT38), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n581), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n678), .B(KEYINPUT39), .Z(new_n689));
  NAND2_X1  g503(.A1(new_n517), .A2(new_n689), .ZN(new_n690));
  AOI211_X1 g504(.A(new_n686), .B(new_n688), .C1(KEYINPUT40), .C2(new_n690), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n691), .B1(KEYINPUT40), .B2(new_n690), .ZN(new_n692));
  INV_X1    g506(.A(G472), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n273), .A2(new_n230), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n284), .B1(new_n267), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n693), .B1(new_n695), .B2(new_n278), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT100), .B1(new_n301), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT100), .ZN(new_n699));
  AOI211_X1 g513(.A(new_n699), .B(new_n696), .C1(new_n291), .C2(new_n300), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n692), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT101), .B(G143), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G45));
  NAND2_X1  g518(.A1(new_n649), .A2(new_n650), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n452), .A3(new_n679), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n706), .A2(new_n673), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n304), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT102), .B(G146), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G48));
  NOR2_X1   g524(.A1(new_n510), .A2(new_n511), .ZN(new_n711));
  OAI21_X1  g525(.A(G469), .B1(new_n711), .B2(G902), .ZN(new_n712));
  INV_X1    g526(.A(new_n467), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n620), .A2(new_n712), .A3(new_n713), .A4(new_n512), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n652), .A2(new_n635), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n304), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT41), .B(G113), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NOR2_X1   g532(.A1(new_n656), .A2(new_n714), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n304), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NAND3_X1  g535(.A1(new_n712), .A2(new_n713), .A3(new_n512), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n668), .A2(new_n635), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n304), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  OAI211_X1 g539(.A(new_n272), .B(new_n253), .C1(new_n274), .C2(new_n275), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n726), .B1(new_n286), .B2(new_n287), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n290), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n623), .A2(new_n728), .A3(new_n620), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT103), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT103), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n623), .A2(new_n728), .A3(new_n731), .A4(new_n620), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n631), .A2(new_n634), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n380), .A3(new_n452), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n722), .A2(new_n463), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n733), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  NAND3_X1  g553(.A1(new_n623), .A2(new_n728), .A3(new_n667), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n740), .A2(new_n706), .ZN(new_n741));
  INV_X1    g555(.A(new_n722), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n734), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  NAND2_X1  g558(.A1(new_n304), .A2(new_n620), .ZN(new_n745));
  INV_X1    g559(.A(new_n517), .ZN(new_n746));
  INV_X1    g560(.A(new_n581), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n518), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n706), .A2(KEYINPUT42), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT104), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n304), .A2(new_n752), .A3(new_n620), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n752), .B1(new_n304), .B2(new_n620), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n748), .A2(new_n746), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n755), .A2(new_n651), .A3(new_n679), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n751), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(KEYINPUT105), .B(G131), .Z(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G33));
  INV_X1    g575(.A(new_n680), .ZN(new_n762));
  AND4_X1   g576(.A1(new_n304), .A2(new_n620), .A3(new_n762), .A4(new_n755), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n190), .ZN(G36));
  INV_X1    g578(.A(G469), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n278), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n515), .A2(KEYINPUT45), .ZN(new_n768));
  OAI21_X1  g582(.A(G469), .B1(new_n515), .B2(KEYINPUT45), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT46), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(KEYINPUT46), .B(new_n767), .C1(new_n768), .C2(new_n769), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n512), .A3(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(new_n713), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n689), .ZN(new_n776));
  AOI211_X1 g590(.A(KEYINPUT43), .B(new_n452), .C1(new_n649), .C2(new_n650), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n638), .B(KEYINPUT106), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n705), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n777), .B1(new_n779), .B2(KEYINPUT43), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n626), .A2(new_n628), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n667), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n748), .B(new_n776), .C1(new_n782), .C2(new_n783), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G137), .ZN(G39));
  NAND2_X1  g601(.A1(new_n775), .A2(KEYINPUT47), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n774), .A2(new_n713), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NOR4_X1   g606(.A1(new_n304), .A2(new_n620), .A3(new_n706), .A4(new_n748), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT107), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G140), .ZN(G42));
  NAND3_X1  g610(.A1(new_n620), .A2(new_n713), .A3(new_n518), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT108), .ZN(new_n798));
  INV_X1    g612(.A(new_n688), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n798), .A2(new_n799), .A3(new_n779), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n712), .A2(new_n512), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT49), .Z(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n701), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n380), .A2(new_n685), .A3(new_n452), .A4(new_n679), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n805), .A2(new_n746), .A3(new_n635), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n698), .B2(new_n700), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n304), .B1(new_n707), .B2(new_n681), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n808), .A3(new_n743), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n807), .A2(new_n808), .A3(KEYINPUT52), .A4(new_n743), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n304), .B1(new_n715), .B2(new_n719), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(new_n738), .A3(new_n724), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT109), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n814), .A2(new_n738), .A3(new_n724), .A4(KEYINPUT109), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n745), .A2(KEYINPUT104), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n304), .A2(new_n752), .A3(new_n620), .ZN(new_n821));
  INV_X1    g635(.A(new_n756), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT42), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT111), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n380), .A2(new_n825), .ZN(new_n826));
  AOI211_X1 g640(.A(new_n632), .B(new_n463), .C1(new_n579), .C2(new_n580), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n377), .A2(new_n379), .A3(KEYINPUT111), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n826), .A2(new_n827), .A3(new_n638), .A4(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n651), .A3(KEYINPUT110), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n827), .A2(new_n651), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT110), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n629), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n670), .A2(new_n621), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n667), .A2(new_n638), .A3(new_n679), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n826), .B2(new_n828), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n304), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(new_n741), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n763), .B1(new_n755), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n824), .A2(new_n837), .A3(new_n751), .A4(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n804), .B1(new_n819), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n670), .A2(new_n621), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n842), .A2(new_n755), .ZN(new_n847));
  INV_X1    g661(.A(new_n629), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n833), .A2(KEYINPUT110), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n849), .B2(new_n831), .ZN(new_n850));
  INV_X1    g664(.A(new_n763), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n846), .A2(new_n847), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n759), .A2(new_n852), .ZN(new_n853));
  AOI211_X1 g667(.A(new_n804), .B(new_n815), .C1(new_n811), .C2(new_n812), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n845), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n817), .A2(new_n818), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n853), .A2(KEYINPUT53), .A3(new_n813), .A4(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n856), .B1(new_n860), .B2(new_n845), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT112), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n733), .ZN(new_n863));
  INV_X1    g677(.A(new_n457), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n780), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(KEYINPUT113), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n780), .A2(new_n867), .A3(new_n864), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n863), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(KEYINPUT114), .A3(new_n734), .A4(new_n742), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n867), .B1(new_n780), .B2(new_n864), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT43), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n778), .B2(new_n705), .ZN(new_n874));
  NOR4_X1   g688(.A1(new_n874), .A2(KEYINPUT113), .A3(new_n777), .A4(new_n457), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n742), .B(new_n733), .C1(new_n872), .C2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n871), .B1(new_n876), .B2(new_n635), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n748), .A2(new_n722), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n872), .B2(new_n875), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n820), .A2(new_n821), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n880), .A2(new_n620), .A3(new_n864), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n884), .A2(new_n698), .A3(new_n700), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n651), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n454), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n881), .A2(new_n882), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT48), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(KEYINPUT115), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n887), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n878), .A2(new_n883), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT116), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n878), .A2(new_n891), .A3(KEYINPUT116), .A4(new_n883), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n799), .A2(new_n518), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n869), .A2(KEYINPUT50), .A3(new_n742), .A4(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT50), .ZN(new_n898));
  INV_X1    g712(.A(new_n896), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n876), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n740), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n902), .B(new_n880), .C1(new_n872), .C2(new_n875), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n885), .A2(new_n638), .A3(new_n649), .A4(new_n650), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n712), .A2(new_n467), .A3(new_n512), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n788), .A2(new_n791), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n748), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n733), .B1(new_n872), .B2(new_n875), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n903), .B(new_n904), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT51), .B1(new_n901), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n910), .B1(new_n900), .B2(new_n897), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT51), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n894), .A2(new_n895), .B1(new_n911), .B2(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n813), .A2(new_n817), .A3(new_n818), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT53), .B1(new_n916), .B2(new_n853), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n819), .A2(new_n844), .A3(new_n804), .ZN(new_n918));
  OAI21_X1  g732(.A(KEYINPUT54), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT112), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n845), .A2(new_n855), .A3(new_n856), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n862), .A2(new_n915), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n453), .A2(new_n354), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n923), .B2(new_n924), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n803), .B1(new_n925), .B2(new_n927), .ZN(G75));
  NOR2_X1   g742(.A1(new_n354), .A2(G952), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n278), .B1(new_n845), .B2(new_n855), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT56), .B1(new_n931), .B2(G210), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n545), .B1(new_n574), .B2(new_n536), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(new_n552), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT55), .Z(new_n935));
  OAI21_X1  g749(.A(new_n930), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n932), .B2(new_n935), .ZN(G51));
  NAND2_X1  g751(.A1(new_n845), .A2(new_n855), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT54), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n939), .A2(KEYINPUT118), .A3(new_n921), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT118), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n938), .A2(new_n941), .A3(KEYINPUT54), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n766), .B(KEYINPUT57), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n711), .B(KEYINPUT119), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n768), .A2(new_n769), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n931), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n929), .B1(new_n946), .B2(new_n948), .ZN(G54));
  NAND3_X1  g763(.A1(new_n931), .A2(KEYINPUT58), .A3(G475), .ZN(new_n950));
  INV_X1    g764(.A(new_n445), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n952), .A2(new_n953), .A3(new_n929), .ZN(G60));
  AND2_X1   g768(.A1(new_n640), .A2(new_n647), .ZN(new_n955));
  NAND2_X1  g769(.A1(G478), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT59), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n940), .A2(new_n942), .A3(new_n958), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n959), .A2(KEYINPUT120), .A3(new_n930), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT120), .B1(new_n959), .B2(new_n930), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n862), .A2(new_n922), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n955), .B1(new_n962), .B2(new_n957), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(G63));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT60), .Z(new_n966));
  AND2_X1   g780(.A1(new_n938), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n665), .B(KEYINPUT121), .Z(new_n968));
  AOI21_X1  g782(.A(new_n929), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n938), .A2(new_n966), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n612), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT122), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n974), .A3(KEYINPUT61), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n969), .B(new_n971), .C1(new_n973), .C2(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n975), .A2(new_n977), .ZN(G66));
  OAI21_X1  g792(.A(new_n461), .B1(G224), .B2(new_n354), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT123), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n859), .A2(new_n837), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n980), .B1(new_n982), .B2(G953), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n933), .B1(new_n459), .B2(G953), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n983), .B(new_n984), .Z(G69));
  NAND2_X1  g799(.A1(new_n808), .A2(new_n743), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n702), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT62), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n826), .A2(new_n638), .A3(new_n828), .ZN(new_n990));
  INV_X1    g804(.A(new_n651), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n690), .B(new_n748), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(new_n304), .A3(new_n620), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n795), .A2(new_n786), .A3(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n354), .B1(new_n989), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n241), .B1(KEYINPUT30), .B2(new_n293), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n434), .B1(new_n433), .B2(new_n394), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT124), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  AOI211_X1 g814(.A(new_n763), .B(new_n986), .C1(new_n784), .C2(new_n785), .ZN(new_n1001));
  INV_X1    g815(.A(new_n759), .ZN(new_n1002));
  OR3_X1    g816(.A1(new_n882), .A2(new_n735), .A3(new_n776), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n1001), .A2(new_n1002), .A3(new_n795), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n674), .B1(new_n1004), .B2(new_n354), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n1000), .B(KEYINPUT125), .C1(new_n1005), .C2(new_n998), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n674), .B1(new_n496), .B2(G953), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1006), .B(new_n1008), .ZN(G72));
  NAND2_X1  g823(.A1(G472), .A2(G902), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT63), .Z(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n917), .A2(new_n918), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n254), .A2(new_n255), .ZN(new_n1014));
  AOI211_X1 g828(.A(new_n1012), .B(new_n1013), .C1(new_n284), .C2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1004), .A2(new_n981), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1016), .A2(new_n1012), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n246), .B(KEYINPUT126), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n253), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n930), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n989), .A2(new_n994), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1011), .B1(new_n1021), .B2(new_n981), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1018), .A2(new_n253), .ZN(new_n1023));
  AOI211_X1 g837(.A(new_n1015), .B(new_n1020), .C1(new_n1022), .C2(new_n1023), .ZN(G57));
endmodule


