

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591;

  XNOR2_X1 U327 ( .A(n298), .B(n332), .ZN(n381) );
  XNOR2_X1 U328 ( .A(n340), .B(n386), .ZN(n410) );
  XNOR2_X1 U329 ( .A(n410), .B(KEYINPUT41), .ZN(n467) );
  NOR2_X1 U330 ( .A1(n571), .A2(n570), .ZN(n573) );
  NOR2_X2 U331 ( .A1(n483), .A2(n462), .ZN(n568) );
  XNOR2_X1 U332 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n418) );
  XNOR2_X1 U333 ( .A(n355), .B(n295), .ZN(n356) );
  XNOR2_X1 U334 ( .A(n394), .B(n345), .ZN(n349) );
  INV_X1 U335 ( .A(KEYINPUT72), .ZN(n343) );
  XNOR2_X1 U336 ( .A(n357), .B(n356), .ZN(n362) );
  XOR2_X1 U337 ( .A(n354), .B(n353), .Z(n295) );
  XOR2_X1 U338 ( .A(n336), .B(n335), .Z(n296) );
  XOR2_X1 U339 ( .A(n401), .B(n400), .Z(n297) );
  XOR2_X1 U340 ( .A(KEYINPUT13), .B(KEYINPUT73), .Z(n298) );
  XNOR2_X1 U341 ( .A(n443), .B(KEYINPUT64), .ZN(n574) );
  XNOR2_X1 U342 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U343 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U344 ( .A(n344), .B(n343), .ZN(n345) );
  INV_X1 U345 ( .A(n574), .ZN(n576) );
  XNOR2_X1 U346 ( .A(n402), .B(n297), .ZN(n403) );
  XNOR2_X1 U347 ( .A(n404), .B(n403), .ZN(n408) );
  XNOR2_X1 U348 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U349 ( .A(n470), .B(n469), .ZN(G1349GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n300) );
  XNOR2_X1 U351 ( .A(G190GAT), .B(KEYINPUT90), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U353 ( .A(n301), .B(KEYINPUT19), .Z(n303) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(G183GAT), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n325) );
  XOR2_X1 U356 ( .A(KEYINPUT88), .B(KEYINPUT0), .Z(n305) );
  XNOR2_X1 U357 ( .A(G113GAT), .B(KEYINPUT87), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n305), .B(n304), .ZN(n434) );
  XOR2_X1 U359 ( .A(G43GAT), .B(G134GAT), .Z(n392) );
  XOR2_X1 U360 ( .A(n434), .B(n392), .Z(n307) );
  NAND2_X1 U361 ( .A1(G227GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U362 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U363 ( .A(G71GAT), .B(KEYINPUT89), .Z(n309) );
  XNOR2_X1 U364 ( .A(G99GAT), .B(KEYINPUT20), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U366 ( .A(n311), .B(n310), .Z(n313) );
  XOR2_X1 U367 ( .A(G15GAT), .B(G127GAT), .Z(n377) );
  XOR2_X1 U368 ( .A(G176GAT), .B(G120GAT), .Z(n339) );
  XNOR2_X1 U369 ( .A(n377), .B(n339), .ZN(n312) );
  XNOR2_X1 U370 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U371 ( .A(n325), .B(n314), .Z(n483) );
  XOR2_X1 U372 ( .A(G36GAT), .B(KEYINPUT80), .Z(n387) );
  XOR2_X1 U373 ( .A(G92GAT), .B(G64GAT), .Z(n335) );
  XNOR2_X1 U374 ( .A(n387), .B(n335), .ZN(n319) );
  XNOR2_X1 U375 ( .A(G8GAT), .B(G211GAT), .ZN(n315) );
  XNOR2_X1 U376 ( .A(n315), .B(KEYINPUT81), .ZN(n375) );
  XOR2_X1 U377 ( .A(n375), .B(G176GAT), .Z(n317) );
  NAND2_X1 U378 ( .A1(G226GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U380 ( .A(n319), .B(n318), .ZN(n327) );
  XOR2_X1 U381 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n321) );
  XNOR2_X1 U382 ( .A(G218GAT), .B(KEYINPUT93), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U384 ( .A(n322), .B(KEYINPUT21), .Z(n324) );
  XNOR2_X1 U385 ( .A(G197GAT), .B(G204GAT), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n324), .B(n323), .ZN(n456) );
  XOR2_X1 U387 ( .A(n325), .B(n456), .Z(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n492) );
  XNOR2_X1 U389 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n407) );
  XOR2_X1 U390 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n329) );
  NAND2_X1 U391 ( .A1(G230GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U392 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U393 ( .A(n330), .B(KEYINPUT33), .Z(n334) );
  XNOR2_X1 U394 ( .A(G106GAT), .B(G78GAT), .ZN(n331) );
  XNOR2_X1 U395 ( .A(n331), .B(G148GAT), .ZN(n455) );
  XNOR2_X1 U396 ( .A(G71GAT), .B(G57GAT), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n455), .B(n381), .ZN(n333) );
  XNOR2_X1 U398 ( .A(n334), .B(n333), .ZN(n336) );
  XNOR2_X1 U399 ( .A(G204GAT), .B(KEYINPUT74), .ZN(n337) );
  XNOR2_X1 U400 ( .A(n296), .B(n337), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U402 ( .A(G99GAT), .B(G85GAT), .ZN(n386) );
  XOR2_X1 U403 ( .A(G29GAT), .B(KEYINPUT69), .Z(n342) );
  XNOR2_X1 U404 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n341) );
  XNOR2_X1 U405 ( .A(n342), .B(n341), .ZN(n394) );
  NAND2_X1 U406 ( .A1(G229GAT), .A2(G233GAT), .ZN(n344) );
  XOR2_X1 U407 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n347) );
  XNOR2_X1 U408 ( .A(G169GAT), .B(G8GAT), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n357) );
  XOR2_X1 U411 ( .A(G50GAT), .B(G43GAT), .Z(n352) );
  XNOR2_X1 U412 ( .A(G1GAT), .B(KEYINPUT70), .ZN(n350) );
  XOR2_X1 U413 ( .A(n350), .B(KEYINPUT71), .Z(n382) );
  XOR2_X1 U414 ( .A(G22GAT), .B(n382), .Z(n351) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n355) );
  XOR2_X1 U416 ( .A(G15GAT), .B(G113GAT), .Z(n354) );
  XNOR2_X1 U417 ( .A(G141GAT), .B(G197GAT), .ZN(n353) );
  XOR2_X1 U418 ( .A(KEYINPUT65), .B(KEYINPUT68), .Z(n359) );
  XNOR2_X1 U419 ( .A(KEYINPUT30), .B(KEYINPUT67), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U421 ( .A(n360), .B(G36GAT), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n577) );
  NAND2_X1 U423 ( .A1(n467), .A2(n577), .ZN(n363) );
  XNOR2_X1 U424 ( .A(n363), .B(KEYINPUT46), .ZN(n384) );
  XOR2_X1 U425 ( .A(KEYINPUT84), .B(KEYINPUT85), .Z(n365) );
  XNOR2_X1 U426 ( .A(G183GAT), .B(G78GAT), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U428 ( .A(KEYINPUT12), .B(KEYINPUT83), .Z(n367) );
  XNOR2_X1 U429 ( .A(KEYINPUT14), .B(KEYINPUT82), .ZN(n366) );
  XNOR2_X1 U430 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U431 ( .A(n369), .B(n368), .Z(n374) );
  XOR2_X1 U432 ( .A(KEYINPUT86), .B(G64GAT), .Z(n371) );
  NAND2_X1 U433 ( .A1(G231GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U435 ( .A(KEYINPUT15), .B(n372), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n376) );
  XOR2_X1 U437 ( .A(n376), .B(n375), .Z(n379) );
  XOR2_X1 U438 ( .A(G22GAT), .B(G155GAT), .Z(n447) );
  XNOR2_X1 U439 ( .A(n377), .B(n447), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n383) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n561) );
  XNOR2_X1 U443 ( .A(KEYINPUT112), .B(n561), .ZN(n570) );
  NAND2_X1 U444 ( .A1(n384), .A2(n570), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n385), .B(KEYINPUT113), .ZN(n405) );
  XNOR2_X1 U446 ( .A(KEYINPUT11), .B(n386), .ZN(n389) );
  XNOR2_X1 U447 ( .A(G218GAT), .B(n387), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U449 ( .A(n390), .B(G92GAT), .Z(n397) );
  AND2_X1 U450 ( .A1(G232GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n395), .B(G190GAT), .ZN(n396) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U453 ( .A(KEYINPUT9), .B(n398), .Z(n404) );
  XNOR2_X1 U454 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n399), .B(G162GAT), .ZN(n450) );
  XNOR2_X1 U456 ( .A(n450), .B(KEYINPUT10), .ZN(n402) );
  XOR2_X1 U457 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n401) );
  XNOR2_X1 U458 ( .A(G106GAT), .B(KEYINPUT79), .ZN(n400) );
  NAND2_X1 U459 ( .A1(n405), .A2(n408), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n416) );
  XNOR2_X1 U461 ( .A(n408), .B(KEYINPUT36), .ZN(n589) );
  NOR2_X1 U462 ( .A1(n561), .A2(n589), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n409), .B(KEYINPUT45), .ZN(n412) );
  INV_X1 U464 ( .A(n577), .ZN(n513) );
  AND2_X1 U465 ( .A1(n410), .A2(n513), .ZN(n411) );
  AND2_X1 U466 ( .A1(n412), .A2(n411), .ZN(n414) );
  INV_X1 U467 ( .A(KEYINPUT115), .ZN(n413) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n415) );
  NOR2_X1 U469 ( .A1(n416), .A2(n415), .ZN(n417) );
  XNOR2_X1 U470 ( .A(n417), .B(KEYINPUT48), .ZN(n537) );
  NOR2_X1 U471 ( .A1(n492), .A2(n537), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n419), .B(n418), .ZN(n442) );
  XOR2_X1 U473 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n421) );
  XNOR2_X1 U474 ( .A(G1GAT), .B(KEYINPUT101), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n427) );
  XOR2_X1 U476 ( .A(KEYINPUT96), .B(KEYINPUT3), .Z(n423) );
  XNOR2_X1 U477 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n453) );
  XOR2_X1 U479 ( .A(n453), .B(KEYINPUT100), .Z(n425) );
  NAND2_X1 U480 ( .A1(G225GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n441) );
  XOR2_X1 U483 ( .A(G155GAT), .B(G148GAT), .Z(n429) );
  XNOR2_X1 U484 ( .A(G127GAT), .B(G120GAT), .ZN(n428) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U486 ( .A(G57GAT), .B(KEYINPUT99), .Z(n431) );
  XNOR2_X1 U487 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U489 ( .A(n433), .B(n432), .Z(n439) );
  XOR2_X1 U490 ( .A(G85GAT), .B(G162GAT), .Z(n436) );
  XNOR2_X1 U491 ( .A(G134GAT), .B(n434), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U493 ( .A(G29GAT), .B(n437), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n480) );
  NAND2_X1 U496 ( .A1(n442), .A2(n480), .ZN(n443) );
  XOR2_X1 U497 ( .A(KEYINPUT24), .B(KEYINPUT97), .Z(n445) );
  XNOR2_X1 U498 ( .A(KEYINPUT22), .B(KEYINPUT92), .ZN(n444) );
  XNOR2_X1 U499 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U500 ( .A(n446), .B(KEYINPUT23), .Z(n449) );
  XNOR2_X1 U501 ( .A(n447), .B(G211GAT), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n460) );
  XOR2_X1 U503 ( .A(n450), .B(KEYINPUT98), .Z(n452) );
  NAND2_X1 U504 ( .A1(G228GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n454) );
  XOR2_X1 U506 ( .A(n454), .B(n453), .Z(n458) );
  XNOR2_X1 U507 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U508 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U509 ( .A(n460), .B(n459), .Z(n479) );
  NOR2_X1 U510 ( .A1(n574), .A2(n479), .ZN(n461) );
  XNOR2_X1 U511 ( .A(n461), .B(KEYINPUT55), .ZN(n462) );
  INV_X1 U512 ( .A(n568), .ZN(n571) );
  NOR2_X1 U513 ( .A1(n571), .A2(n408), .ZN(n466) );
  XNOR2_X1 U514 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n464) );
  INV_X1 U515 ( .A(G190GAT), .ZN(n463) );
  XNOR2_X1 U516 ( .A(n466), .B(n465), .ZN(G1351GAT) );
  BUF_X1 U517 ( .A(n467), .Z(n557) );
  NAND2_X1 U518 ( .A1(n568), .A2(n557), .ZN(n470) );
  XOR2_X1 U519 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n468) );
  XNOR2_X1 U520 ( .A(n468), .B(G176GAT), .ZN(n469) );
  XOR2_X1 U521 ( .A(KEYINPUT103), .B(KEYINPUT34), .Z(n490) );
  NAND2_X1 U522 ( .A1(n410), .A2(n577), .ZN(n471) );
  XOR2_X1 U523 ( .A(KEYINPUT75), .B(n471), .Z(n501) );
  INV_X1 U524 ( .A(n408), .ZN(n563) );
  NOR2_X1 U525 ( .A1(n563), .A2(n561), .ZN(n472) );
  XNOR2_X1 U526 ( .A(n472), .B(KEYINPUT16), .ZN(n488) );
  NOR2_X1 U527 ( .A1(n483), .A2(n492), .ZN(n473) );
  NOR2_X1 U528 ( .A1(n479), .A2(n473), .ZN(n474) );
  XNOR2_X1 U529 ( .A(n474), .B(KEYINPUT25), .ZN(n477) );
  XOR2_X1 U530 ( .A(KEYINPUT27), .B(n492), .Z(n481) );
  NAND2_X1 U531 ( .A1(n479), .A2(n483), .ZN(n475) );
  XOR2_X1 U532 ( .A(n475), .B(KEYINPUT26), .Z(n575) );
  NAND2_X1 U533 ( .A1(n481), .A2(n575), .ZN(n476) );
  NAND2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U535 ( .A1(n480), .A2(n478), .ZN(n487) );
  XNOR2_X1 U536 ( .A(n479), .B(KEYINPUT28), .ZN(n542) );
  INV_X1 U537 ( .A(n480), .ZN(n527) );
  NAND2_X1 U538 ( .A1(n527), .A2(n481), .ZN(n538) );
  NOR2_X1 U539 ( .A1(n542), .A2(n538), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n482), .B(KEYINPUT102), .ZN(n485) );
  INV_X1 U541 ( .A(n483), .ZN(n539) );
  XNOR2_X1 U542 ( .A(n539), .B(KEYINPUT91), .ZN(n484) );
  NAND2_X1 U543 ( .A1(n485), .A2(n484), .ZN(n486) );
  NAND2_X1 U544 ( .A1(n487), .A2(n486), .ZN(n498) );
  NAND2_X1 U545 ( .A1(n488), .A2(n498), .ZN(n515) );
  NOR2_X1 U546 ( .A1(n501), .A2(n515), .ZN(n496) );
  NAND2_X1 U547 ( .A1(n496), .A2(n527), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n491), .ZN(G1324GAT) );
  INV_X1 U550 ( .A(n492), .ZN(n529) );
  NAND2_X1 U551 ( .A1(n496), .A2(n529), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n493), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .Z(n495) );
  NAND2_X1 U554 ( .A1(n496), .A2(n539), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NAND2_X1 U556 ( .A1(n542), .A2(n496), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n497), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT39), .B(KEYINPUT104), .Z(n504) );
  NAND2_X1 U559 ( .A1(n561), .A2(n498), .ZN(n499) );
  NOR2_X1 U560 ( .A1(n499), .A2(n589), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n500), .B(KEYINPUT37), .ZN(n526) );
  NOR2_X1 U562 ( .A1(n526), .A2(n501), .ZN(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT38), .B(n502), .ZN(n511) );
  NAND2_X1 U564 ( .A1(n511), .A2(n527), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G29GAT), .B(n505), .ZN(G1328GAT) );
  XOR2_X1 U567 ( .A(G36GAT), .B(KEYINPUT105), .Z(n507) );
  NAND2_X1 U568 ( .A1(n529), .A2(n511), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(G1329GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n509) );
  NAND2_X1 U571 ( .A1(n511), .A2(n539), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U573 ( .A(G43GAT), .B(n510), .Z(G1330GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n542), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n512), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n518) );
  NAND2_X1 U577 ( .A1(n513), .A2(n557), .ZN(n514) );
  XOR2_X1 U578 ( .A(KEYINPUT107), .B(n514), .Z(n525) );
  NOR2_X1 U579 ( .A1(n515), .A2(n525), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n516), .B(KEYINPUT108), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n527), .A2(n521), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1332GAT) );
  NAND2_X1 U583 ( .A1(n521), .A2(n529), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n539), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n523) );
  NAND2_X1 U588 ( .A1(n521), .A2(n542), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U590 ( .A(G78GAT), .B(n524), .Z(G1335GAT) );
  NOR2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n533), .A2(n527), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NAND2_X1 U594 ( .A1(n533), .A2(n529), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(KEYINPUT110), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G92GAT), .B(n531), .ZN(G1337GAT) );
  NAND2_X1 U597 ( .A1(n539), .A2(n533), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n532), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n535) );
  NAND2_X1 U600 ( .A1(n533), .A2(n542), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  XOR2_X1 U603 ( .A(G113GAT), .B(KEYINPUT117), .Z(n544) );
  NOR2_X1 U604 ( .A1(n537), .A2(n538), .ZN(n554) );
  NAND2_X1 U605 ( .A1(n554), .A2(n539), .ZN(n540) );
  XNOR2_X1 U606 ( .A(KEYINPUT116), .B(n540), .ZN(n541) );
  NOR2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n548), .A2(n577), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U611 ( .A1(n548), .A2(n557), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G120GAT), .B(n547), .ZN(G1341GAT) );
  INV_X1 U614 ( .A(n548), .ZN(n551) );
  NOR2_X1 U615 ( .A1(n570), .A2(n551), .ZN(n549) );
  XOR2_X1 U616 ( .A(KEYINPUT50), .B(n549), .Z(n550) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  NOR2_X1 U618 ( .A1(n408), .A2(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  XOR2_X1 U621 ( .A(G141GAT), .B(KEYINPUT119), .Z(n556) );
  AND2_X1 U622 ( .A1(n575), .A2(n554), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n564), .A2(n577), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(G1344GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n559) );
  NAND2_X1 U626 ( .A1(n564), .A2(n557), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(n560), .ZN(G1345GAT) );
  INV_X1 U629 ( .A(n561), .ZN(n585) );
  NAND2_X1 U630 ( .A1(n564), .A2(n585), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n562), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n566) );
  NAND2_X1 U633 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(G162GAT), .B(n567), .ZN(G1347GAT) );
  NAND2_X1 U636 ( .A1(n568), .A2(n577), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n569), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U638 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1350GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n579) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n588) );
  INV_X1 U642 ( .A(n588), .ZN(n584) );
  NAND2_X1 U643 ( .A1(n584), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n582) );
  OR2_X1 U647 ( .A1(n588), .A2(n410), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U649 ( .A(G204GAT), .B(n583), .Z(G1353GAT) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT126), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

