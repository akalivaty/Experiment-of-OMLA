

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776;

  NAND2_X1 U368 ( .A1(n411), .A2(n409), .ZN(n460) );
  XNOR2_X1 U369 ( .A(n608), .B(n609), .ZN(n356) );
  AND2_X1 U370 ( .A1(n352), .A2(n370), .ZN(n627) );
  XNOR2_X1 U371 ( .A(n577), .B(KEYINPUT77), .ZN(n586) );
  AND2_X1 U372 ( .A1(n618), .A2(n695), .ZN(n605) );
  BUF_X1 U373 ( .A(n617), .Z(n618) );
  NOR2_X1 U374 ( .A1(n698), .A2(n699), .ZN(n695) );
  XNOR2_X1 U375 ( .A(n357), .B(n534), .ZN(n698) );
  XNOR2_X1 U376 ( .A(n347), .B(n545), .ZN(n348) );
  XNOR2_X1 U377 ( .A(G140), .B(n490), .ZN(n763) );
  XNOR2_X1 U378 ( .A(n498), .B(n462), .ZN(n347) );
  XNOR2_X1 U379 ( .A(G125), .B(KEYINPUT10), .ZN(n489) );
  INV_X1 U380 ( .A(G902), .ZN(n538) );
  XNOR2_X2 U381 ( .A(n611), .B(KEYINPUT40), .ZN(n623) );
  INV_X2 U382 ( .A(KEYINPUT69), .ZN(n463) );
  AND2_X1 U383 ( .A1(n446), .A2(n445), .ZN(n441) );
  XNOR2_X2 U384 ( .A(n585), .B(KEYINPUT108), .ZN(n405) );
  AND2_X2 U385 ( .A1(n414), .A2(n412), .ZN(n411) );
  NOR2_X1 U386 ( .A1(n732), .A2(n731), .ZN(n363) );
  NAND2_X1 U387 ( .A1(n443), .A2(n642), .ZN(n442) );
  XNOR2_X1 U388 ( .A(n544), .B(n469), .ZN(n507) );
  INV_X1 U389 ( .A(KEYINPUT2), .ZN(n350) );
  INV_X1 U390 ( .A(KEYINPUT121), .ZN(n362) );
  XNOR2_X1 U391 ( .A(n363), .B(n362), .ZN(n361) );
  NOR2_X1 U392 ( .A1(n442), .A2(n350), .ZN(n349) );
  AND2_X1 U393 ( .A1(n379), .A2(KEYINPUT44), .ZN(n378) );
  XNOR2_X1 U394 ( .A(n624), .B(KEYINPUT46), .ZN(n403) );
  NAND2_X1 U395 ( .A1(n410), .A2(n581), .ZN(n409) );
  XNOR2_X1 U396 ( .A(n353), .B(n452), .ZN(n352) );
  XNOR2_X1 U397 ( .A(n447), .B(KEYINPUT111), .ZN(n715) );
  XNOR2_X1 U398 ( .A(n558), .B(n448), .ZN(n711) );
  NOR2_X1 U399 ( .A1(n745), .A2(G902), .ZN(n357) );
  XNOR2_X1 U400 ( .A(n401), .B(n367), .ZN(n615) );
  XNOR2_X1 U401 ( .A(n529), .B(n528), .ZN(n745) );
  XNOR2_X1 U402 ( .A(n459), .B(n506), .ZN(n526) );
  INV_X1 U403 ( .A(KEYINPUT64), .ZN(n471) );
  XNOR2_X2 U404 ( .A(n762), .B(n477), .ZN(n734) );
  XNOR2_X2 U405 ( .A(n383), .B(n470), .ZN(n762) );
  XNOR2_X2 U406 ( .A(n348), .B(n507), .ZN(n383) );
  NAND2_X1 U407 ( .A1(n351), .A2(n349), .ZN(n649) );
  INV_X1 U408 ( .A(n444), .ZN(n351) );
  NOR2_X1 U409 ( .A1(n444), .A2(n442), .ZN(n765) );
  NAND2_X1 U410 ( .A1(n354), .A2(n606), .ZN(n353) );
  XNOR2_X1 U411 ( .A(n605), .B(n453), .ZN(n354) );
  NAND2_X1 U412 ( .A1(n355), .A2(n441), .ZN(n440) );
  INV_X1 U413 ( .A(n403), .ZN(n355) );
  NAND2_X1 U414 ( .A1(n356), .A2(n610), .ZN(n611) );
  NAND2_X1 U415 ( .A1(n356), .A2(n638), .ZN(n640) );
  XNOR2_X1 U416 ( .A(n359), .B(n358), .ZN(G75) );
  INV_X1 U417 ( .A(KEYINPUT53), .ZN(n358) );
  NAND2_X1 U418 ( .A1(n361), .A2(n360), .ZN(n359) );
  INV_X1 U419 ( .A(G953), .ZN(n360) );
  XNOR2_X2 U420 ( .A(n408), .B(G143), .ZN(n544) );
  NAND2_X1 U421 ( .A1(n366), .A2(n644), .ZN(n437) );
  INV_X1 U422 ( .A(G137), .ZN(n462) );
  NAND2_X1 U423 ( .A1(n711), .A2(n612), .ZN(n447) );
  NOR2_X1 U424 ( .A1(n392), .A2(n690), .ZN(n397) );
  INV_X1 U425 ( .A(G237), .ZN(n537) );
  NAND2_X1 U426 ( .A1(n437), .A2(n436), .ZN(n424) );
  OR2_X1 U427 ( .A1(n660), .A2(n425), .ZN(n421) );
  INV_X1 U428 ( .A(n437), .ZN(n425) );
  NAND2_X1 U429 ( .A1(n436), .A2(n553), .ZN(n435) );
  NAND2_X1 U430 ( .A1(n390), .A2(n389), .ZN(n521) );
  INV_X1 U431 ( .A(KEYINPUT38), .ZN(n448) );
  INV_X1 U432 ( .A(KEYINPUT109), .ZN(n453) );
  INV_X1 U433 ( .A(KEYINPUT78), .ZN(n452) );
  NAND2_X1 U434 ( .A1(n422), .A2(n437), .ZN(n407) );
  INV_X1 U435 ( .A(n615), .ZN(n702) );
  XNOR2_X1 U436 ( .A(n418), .B(n567), .ZN(n406) );
  OR2_X1 U437 ( .A1(n377), .A2(n373), .ZN(n418) );
  XNOR2_X1 U438 ( .A(n486), .B(n485), .ZN(n550) );
  XNOR2_X1 U439 ( .A(G116), .B(KEYINPUT71), .ZN(n485) );
  XNOR2_X1 U440 ( .A(n464), .B(G119), .ZN(n486) );
  XNOR2_X1 U441 ( .A(G113), .B(KEYINPUT3), .ZN(n464) );
  XNOR2_X1 U442 ( .A(n527), .B(n457), .ZN(n456) );
  INV_X1 U443 ( .A(KEYINPUT24), .ZN(n457) );
  XNOR2_X1 U444 ( .A(G128), .B(G137), .ZN(n527) );
  XNOR2_X1 U445 ( .A(G110), .B(G119), .ZN(n455) );
  XNOR2_X1 U446 ( .A(KEYINPUT85), .B(KEYINPUT8), .ZN(n506) );
  XNOR2_X1 U447 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U448 ( .A(KEYINPUT9), .B(G107), .Z(n509) );
  XNOR2_X1 U449 ( .A(n756), .B(KEYINPUT72), .ZN(n551) );
  INV_X1 U450 ( .A(KEYINPUT88), .ZN(n466) );
  XNOR2_X1 U451 ( .A(n533), .B(n532), .ZN(n534) );
  BUF_X1 U452 ( .A(n576), .Z(n696) );
  NAND2_X1 U453 ( .A1(n381), .A2(n384), .ZN(n379) );
  INV_X1 U454 ( .A(KEYINPUT70), .ZN(n400) );
  AND2_X1 U455 ( .A1(n396), .A2(n395), .ZN(n394) );
  INV_X1 U456 ( .A(n561), .ZN(n390) );
  XNOR2_X1 U457 ( .A(KEYINPUT93), .B(KEYINPUT15), .ZN(n514) );
  INV_X1 U458 ( .A(KEYINPUT89), .ZN(n598) );
  XNOR2_X1 U459 ( .A(n592), .B(KEYINPUT106), .ZN(n716) );
  NOR2_X1 U460 ( .A1(G953), .A2(G237), .ZN(n491) );
  NAND2_X1 U461 ( .A1(G234), .A2(G237), .ZN(n518) );
  NAND2_X1 U462 ( .A1(n428), .A2(n426), .ZN(n558) );
  NAND2_X1 U463 ( .A1(n432), .A2(n560), .ZN(n431) );
  NAND2_X1 U464 ( .A1(n421), .A2(n423), .ZN(n420) );
  AND2_X1 U465 ( .A1(n424), .A2(n371), .ZN(n423) );
  INV_X1 U466 ( .A(n434), .ZN(n428) );
  XNOR2_X1 U467 ( .A(n531), .B(KEYINPUT98), .ZN(n533) );
  XNOR2_X1 U468 ( .A(G143), .B(G113), .ZN(n494) );
  XNOR2_X1 U469 ( .A(n468), .B(G146), .ZN(n545) );
  XNOR2_X1 U470 ( .A(G125), .B(KEYINPUT80), .ZN(n541) );
  AND2_X1 U471 ( .A1(n413), .A2(n461), .ZN(n412) );
  INV_X1 U472 ( .A(n625), .ZN(n461) );
  NAND2_X1 U473 ( .A1(n387), .A2(n386), .ZN(n629) );
  NAND2_X1 U474 ( .A1(n427), .A2(n428), .ZN(n386) );
  NOR2_X1 U475 ( .A1(n430), .A2(n429), .ZN(n387) );
  NOR2_X1 U476 ( .A1(n407), .A2(n433), .ZN(n427) );
  NAND2_X1 U477 ( .A1(n652), .A2(n538), .ZN(n401) );
  XNOR2_X1 U478 ( .A(n475), .B(n474), .ZN(n756) );
  XNOR2_X1 U479 ( .A(G101), .B(G110), .ZN(n474) );
  XNOR2_X1 U480 ( .A(n550), .B(n549), .ZN(n757) );
  XNOR2_X1 U481 ( .A(n458), .B(n454), .ZN(n528) );
  XNOR2_X1 U482 ( .A(n456), .B(n455), .ZN(n454) );
  XNOR2_X1 U483 ( .A(n510), .B(G116), .ZN(n416) );
  NOR2_X1 U484 ( .A1(n694), .A2(n628), .ZN(n621) );
  NAND2_X1 U485 ( .A1(n620), .A2(n402), .ZN(n680) );
  AND2_X1 U486 ( .A1(n619), .A2(n629), .ZN(n402) );
  INV_X1 U487 ( .A(n638), .ZN(n687) );
  INV_X1 U488 ( .A(G101), .ZN(n571) );
  XNOR2_X1 U489 ( .A(n467), .B(n466), .ZN(n465) );
  NOR2_X1 U490 ( .A1(n377), .A2(n581), .ZN(n365) );
  XOR2_X1 U491 ( .A(n555), .B(KEYINPUT94), .Z(n366) );
  XNOR2_X1 U492 ( .A(G472), .B(KEYINPUT75), .ZN(n367) );
  OR2_X1 U493 ( .A1(G902), .A2(n740), .ZN(n368) );
  AND2_X1 U494 ( .A1(n716), .A2(n415), .ZN(n369) );
  XOR2_X1 U495 ( .A(n607), .B(KEYINPUT30), .Z(n370) );
  AND2_X1 U496 ( .A1(n612), .A2(n433), .ZN(n371) );
  INV_X1 U497 ( .A(n366), .ZN(n436) );
  NOR2_X1 U498 ( .A1(n376), .A2(n589), .ZN(n372) );
  NAND2_X1 U499 ( .A1(n714), .A2(n566), .ZN(n373) );
  XNOR2_X1 U500 ( .A(n565), .B(KEYINPUT0), .ZN(n374) );
  INV_X1 U501 ( .A(KEYINPUT90), .ZN(n384) );
  INV_X1 U502 ( .A(KEYINPUT48), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n399), .B(n400), .ZN(n446) );
  NAND2_X1 U504 ( .A1(n397), .A2(n394), .ZN(n399) );
  XNOR2_X1 U505 ( .A(n507), .B(n416), .ZN(n511) );
  XNOR2_X1 U506 ( .A(n623), .B(G131), .ZN(G33) );
  AND2_X1 U507 ( .A1(n406), .A2(n698), .ZN(n584) );
  XNOR2_X1 U508 ( .A(n617), .B(n481), .ZN(n576) );
  AND2_X1 U509 ( .A1(n434), .A2(n371), .ZN(n429) );
  AND2_X1 U510 ( .A1(n651), .A2(n375), .ZN(n662) );
  AND2_X1 U511 ( .A1(n438), .A2(G210), .ZN(n375) );
  BUF_X1 U512 ( .A(n377), .Z(n376) );
  XNOR2_X1 U513 ( .A(n385), .B(n374), .ZN(n377) );
  BUF_X1 U514 ( .A(n733), .Z(n743) );
  NAND2_X1 U515 ( .A1(n576), .A2(n695), .ZN(n577) );
  NAND2_X1 U516 ( .A1(n376), .A2(n581), .ZN(n413) );
  NOR2_X1 U517 ( .A1(n706), .A2(n376), .ZN(n588) );
  NAND2_X1 U518 ( .A1(n378), .A2(n380), .ZN(n449) );
  NAND2_X1 U519 ( .A1(n380), .A2(n379), .ZN(n419) );
  NAND2_X1 U520 ( .A1(n382), .A2(n405), .ZN(n380) );
  NAND2_X1 U521 ( .A1(n405), .A2(n388), .ZN(n381) );
  AND2_X1 U522 ( .A1(n388), .A2(KEYINPUT90), .ZN(n382) );
  XNOR2_X1 U523 ( .A(n383), .B(n488), .ZN(n652) );
  NAND2_X1 U524 ( .A1(n629), .A2(n564), .ZN(n385) );
  XNOR2_X1 U525 ( .A(n388), .B(G119), .ZN(G21) );
  XNOR2_X2 U526 ( .A(n575), .B(n574), .ZN(n388) );
  NAND2_X1 U527 ( .A1(n391), .A2(G224), .ZN(n546) );
  NAND2_X1 U528 ( .A1(n391), .A2(G234), .ZN(n459) );
  NAND2_X1 U529 ( .A1(n391), .A2(G227), .ZN(n472) );
  OR2_X1 U530 ( .A1(n391), .A2(G952), .ZN(n663) );
  INV_X1 U531 ( .A(n391), .ZN(n389) );
  NAND2_X1 U532 ( .A1(n766), .A2(n391), .ZN(n772) );
  XNOR2_X2 U533 ( .A(n471), .B(G953), .ZN(n391) );
  NOR2_X1 U534 ( .A1(n631), .A2(n393), .ZN(n392) );
  NAND2_X1 U535 ( .A1(n398), .A2(n632), .ZN(n393) );
  INV_X1 U536 ( .A(n679), .ZN(n398) );
  NAND2_X1 U537 ( .A1(n679), .A2(KEYINPUT76), .ZN(n395) );
  NAND2_X1 U538 ( .A1(n631), .A2(KEYINPUT76), .ZN(n396) );
  INV_X1 U539 ( .A(n680), .ZN(n415) );
  NAND2_X1 U540 ( .A1(n620), .A2(n619), .ZN(n628) );
  NAND2_X1 U541 ( .A1(n403), .A2(KEYINPUT48), .ZN(n439) );
  NAND2_X1 U542 ( .A1(n627), .A2(n711), .ZN(n608) );
  XNOR2_X2 U543 ( .A(n404), .B(n757), .ZN(n660) );
  XNOR2_X1 U544 ( .A(n552), .B(n551), .ZN(n404) );
  XNOR2_X1 U545 ( .A(n405), .B(G110), .ZN(G12) );
  NAND2_X1 U546 ( .A1(n406), .A2(n568), .ZN(n467) );
  INV_X1 U547 ( .A(n407), .ZN(n426) );
  XNOR2_X2 U548 ( .A(G128), .B(KEYINPUT83), .ZN(n408) );
  INV_X1 U549 ( .A(n710), .ZN(n410) );
  NAND2_X1 U550 ( .A1(n710), .A2(n365), .ZN(n414) );
  XNOR2_X2 U551 ( .A(n579), .B(KEYINPUT33), .ZN(n710) );
  AND2_X1 U552 ( .A1(n417), .A2(n449), .ZN(n601) );
  NAND2_X1 U553 ( .A1(n450), .A2(n419), .ZN(n417) );
  XNOR2_X1 U554 ( .A(n602), .B(KEYINPUT45), .ZN(n647) );
  NAND2_X1 U555 ( .A1(n420), .A2(n431), .ZN(n430) );
  NAND2_X1 U556 ( .A1(n660), .A2(n366), .ZN(n422) );
  INV_X1 U557 ( .A(n612), .ZN(n432) );
  INV_X1 U558 ( .A(n560), .ZN(n433) );
  NOR2_X1 U559 ( .A1(n660), .A2(n435), .ZN(n434) );
  AND2_X1 U560 ( .A1(n438), .A2(n693), .ZN(n732) );
  AND2_X2 U561 ( .A1(n651), .A2(n438), .ZN(n733) );
  NAND2_X1 U562 ( .A1(n650), .A2(n648), .ZN(n438) );
  NAND2_X1 U563 ( .A1(n440), .A2(n439), .ZN(n444) );
  OR2_X1 U564 ( .A1(n446), .A2(n445), .ZN(n443) );
  INV_X1 U565 ( .A(n558), .ZN(n633) );
  XNOR2_X1 U566 ( .A(n451), .B(KEYINPUT68), .ZN(n450) );
  NOR2_X2 U567 ( .A1(n773), .A2(KEYINPUT44), .ZN(n451) );
  NOR2_X2 U568 ( .A1(n664), .A2(n747), .ZN(n665) );
  NAND2_X1 U569 ( .A1(n526), .A2(G221), .ZN(n458) );
  XNOR2_X2 U570 ( .A(n460), .B(KEYINPUT35), .ZN(n773) );
  XNOR2_X2 U571 ( .A(n463), .B(G131), .ZN(n498) );
  NAND2_X1 U572 ( .A1(n465), .A2(n569), .ZN(n570) );
  BUF_X1 U573 ( .A(n762), .Z(n764) );
  INV_X1 U574 ( .A(KEYINPUT47), .ZN(n630) );
  INV_X1 U575 ( .A(KEYINPUT76), .ZN(n632) );
  INV_X1 U576 ( .A(n775), .ZN(n622) );
  INV_X1 U577 ( .A(KEYINPUT4), .ZN(n468) );
  XNOR2_X1 U578 ( .A(n476), .B(n551), .ZN(n477) );
  XNOR2_X1 U579 ( .A(n580), .B(KEYINPUT34), .ZN(n581) );
  BUF_X1 U580 ( .A(n773), .Z(n774) );
  INV_X1 U581 ( .A(G134), .ZN(n469) );
  INV_X1 U582 ( .A(KEYINPUT97), .ZN(n470) );
  XOR2_X1 U583 ( .A(G140), .B(KEYINPUT79), .Z(n473) );
  XNOR2_X1 U584 ( .A(n473), .B(n472), .ZN(n476) );
  XOR2_X1 U585 ( .A(G104), .B(G107), .Z(n475) );
  NOR2_X2 U586 ( .A1(n734), .A2(G902), .ZN(n479) );
  INV_X1 U587 ( .A(G469), .ZN(n478) );
  XNOR2_X2 U588 ( .A(n479), .B(n478), .ZN(n617) );
  INV_X1 U589 ( .A(KEYINPUT65), .ZN(n480) );
  XNOR2_X1 U590 ( .A(n480), .B(KEYINPUT1), .ZN(n481) );
  NAND2_X1 U591 ( .A1(n491), .A2(G210), .ZN(n482) );
  XNOR2_X1 U592 ( .A(n482), .B(n571), .ZN(n484) );
  XOR2_X1 U593 ( .A(KEYINPUT100), .B(KEYINPUT5), .Z(n483) );
  XNOR2_X1 U594 ( .A(n484), .B(n483), .ZN(n487) );
  XNOR2_X1 U595 ( .A(n487), .B(n550), .ZN(n488) );
  XNOR2_X1 U596 ( .A(n702), .B(KEYINPUT6), .ZN(n568) );
  INV_X1 U597 ( .A(n489), .ZN(n490) );
  XNOR2_X1 U598 ( .A(n763), .B(G146), .ZN(n525) );
  XOR2_X1 U599 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n493) );
  NAND2_X1 U600 ( .A1(G214), .A2(n491), .ZN(n492) );
  XNOR2_X1 U601 ( .A(n493), .B(n492), .ZN(n497) );
  XOR2_X1 U602 ( .A(G122), .B(G104), .Z(n495) );
  XNOR2_X1 U603 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U604 ( .A(n497), .B(n496), .ZN(n500) );
  XOR2_X1 U605 ( .A(n498), .B(KEYINPUT102), .Z(n499) );
  XNOR2_X1 U606 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U607 ( .A(n525), .B(n501), .ZN(n667) );
  NAND2_X1 U608 ( .A1(n667), .A2(n538), .ZN(n505) );
  XOR2_X1 U609 ( .A(KEYINPUT104), .B(KEYINPUT13), .Z(n503) );
  XNOR2_X1 U610 ( .A(KEYINPUT103), .B(G475), .ZN(n502) );
  XNOR2_X1 U611 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U612 ( .A(n505), .B(n504), .ZN(n591) );
  XNOR2_X1 U613 ( .A(KEYINPUT105), .B(G478), .ZN(n513) );
  NAND2_X1 U614 ( .A1(n526), .A2(G217), .ZN(n512) );
  XOR2_X1 U615 ( .A(G122), .B(KEYINPUT7), .Z(n508) );
  XNOR2_X1 U616 ( .A(n512), .B(n511), .ZN(n740) );
  XNOR2_X1 U617 ( .A(n513), .B(n368), .ZN(n582) );
  INV_X1 U618 ( .A(n582), .ZN(n590) );
  OR2_X1 U619 ( .A1(n591), .A2(n590), .ZN(n684) );
  XNOR2_X1 U620 ( .A(n514), .B(n538), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n553), .A2(G234), .ZN(n515) );
  XNOR2_X1 U622 ( .A(n515), .B(KEYINPUT20), .ZN(n530) );
  AND2_X1 U623 ( .A1(n530), .A2(G221), .ZN(n517) );
  XNOR2_X1 U624 ( .A(KEYINPUT99), .B(KEYINPUT21), .ZN(n516) );
  XNOR2_X1 U625 ( .A(n517), .B(n516), .ZN(n699) );
  XOR2_X1 U626 ( .A(KEYINPUT14), .B(KEYINPUT95), .Z(n519) );
  XNOR2_X1 U627 ( .A(n519), .B(n518), .ZN(n520) );
  NAND2_X1 U628 ( .A1(G952), .A2(n520), .ZN(n725) );
  NOR2_X1 U629 ( .A1(n725), .A2(G953), .ZN(n563) );
  NAND2_X1 U630 ( .A1(G902), .A2(n520), .ZN(n561) );
  NOR2_X1 U631 ( .A1(G900), .A2(n521), .ZN(n522) );
  NOR2_X1 U632 ( .A1(n563), .A2(n522), .ZN(n523) );
  XOR2_X1 U633 ( .A(KEYINPUT84), .B(n523), .Z(n606) );
  INV_X1 U634 ( .A(n606), .ZN(n524) );
  NOR2_X1 U635 ( .A1(n699), .A2(n524), .ZN(n535) );
  XNOR2_X1 U636 ( .A(n525), .B(KEYINPUT23), .ZN(n529) );
  NAND2_X1 U637 ( .A1(G217), .A2(n530), .ZN(n531) );
  INV_X1 U638 ( .A(KEYINPUT25), .ZN(n532) );
  NAND2_X1 U639 ( .A1(n535), .A2(n698), .ZN(n614) );
  OR2_X1 U640 ( .A1(n684), .A2(n614), .ZN(n536) );
  NOR2_X1 U641 ( .A1(n568), .A2(n536), .ZN(n539) );
  NAND2_X1 U642 ( .A1(n538), .A2(n537), .ZN(n554) );
  NAND2_X1 U643 ( .A1(n554), .A2(G214), .ZN(n612) );
  NAND2_X1 U644 ( .A1(n539), .A2(n612), .ZN(n634) );
  OR2_X1 U645 ( .A1(n696), .A2(n634), .ZN(n540) );
  XNOR2_X1 U646 ( .A(KEYINPUT43), .B(n540), .ZN(n556) );
  XNOR2_X1 U647 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n542) );
  XNOR2_X1 U648 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U649 ( .A(n544), .B(n543), .ZN(n548) );
  XNOR2_X1 U650 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U651 ( .A(n548), .B(n547), .ZN(n552) );
  XNOR2_X1 U652 ( .A(KEYINPUT16), .B(G122), .ZN(n549) );
  INV_X1 U653 ( .A(n553), .ZN(n644) );
  NAND2_X1 U654 ( .A1(n554), .A2(G210), .ZN(n555) );
  AND2_X1 U655 ( .A1(n556), .A2(n633), .ZN(n641) );
  XOR2_X1 U656 ( .A(G140), .B(KEYINPUT117), .Z(n557) );
  XOR2_X1 U657 ( .A(n641), .B(n557), .Z(G42) );
  INV_X1 U658 ( .A(KEYINPUT67), .ZN(n559) );
  XNOR2_X1 U659 ( .A(n559), .B(KEYINPUT19), .ZN(n560) );
  XOR2_X1 U660 ( .A(KEYINPUT96), .B(G898), .Z(n751) );
  NAND2_X1 U661 ( .A1(G953), .A2(n751), .ZN(n758) );
  NOR2_X1 U662 ( .A1(n561), .A2(n758), .ZN(n562) );
  OR2_X1 U663 ( .A1(n563), .A2(n562), .ZN(n564) );
  INV_X1 U664 ( .A(KEYINPUT91), .ZN(n565) );
  AND2_X1 U665 ( .A1(n591), .A2(n582), .ZN(n714) );
  INV_X1 U666 ( .A(n699), .ZN(n566) );
  INV_X1 U667 ( .A(KEYINPUT22), .ZN(n567) );
  INV_X1 U668 ( .A(n568), .ZN(n578) );
  NOR2_X1 U669 ( .A1(n696), .A2(n698), .ZN(n569) );
  XNOR2_X1 U670 ( .A(n570), .B(KEYINPUT107), .ZN(n596) );
  XNOR2_X1 U671 ( .A(n596), .B(n571), .ZN(G3) );
  INV_X1 U672 ( .A(KEYINPUT92), .ZN(n572) );
  XNOR2_X1 U673 ( .A(n696), .B(n572), .ZN(n637) );
  NOR2_X1 U674 ( .A1(n637), .A2(n578), .ZN(n573) );
  NAND2_X1 U675 ( .A1(n584), .A2(n573), .ZN(n575) );
  XNOR2_X1 U676 ( .A(KEYINPUT82), .B(KEYINPUT32), .ZN(n574) );
  NAND2_X1 U677 ( .A1(n586), .A2(n578), .ZN(n579) );
  XOR2_X1 U678 ( .A(KEYINPUT81), .B(KEYINPUT74), .Z(n580) );
  OR2_X1 U679 ( .A1(n591), .A2(n582), .ZN(n625) );
  NOR2_X1 U680 ( .A1(n696), .A2(n702), .ZN(n583) );
  NAND2_X1 U681 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U682 ( .A1(n773), .A2(KEYINPUT44), .ZN(n595) );
  BUF_X1 U683 ( .A(n586), .Z(n587) );
  NAND2_X1 U684 ( .A1(n587), .A2(n702), .ZN(n706) );
  XNOR2_X1 U685 ( .A(n588), .B(KEYINPUT31), .ZN(n686) );
  NAND2_X1 U686 ( .A1(n605), .A2(n615), .ZN(n589) );
  XNOR2_X1 U687 ( .A(n372), .B(KEYINPUT101), .ZN(n673) );
  NAND2_X1 U688 ( .A1(n686), .A2(n673), .ZN(n593) );
  AND2_X1 U689 ( .A1(n591), .A2(n590), .ZN(n638) );
  NAND2_X1 U690 ( .A1(n687), .A2(n684), .ZN(n592) );
  NAND2_X1 U691 ( .A1(n593), .A2(n716), .ZN(n594) );
  NAND2_X1 U692 ( .A1(n595), .A2(n594), .ZN(n597) );
  NOR2_X1 U693 ( .A1(n597), .A2(n596), .ZN(n599) );
  XNOR2_X1 U694 ( .A(n599), .B(n598), .ZN(n600) );
  NAND2_X1 U695 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U696 ( .A1(n647), .A2(n644), .ZN(n604) );
  INV_X1 U697 ( .A(KEYINPUT86), .ZN(n603) );
  XNOR2_X1 U698 ( .A(n604), .B(n603), .ZN(n643) );
  XOR2_X1 U699 ( .A(KEYINPUT73), .B(KEYINPUT39), .Z(n609) );
  NAND2_X1 U700 ( .A1(n612), .A2(n702), .ZN(n607) );
  INV_X1 U701 ( .A(n684), .ZN(n610) );
  NAND2_X1 U702 ( .A1(n714), .A2(n715), .ZN(n613) );
  XOR2_X1 U703 ( .A(KEYINPUT41), .B(n613), .Z(n694) );
  NOR2_X1 U704 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U705 ( .A(KEYINPUT28), .B(n616), .ZN(n620) );
  XNOR2_X1 U706 ( .A(n618), .B(KEYINPUT110), .ZN(n619) );
  XNOR2_X1 U707 ( .A(n621), .B(KEYINPUT42), .ZN(n775) );
  NAND2_X1 U708 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U709 ( .A1(n633), .A2(n625), .ZN(n626) );
  AND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(n679) );
  XNOR2_X1 U711 ( .A(n369), .B(n630), .ZN(n631) );
  NOR2_X1 U712 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U713 ( .A(KEYINPUT36), .B(n635), .Z(n636) );
  NOR2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n690) );
  INV_X1 U715 ( .A(KEYINPUT112), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n640), .B(n639), .ZN(n776) );
  NOR2_X1 U717 ( .A1(n776), .A2(n641), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n765), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n644), .A2(KEYINPUT2), .ZN(n645) );
  NAND2_X1 U720 ( .A1(n646), .A2(n645), .ZN(n651) );
  BUF_X1 U721 ( .A(n647), .Z(n648) );
  XNOR2_X1 U722 ( .A(n649), .B(KEYINPUT87), .ZN(n650) );
  NAND2_X1 U723 ( .A1(n733), .A2(G472), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n652), .B(KEYINPUT62), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n654), .B(n653), .ZN(n655) );
  NAND2_X1 U726 ( .A1(n655), .A2(n663), .ZN(n657) );
  XOR2_X1 U727 ( .A(KEYINPUT113), .B(KEYINPUT63), .Z(n656) );
  XNOR2_X1 U728 ( .A(n657), .B(n656), .ZN(G57) );
  XOR2_X1 U729 ( .A(KEYINPUT122), .B(KEYINPUT54), .Z(n658) );
  XNOR2_X1 U730 ( .A(n658), .B(KEYINPUT55), .ZN(n659) );
  XOR2_X1 U731 ( .A(n660), .B(n659), .Z(n661) );
  XNOR2_X1 U732 ( .A(n662), .B(n661), .ZN(n664) );
  INV_X1 U733 ( .A(n663), .ZN(n747) );
  XNOR2_X1 U734 ( .A(n665), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U735 ( .A1(n733), .A2(G475), .ZN(n669) );
  XNOR2_X1 U736 ( .A(KEYINPUT66), .B(KEYINPUT59), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X2 U739 ( .A1(n670), .A2(n747), .ZN(n671) );
  XNOR2_X1 U740 ( .A(n671), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X1 U741 ( .A1(n684), .A2(n673), .ZN(n672) );
  XOR2_X1 U742 ( .A(G104), .B(n672), .Z(G6) );
  NOR2_X1 U743 ( .A1(n687), .A2(n673), .ZN(n675) );
  XNOR2_X1 U744 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U746 ( .A(G107), .B(n676), .ZN(G9) );
  NOR2_X1 U747 ( .A1(n680), .A2(n687), .ZN(n678) );
  XNOR2_X1 U748 ( .A(G128), .B(KEYINPUT29), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n678), .B(n677), .ZN(G30) );
  XOR2_X1 U750 ( .A(G143), .B(n679), .Z(G45) );
  NOR2_X1 U751 ( .A1(n680), .A2(n684), .ZN(n682) );
  XNOR2_X1 U752 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n681) );
  XNOR2_X1 U753 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U754 ( .A(G146), .B(n683), .ZN(G48) );
  NOR2_X1 U755 ( .A1(n684), .A2(n686), .ZN(n685) );
  XOR2_X1 U756 ( .A(G113), .B(n685), .Z(G15) );
  NOR2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U758 ( .A(KEYINPUT116), .B(n688), .Z(n689) );
  XNOR2_X1 U759 ( .A(G116), .B(n689), .ZN(G18) );
  XNOR2_X1 U760 ( .A(G125), .B(n690), .ZN(n691) );
  XNOR2_X1 U761 ( .A(n691), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U762 ( .A1(n648), .A2(n765), .ZN(n692) );
  NAND2_X1 U763 ( .A1(n692), .A2(n350), .ZN(n693) );
  INV_X1 U764 ( .A(n694), .ZN(n727) );
  OR2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U766 ( .A(KEYINPUT50), .B(n697), .ZN(n704) );
  NAND2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U768 ( .A(KEYINPUT49), .B(n700), .ZN(n701) );
  NOR2_X1 U769 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U770 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U771 ( .A(n705), .B(KEYINPUT118), .ZN(n707) );
  NAND2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U773 ( .A(KEYINPUT51), .B(n708), .Z(n709) );
  NAND2_X1 U774 ( .A1(n727), .A2(n709), .ZN(n721) );
  BUF_X1 U775 ( .A(n710), .Z(n726) );
  INV_X1 U776 ( .A(n711), .ZN(n712) );
  NAND2_X1 U777 ( .A1(n712), .A2(n432), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n714), .A2(n713), .ZN(n718) );
  NAND2_X1 U779 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U780 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U781 ( .A1(n726), .A2(n719), .ZN(n720) );
  NAND2_X1 U782 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U783 ( .A(n722), .B(KEYINPUT119), .ZN(n723) );
  XNOR2_X1 U784 ( .A(n723), .B(KEYINPUT52), .ZN(n724) );
  NOR2_X1 U785 ( .A1(n725), .A2(n724), .ZN(n729) );
  AND2_X1 U786 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U787 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U788 ( .A(KEYINPUT120), .B(n730), .Z(n731) );
  NAND2_X1 U789 ( .A1(n743), .A2(G469), .ZN(n738) );
  XNOR2_X1 U790 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n736) );
  XNOR2_X1 U791 ( .A(n734), .B(KEYINPUT57), .ZN(n735) );
  XNOR2_X1 U792 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U793 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U794 ( .A1(n747), .A2(n739), .ZN(G54) );
  NAND2_X1 U795 ( .A1(n743), .A2(G478), .ZN(n741) );
  XNOR2_X1 U796 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U797 ( .A1(n747), .A2(n742), .ZN(G63) );
  NAND2_X1 U798 ( .A1(n743), .A2(G217), .ZN(n744) );
  XNOR2_X1 U799 ( .A(n744), .B(n745), .ZN(n746) );
  NOR2_X1 U800 ( .A1(n747), .A2(n746), .ZN(G66) );
  INV_X1 U801 ( .A(n648), .ZN(n748) );
  NOR2_X1 U802 ( .A1(n748), .A2(G953), .ZN(n754) );
  NAND2_X1 U803 ( .A1(G953), .A2(G224), .ZN(n749) );
  XOR2_X1 U804 ( .A(KEYINPUT61), .B(n749), .Z(n750) );
  NOR2_X1 U805 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U806 ( .A(n752), .B(KEYINPUT124), .ZN(n753) );
  NOR2_X1 U807 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U808 ( .A(n755), .B(KEYINPUT125), .Z(n761) );
  XOR2_X1 U809 ( .A(n757), .B(n756), .Z(n759) );
  NAND2_X1 U810 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U811 ( .A(n761), .B(n760), .ZN(G69) );
  XOR2_X1 U812 ( .A(n764), .B(n763), .Z(n767) );
  XNOR2_X1 U813 ( .A(n765), .B(n767), .ZN(n766) );
  XOR2_X1 U814 ( .A(n767), .B(G227), .Z(n768) );
  XNOR2_X1 U815 ( .A(n768), .B(KEYINPUT126), .ZN(n769) );
  NAND2_X1 U816 ( .A1(n769), .A2(G900), .ZN(n770) );
  NAND2_X1 U817 ( .A1(G953), .A2(n770), .ZN(n771) );
  NAND2_X1 U818 ( .A1(n772), .A2(n771), .ZN(G72) );
  XOR2_X1 U819 ( .A(n774), .B(G122), .Z(G24) );
  XOR2_X1 U820 ( .A(G137), .B(n775), .Z(G39) );
  XOR2_X1 U821 ( .A(G134), .B(n776), .Z(G36) );
endmodule

