//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n528, new_n529, new_n530, new_n531, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1266, new_n1267, new_n1268;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT64), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  OR2_X1    g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  AOI21_X1  g035(.A(G2105), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G137), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n463), .B1(G2104), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR3_X1   g041(.A1(new_n466), .A2(KEYINPUT65), .A3(G2105), .ZN(new_n467));
  OAI21_X1  g042(.A(G101), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n464), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n469), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n461), .A2(G136), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n464), .B1(new_n459), .B2(new_n460), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G126), .B(G2105), .C1(new_n470), .C2(new_n471), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g062(.A(G138), .B(new_n464), .C1(new_n470), .C2(new_n471), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n459), .A2(new_n460), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n464), .A2(G138), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n487), .B1(new_n489), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G543), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT5), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n495), .A2(KEYINPUT66), .A3(G543), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  AND2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n502), .A2(G543), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n503), .A2(G88), .B1(G50), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(G62), .ZN(new_n506));
  NAND2_X1  g081(.A1(G75), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G651), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT67), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n505), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n501), .A2(new_n502), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n502), .A2(G543), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n517), .B1(new_n506), .B2(new_n507), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT67), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n511), .A2(new_n519), .ZN(G166));
  NAND2_X1  g095(.A1(new_n503), .A2(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n501), .A2(G63), .A3(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n504), .A2(G51), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n521), .A2(new_n522), .A3(new_n524), .A4(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  XOR2_X1   g102(.A(KEYINPUT68), .B(G90), .Z(new_n528));
  NAND2_X1  g103(.A1(new_n503), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n501), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  OAI221_X1 g106(.A(new_n529), .B1(new_n530), .B2(new_n515), .C1(new_n517), .C2(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  NAND2_X1  g108(.A1(new_n504), .A2(G43), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT70), .B(G81), .Z(new_n535));
  NAND3_X1  g110(.A1(new_n501), .A2(new_n502), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n538));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n540), .B1(new_n501), .B2(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n538), .B1(new_n541), .B2(new_n517), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n495), .A2(KEYINPUT66), .A3(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(KEYINPUT66), .B1(new_n495), .B2(G543), .ZN(new_n545));
  OAI211_X1 g120(.A(G56), .B(new_n543), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(new_n539), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n547), .A2(KEYINPUT69), .A3(G651), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n537), .B1(new_n542), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND3_X1  g129(.A1(new_n501), .A2(G91), .A3(new_n502), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT74), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n501), .A2(new_n557), .A3(G91), .A4(new_n502), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n499), .A2(new_n500), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n559), .A2(G65), .A3(new_n543), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n556), .A2(new_n558), .B1(new_n562), .B2(G651), .ZN(new_n563));
  AND2_X1   g138(.A1(G53), .A2(G543), .ZN(new_n564));
  AND2_X1   g139(.A1(KEYINPUT6), .A2(G651), .ZN(new_n565));
  NOR2_X1   g140(.A1(KEYINPUT6), .A2(G651), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n568));
  AND2_X1   g143(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n569));
  NOR2_X1   g144(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n568), .B(KEYINPUT72), .C1(new_n567), .C2(new_n571), .ZN(new_n572));
  XNOR2_X1  g147(.A(KEYINPUT71), .B(KEYINPUT9), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n502), .A2(new_n573), .A3(new_n574), .A4(new_n564), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT73), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT72), .B1(new_n567), .B2(new_n571), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n502), .B2(new_n564), .ZN(new_n579));
  OAI211_X1 g154(.A(KEYINPUT73), .B(new_n575), .C1(new_n577), .C2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n563), .B1(new_n576), .B2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G166), .ZN(G303));
  NAND2_X1  g158(.A1(new_n504), .A2(G49), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n501), .B2(G74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n501), .A2(G87), .A3(new_n502), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(new_n501), .A2(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT75), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n517), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n501), .A2(G86), .A3(new_n502), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n502), .A2(G48), .A3(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n501), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n517), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  XOR2_X1   g174(.A(KEYINPUT76), .B(G47), .Z(new_n600));
  OAI22_X1  g175(.A1(new_n512), .A2(new_n599), .B1(new_n515), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G290));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NOR2_X1   g179(.A1(G301), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n501), .A2(G66), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n504), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n512), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n501), .A2(KEYINPUT10), .A3(G92), .A4(new_n502), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n609), .A2(new_n614), .A3(KEYINPUT77), .ZN(new_n618));
  AND2_X1   g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n605), .B1(new_n619), .B2(new_n604), .ZN(G284));
  AOI21_X1  g195(.A(new_n605), .B1(new_n619), .B2(new_n604), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  INV_X1    g197(.A(G299), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G868), .ZN(G297));
  XNOR2_X1  g199(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(G860), .ZN(G148));
  AND2_X1   g202(.A1(new_n534), .A2(new_n536), .ZN(new_n628));
  AOI21_X1  g203(.A(KEYINPUT69), .B1(new_n547), .B2(G651), .ZN(new_n629));
  AOI211_X1 g204(.A(new_n538), .B(new_n517), .C1(new_n546), .C2(new_n539), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(new_n604), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n617), .A2(new_n626), .A3(new_n618), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n632), .B1(new_n634), .B2(new_n604), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g211(.A1(new_n465), .A2(new_n467), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(new_n490), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT13), .Z(new_n641));
  INV_X1    g216(.A(G2100), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n461), .A2(G135), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n477), .A2(G123), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n464), .A2(G111), .ZN(new_n647));
  OAI21_X1  g222(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n645), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(G2096), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n643), .A2(new_n644), .A3(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(KEYINPUT14), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2451), .B(G2454), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n652), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT80), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n663), .A2(new_n664), .A3(new_n652), .ZN(new_n667));
  INV_X1    g242(.A(G14), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n666), .A2(new_n669), .ZN(G401));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT81), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT17), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2084), .B(G2090), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n675), .B1(new_n672), .B2(new_n674), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n673), .B2(new_n674), .ZN(new_n678));
  INV_X1    g253(.A(new_n674), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n679), .A2(new_n675), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n672), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT18), .ZN(new_n682));
  OR3_X1    g257(.A1(new_n676), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT83), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G1986), .ZN(new_n690));
  XOR2_X1   g265(.A(G1971), .B(G1976), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT19), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT82), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n693), .A2(new_n694), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(new_n695), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n697), .B1(new_n692), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n692), .A2(new_n698), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT20), .Z(new_n702));
  OAI21_X1  g277(.A(G1981), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n700), .A2(G1981), .A3(new_n702), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n690), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n705), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n707), .A2(G1986), .A3(new_n703), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n689), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1991), .B(G1996), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n706), .A2(new_n708), .A3(new_n689), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n711), .ZN(new_n714));
  INV_X1    g289(.A(new_n712), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n709), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n713), .A2(new_n716), .ZN(G229));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NOR2_X1   g293(.A1(G168), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n718), .B2(G21), .ZN(new_n720));
  INV_X1    g295(.A(G1966), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT30), .B(G28), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  OR2_X1    g300(.A1(KEYINPUT31), .A2(G11), .ZN(new_n726));
  NAND2_X1  g301(.A1(KEYINPUT31), .A2(G11), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n724), .A2(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n649), .B2(new_n725), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n725), .B1(KEYINPUT24), .B2(G34), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(KEYINPUT24), .B2(G34), .ZN(new_n731));
  INV_X1    g306(.A(G160), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G29), .ZN(new_n733));
  INV_X1    g308(.A(G2084), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n729), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n722), .A2(new_n723), .A3(new_n735), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n637), .A2(G105), .B1(G141), .B2(new_n461), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT26), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G129), .B2(new_n477), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(new_n725), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n725), .B2(G32), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(G29), .A2(G33), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT25), .Z(new_n749));
  NAND2_X1  g324(.A1(new_n461), .A2(G139), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n490), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n749), .B(new_n750), .C1(new_n464), .C2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n747), .B1(new_n752), .B2(new_n725), .ZN(new_n753));
  INV_X1    g328(.A(G2072), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n744), .A2(new_n745), .ZN(new_n756));
  NAND2_X1  g331(.A1(G164), .A2(G29), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G27), .B2(G29), .ZN(new_n758));
  INV_X1    g333(.A(G2078), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n746), .A2(new_n755), .A3(new_n756), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n725), .A2(G35), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G162), .B2(new_n725), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT29), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n764), .A2(G2090), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n753), .A2(new_n754), .ZN(new_n766));
  OAI221_X1 g341(.A(new_n766), .B1(new_n759), .B2(new_n758), .C1(new_n734), .C2(new_n733), .ZN(new_n767));
  OR4_X1    g342(.A1(new_n736), .A2(new_n761), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G1961), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(KEYINPUT93), .ZN(new_n770));
  NOR2_X1   g345(.A1(G171), .A2(new_n718), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n718), .A2(G5), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n769), .A2(KEYINPUT93), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n718), .A2(G19), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(KEYINPUT88), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(KEYINPUT88), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n777), .B(new_n778), .C1(new_n549), .C2(new_n718), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT89), .B(G1341), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n775), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n725), .A2(G26), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n461), .A2(G140), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n477), .A2(G128), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n464), .A2(G116), .ZN(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n788), .B(new_n789), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT90), .Z(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n787), .B1(new_n794), .B2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT92), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2067), .ZN(new_n797));
  NOR3_X1   g372(.A1(new_n768), .A2(new_n784), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n718), .A2(G4), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n619), .B2(new_n718), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT87), .B(G1348), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n718), .A2(G20), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT23), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n623), .B2(new_n718), .ZN(new_n805));
  INV_X1    g380(.A(G1956), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n764), .A2(G2090), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT94), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n798), .A2(new_n802), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G303), .A2(new_n718), .ZN(new_n812));
  NOR2_X1   g387(.A1(G16), .A2(G22), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT86), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G1971), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n812), .A2(KEYINPUT86), .A3(new_n813), .ZN(new_n818));
  OR3_X1    g393(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT34), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n817), .B1(new_n816), .B2(new_n818), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n718), .A2(G23), .ZN(new_n822));
  INV_X1    g397(.A(G288), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(new_n718), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT33), .B(G1976), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(G6), .A2(G16), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n595), .B2(G16), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT32), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G1981), .ZN(new_n833));
  INV_X1    g408(.A(G1981), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n830), .A2(new_n834), .A3(new_n831), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n826), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n461), .A2(G131), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n477), .A2(G119), .ZN(new_n839));
  OR2_X1    g414(.A1(G95), .A2(G2105), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n840), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  MUX2_X1   g417(.A(G25), .B(new_n842), .S(G29), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT84), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT35), .B(G1991), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n718), .A2(G24), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n602), .A2(KEYINPUT85), .ZN(new_n848));
  OAI21_X1  g423(.A(G16), .B1(new_n602), .B2(KEYINPUT85), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n846), .B1(G1986), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G1986), .B2(new_n850), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n837), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n819), .A2(new_n821), .A3(new_n836), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(KEYINPUT34), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT36), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT36), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n853), .A2(new_n858), .A3(new_n855), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n811), .B1(new_n857), .B2(new_n859), .ZN(G311));
  INV_X1    g435(.A(new_n811), .ZN(new_n861));
  INV_X1    g436(.A(new_n859), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n858), .B1(new_n853), .B2(new_n855), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(G150));
  NAND2_X1  g439(.A1(new_n501), .A2(G67), .ZN(new_n865));
  NAND2_X1  g440(.A1(G80), .A2(G543), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n517), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n559), .A2(G93), .A3(new_n543), .A4(new_n502), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n502), .A2(G55), .A3(G543), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT95), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT95), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n868), .A2(new_n872), .A3(new_n869), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n867), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT96), .B(G860), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n619), .A2(G559), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT38), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n865), .A2(new_n866), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(G651), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n868), .A2(new_n872), .A3(new_n869), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n872), .B1(new_n868), .B2(new_n869), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n631), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n549), .A2(new_n874), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n880), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n878), .B(KEYINPUT38), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n887), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n891), .A3(KEYINPUT39), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT97), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT97), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n888), .A2(new_n891), .A3(new_n894), .A4(KEYINPUT39), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT39), .B1(new_n888), .B2(new_n891), .ZN(new_n897));
  INV_X1    g472(.A(new_n875), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n896), .A2(KEYINPUT98), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT98), .B1(new_n896), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n877), .B1(new_n900), .B2(new_n901), .ZN(G145));
  NAND2_X1  g477(.A1(new_n489), .A2(new_n493), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n483), .A2(new_n486), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n741), .B(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n906), .A2(new_n793), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n906), .A2(new_n793), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n752), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT99), .ZN(new_n911));
  OR3_X1    g486(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n911), .B1(new_n907), .B2(new_n908), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n461), .A2(G142), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n477), .A2(G130), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n464), .A2(G118), .ZN(new_n917));
  OAI21_X1  g492(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n915), .B(new_n916), .C1(new_n917), .C2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT102), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n920), .A2(new_n640), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n842), .B(KEYINPUT101), .Z(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n640), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n922), .B2(new_n924), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n914), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n912), .B(new_n913), .C1(new_n925), .C2(new_n926), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(G160), .B(new_n649), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(G162), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n914), .A2(KEYINPUT103), .A3(new_n927), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G37), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n914), .B2(new_n927), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n937), .A2(KEYINPUT104), .A3(new_n930), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT104), .B1(new_n937), .B2(new_n930), .ZN(new_n939));
  OAI211_X1 g514(.A(new_n935), .B(new_n936), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g516(.A1(G166), .A2(new_n823), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(G166), .A2(new_n823), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n602), .B(new_n595), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n943), .B2(new_n944), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  XOR2_X1   g524(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(G299), .A2(new_n615), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n575), .B1(new_n577), .B2(new_n579), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT73), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n580), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n956), .A2(new_n563), .B1(new_n614), .B2(new_n609), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT41), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n609), .A2(new_n614), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n959), .A2(new_n563), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g535(.A1(G299), .A2(new_n615), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT41), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n958), .A2(KEYINPUT105), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n960), .A2(new_n961), .A3(new_n965), .A4(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n634), .A2(new_n890), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n633), .A2(new_n886), .A3(new_n887), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n952), .A2(new_n957), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n968), .A2(new_n973), .A3(new_n969), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n951), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n964), .A2(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n968), .A2(new_n973), .A3(new_n969), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n976), .A2(new_n977), .A3(new_n950), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n949), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n971), .A2(new_n951), .A3(new_n974), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n950), .B1(new_n976), .B2(new_n977), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n981), .A3(new_n948), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n604), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n874), .A2(G868), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n983), .A2(KEYINPUT107), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n980), .A2(new_n981), .A3(new_n948), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n948), .B1(new_n980), .B2(new_n981), .ZN(new_n988));
  OAI21_X1  g563(.A(G868), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n984), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n985), .A2(new_n991), .ZN(G295));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n990), .ZN(G331));
  AND3_X1   g568(.A1(new_n886), .A2(new_n887), .A3(G301), .ZN(new_n994));
  AOI21_X1  g569(.A(G301), .B1(new_n886), .B2(new_n887), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n994), .A2(new_n995), .A3(G286), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n549), .A2(new_n874), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n631), .A2(new_n885), .ZN(new_n998));
  OAI21_X1  g573(.A(G171), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n886), .A2(new_n887), .A3(G301), .ZN(new_n1000));
  AOI21_X1  g575(.A(G168), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n972), .B1(new_n996), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(G286), .B1(new_n994), .B2(new_n995), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n999), .A2(G168), .A3(new_n1000), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n964), .A2(new_n1003), .A3(new_n1004), .A4(new_n966), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1005), .A3(new_n948), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT108), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n949), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1002), .A2(new_n1005), .A3(new_n1010), .A4(new_n948), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1007), .A2(new_n1009), .A3(new_n936), .A4(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT43), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(G37), .B1(new_n1006), .B2(KEYINPUT108), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n973), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n958), .A2(new_n1017), .A3(new_n963), .ZN(new_n1018));
  AND4_X1   g593(.A1(new_n1004), .A2(new_n1016), .A3(new_n1003), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1002), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n949), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AND4_X1   g596(.A1(KEYINPUT43), .A2(new_n1015), .A3(new_n1011), .A4(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT44), .B1(new_n1014), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1015), .A2(new_n1021), .A3(new_n1013), .A4(new_n1011), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1023), .A2(new_n1028), .ZN(G397));
  XNOR2_X1  g604(.A(new_n793), .B(G2067), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(G164), .B2(G1384), .ZN(new_n1032));
  INV_X1    g607(.A(new_n469), .ZN(new_n1033));
  INV_X1    g608(.A(new_n474), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(G40), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1030), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT111), .ZN(new_n1039));
  INV_X1    g614(.A(new_n845), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n842), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n842), .A2(new_n1040), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1036), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1036), .A2(G1996), .A3(new_n741), .ZN(new_n1044));
  OR3_X1    g619(.A1(new_n1032), .A2(new_n1035), .A3(G1996), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n1045), .B(KEYINPUT110), .Z(new_n1046));
  AOI21_X1  g621(.A(new_n1044), .B1(new_n1046), .B2(new_n742), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1039), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1048));
  NOR2_X1   g623(.A1(G290), .A2(G1986), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G290), .A2(G1986), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1037), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n511), .A2(G8), .A3(new_n519), .ZN(new_n1054));
  NAND2_X1  g629(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1055));
  NOR2_X1   g630(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT114), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1057), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1384), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n905), .A2(KEYINPUT112), .A3(KEYINPUT45), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(KEYINPUT45), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1063), .B1(G164), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G40), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n469), .A2(new_n1066), .A3(new_n474), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1062), .A2(new_n1032), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1068), .A2(new_n817), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT50), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n905), .A2(new_n1070), .A3(new_n1061), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(G1384), .B1(new_n903), .B2(new_n904), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(KEYINPUT118), .A3(new_n1070), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1067), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(KEYINPUT117), .A3(new_n1067), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1076), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G2090), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1069), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G8), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1060), .B(KEYINPUT119), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n1087));
  NOR4_X1   g662(.A1(G164), .A2(new_n1072), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1088));
  AOI21_X1  g663(.A(KEYINPUT118), .B1(new_n1074), .B2(new_n1070), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1081), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT117), .B1(new_n1077), .B2(new_n1067), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1090), .B(new_n1083), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1068), .A2(new_n817), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1085), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1087), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT49), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n588), .A2(new_n590), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(G651), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n592), .A2(new_n593), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n834), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n591), .A2(new_n594), .A3(G1981), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1098), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1085), .B1(new_n1067), .B2(new_n1074), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(new_n1101), .A3(new_n834), .ZN(new_n1106));
  OAI21_X1  g681(.A(G1981), .B1(new_n591), .B2(new_n594), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(KEYINPUT49), .A3(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n1105), .A3(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n584), .A2(new_n585), .A3(G1976), .A4(new_n586), .ZN(new_n1110));
  INV_X1    g685(.A(G1976), .ZN(new_n1111));
  AOI21_X1  g686(.A(KEYINPUT52), .B1(G288), .B2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1105), .A2(KEYINPUT115), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n905), .A2(new_n1061), .ZN(new_n1115));
  OAI211_X1 g690(.A(G8), .B(new_n1110), .C1(new_n1115), .C2(new_n1035), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1114), .B1(new_n1116), .B2(KEYINPUT52), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1105), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1109), .B(new_n1113), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1077), .A2(new_n1071), .A3(new_n1067), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1083), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1085), .B1(new_n1121), .B2(new_n1094), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1119), .B1(new_n1096), .B2(new_n1122), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1086), .A2(new_n1097), .A3(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(G301), .B(KEYINPUT54), .Z(new_n1125));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1035), .B1(new_n1115), .B2(KEYINPUT50), .ZN(new_n1127));
  AOI21_X1  g702(.A(G1961), .B1(new_n1127), .B2(new_n1071), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n905), .A2(KEYINPUT45), .A3(new_n1061), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1130), .A2(G2078), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1032), .A2(new_n1129), .A3(new_n1067), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1126), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT126), .B(new_n1132), .C1(new_n1120), .C2(G1961), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1130), .B1(new_n1068), .B2(G2078), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1125), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1128), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1033), .A2(G40), .A3(new_n1131), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n472), .A2(new_n473), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1141), .A2(KEYINPUT127), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n464), .B1(new_n1141), .B2(KEYINPUT127), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1140), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1144), .A2(new_n1062), .A3(new_n1032), .A4(new_n1065), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1125), .A2(new_n1139), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1138), .B1(new_n1137), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(G286), .A2(G8), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1067), .B1(G164), .B2(new_n1064), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1074), .A2(KEYINPUT45), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT120), .B(new_n721), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1077), .A2(new_n1071), .A3(new_n734), .A4(new_n1067), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1032), .A2(new_n1129), .A3(new_n1067), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT120), .B1(new_n1155), .B2(new_n721), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1149), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n721), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1160), .A2(KEYINPUT125), .A3(new_n1153), .A4(new_n1152), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1148), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1157), .A2(G168), .A3(new_n1161), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT51), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1164), .A2(new_n1085), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1160), .A2(new_n1153), .A3(new_n1152), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(G8), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1163), .A2(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1124), .B(new_n1147), .C1(new_n1162), .C2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n1171));
  INV_X1    g746(.A(new_n953), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n563), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT57), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT123), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1175), .B(new_n1176), .C1(new_n1174), .C2(G299), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n623), .A2(KEYINPUT123), .A3(KEYINPUT57), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT122), .B1(new_n1082), .B2(G1956), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1182), .A2(new_n1183), .A3(new_n806), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  XOR2_X1   g760(.A(KEYINPUT56), .B(G2072), .Z(new_n1186));
  NOR2_X1   g761(.A1(new_n1068), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1180), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  AOI211_X1 g764(.A(new_n1187), .B(new_n1179), .C1(new_n1181), .C2(new_n1184), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1171), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1082), .A2(KEYINPUT122), .A3(G1956), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1183), .B1(new_n1182), .B2(new_n806), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1188), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1194), .A2(new_n1179), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1185), .A2(new_n1180), .A3(new_n1188), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1195), .A2(KEYINPUT61), .A3(new_n1196), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1115), .A2(new_n1035), .ZN(new_n1198));
  XNOR2_X1  g773(.A(KEYINPUT58), .B(G1341), .ZN(new_n1199));
  OAI22_X1  g774(.A1(new_n1068), .A2(G1996), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n549), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT59), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1201), .B(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(G2067), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1198), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1205), .B1(new_n1120), .B2(G1348), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1207), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT60), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1209), .B1(new_n1206), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n615), .B1(new_n1206), .B2(new_n1210), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1213), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1215), .A2(new_n1211), .A3(new_n1208), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1203), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1191), .A2(new_n1197), .A3(new_n1217), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1207), .A2(new_n615), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1196), .B1(new_n1189), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1170), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g799(.A(new_n1162), .ZN(new_n1225));
  INV_X1    g800(.A(KEYINPUT62), .ZN(new_n1226));
  NAND3_X1  g801(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OAI21_X1  g802(.A(KEYINPUT62), .B1(new_n1169), .B2(new_n1162), .ZN(new_n1228));
  AOI21_X1  g803(.A(G301), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1229));
  AND4_X1   g804(.A1(new_n1097), .A2(new_n1086), .A3(new_n1229), .A4(new_n1123), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1227), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  NAND3_X1  g806(.A1(new_n1166), .A2(G8), .A3(G168), .ZN(new_n1232));
  INV_X1    g807(.A(new_n1232), .ZN(new_n1233));
  NAND4_X1  g808(.A1(new_n1086), .A2(new_n1097), .A3(new_n1123), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g809(.A(KEYINPUT63), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OR2_X1    g811(.A1(new_n1122), .A2(KEYINPUT121), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1122), .A2(KEYINPUT121), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n1237), .A2(new_n1060), .A3(new_n1238), .ZN(new_n1239));
  NAND4_X1  g814(.A1(new_n1239), .A2(KEYINPUT63), .A3(new_n1123), .A4(new_n1233), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1236), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g816(.A(new_n1122), .ZN(new_n1242));
  NOR3_X1   g817(.A1(new_n1060), .A2(new_n1242), .A3(new_n1119), .ZN(new_n1243));
  NAND3_X1  g818(.A1(new_n1109), .A2(new_n1111), .A3(new_n823), .ZN(new_n1244));
  XNOR2_X1  g819(.A(new_n1106), .B(KEYINPUT116), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g821(.A(new_n1243), .B1(new_n1105), .B2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g822(.A1(new_n1231), .A2(new_n1241), .A3(new_n1247), .ZN(new_n1248));
  OAI21_X1  g823(.A(new_n1053), .B1(new_n1221), .B2(new_n1248), .ZN(new_n1249));
  INV_X1    g824(.A(KEYINPUT46), .ZN(new_n1250));
  XNOR2_X1  g825(.A(new_n1046), .B(new_n1250), .ZN(new_n1251));
  INV_X1    g826(.A(new_n1030), .ZN(new_n1252));
  OAI21_X1  g827(.A(new_n1036), .B1(new_n1252), .B2(new_n741), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1251), .A2(new_n1253), .ZN(new_n1254));
  AND2_X1   g829(.A1(new_n1254), .A2(KEYINPUT47), .ZN(new_n1255));
  NOR2_X1   g830(.A1(new_n1254), .A2(KEYINPUT47), .ZN(new_n1256));
  NAND2_X1  g831(.A1(new_n1049), .A2(new_n1036), .ZN(new_n1257));
  XOR2_X1   g832(.A(new_n1257), .B(KEYINPUT48), .Z(new_n1258));
  OAI22_X1  g833(.A1(new_n1255), .A2(new_n1256), .B1(new_n1048), .B2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g834(.A1(new_n1039), .A2(new_n1042), .A3(new_n1047), .ZN(new_n1260));
  NAND2_X1  g835(.A1(new_n793), .A2(new_n1204), .ZN(new_n1261));
  AOI21_X1  g836(.A(new_n1037), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g837(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g838(.A1(new_n1249), .A2(new_n1263), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g839(.A1(new_n685), .A2(G319), .ZN(new_n1266));
  AOI21_X1  g840(.A(new_n1266), .B1(new_n666), .B2(new_n669), .ZN(new_n1267));
  AND3_X1   g841(.A1(new_n713), .A2(new_n716), .A3(new_n1267), .ZN(new_n1268));
  NAND3_X1  g842(.A1(new_n1026), .A2(new_n940), .A3(new_n1268), .ZN(G225));
  INV_X1    g843(.A(G225), .ZN(G308));
endmodule


