

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n731), .A2(n730), .ZN(n732) );
  INV_X1 U549 ( .A(n676), .ZN(n704) );
  INV_X1 U550 ( .A(KEYINPUT29), .ZN(n702) );
  XNOR2_X1 U551 ( .A(n703), .B(n702), .ZN(n709) );
  BUF_X1 U552 ( .A(n676), .Z(n720) );
  NOR2_X1 U553 ( .A1(G651), .A2(n621), .ZN(n631) );
  XOR2_X1 U554 ( .A(KEYINPUT17), .B(n530), .Z(n876) );
  NOR2_X1 U555 ( .A1(n538), .A2(n537), .ZN(G160) );
  INV_X1 U556 ( .A(G651), .ZN(n521) );
  XOR2_X1 U557 ( .A(KEYINPUT0), .B(G543), .Z(n621) );
  OR2_X1 U558 ( .A1(n521), .A2(n621), .ZN(n515) );
  XNOR2_X1 U559 ( .A(KEYINPUT65), .B(n515), .ZN(n634) );
  NAND2_X1 U560 ( .A1(n634), .A2(G76), .ZN(n516) );
  XNOR2_X1 U561 ( .A(KEYINPUT70), .B(n516), .ZN(n519) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n630) );
  NAND2_X1 U563 ( .A1(n630), .A2(G89), .ZN(n517) );
  XNOR2_X1 U564 ( .A(KEYINPUT4), .B(n517), .ZN(n518) );
  NAND2_X1 U565 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U566 ( .A(n520), .B(KEYINPUT5), .ZN(n528) );
  XNOR2_X1 U567 ( .A(KEYINPUT71), .B(KEYINPUT6), .ZN(n526) );
  NOR2_X1 U568 ( .A1(G543), .A2(n521), .ZN(n522) );
  XOR2_X1 U569 ( .A(KEYINPUT1), .B(n522), .Z(n636) );
  NAND2_X1 U570 ( .A1(G63), .A2(n636), .ZN(n524) );
  NAND2_X1 U571 ( .A1(G51), .A2(n631), .ZN(n523) );
  NAND2_X1 U572 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U573 ( .A(n526), .B(n525), .ZN(n527) );
  NAND2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U575 ( .A(KEYINPUT7), .B(n529), .ZN(G168) );
  XOR2_X1 U576 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  NAND2_X1 U578 ( .A1(n876), .A2(G137), .ZN(n533) );
  XOR2_X1 U579 ( .A(G2104), .B(KEYINPUT64), .Z(n534) );
  NOR2_X4 U580 ( .A1(G2105), .A2(n534), .ZN(n877) );
  NAND2_X1 U581 ( .A1(G101), .A2(n877), .ZN(n531) );
  XOR2_X1 U582 ( .A(KEYINPUT23), .B(n531), .Z(n532) );
  NAND2_X1 U583 ( .A1(n533), .A2(n532), .ZN(n538) );
  AND2_X1 U584 ( .A1(G2105), .A2(n534), .ZN(n880) );
  NAND2_X1 U585 ( .A1(G125), .A2(n880), .ZN(n536) );
  AND2_X1 U586 ( .A1(G2105), .A2(G2104), .ZN(n881) );
  NAND2_X1 U587 ( .A1(G113), .A2(n881), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U589 ( .A1(G64), .A2(n636), .ZN(n540) );
  NAND2_X1 U590 ( .A1(G52), .A2(n631), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n545) );
  NAND2_X1 U592 ( .A1(G90), .A2(n630), .ZN(n542) );
  NAND2_X1 U593 ( .A1(G77), .A2(n634), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U595 ( .A(KEYINPUT9), .B(n543), .Z(n544) );
  NOR2_X1 U596 ( .A1(n545), .A2(n544), .ZN(G171) );
  AND2_X1 U597 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U598 ( .A(G57), .ZN(G237) );
  INV_X1 U599 ( .A(G132), .ZN(G219) );
  INV_X1 U600 ( .A(G82), .ZN(G220) );
  NAND2_X1 U601 ( .A1(G7), .A2(G661), .ZN(n546) );
  XNOR2_X1 U602 ( .A(n546), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U603 ( .A(G223), .ZN(n821) );
  NAND2_X1 U604 ( .A1(n821), .A2(G567), .ZN(n547) );
  XOR2_X1 U605 ( .A(KEYINPUT11), .B(n547), .Z(G234) );
  NAND2_X1 U606 ( .A1(G56), .A2(n636), .ZN(n548) );
  XOR2_X1 U607 ( .A(KEYINPUT14), .B(n548), .Z(n554) );
  NAND2_X1 U608 ( .A1(n630), .A2(G81), .ZN(n549) );
  XNOR2_X1 U609 ( .A(n549), .B(KEYINPUT12), .ZN(n551) );
  NAND2_X1 U610 ( .A1(G68), .A2(n634), .ZN(n550) );
  NAND2_X1 U611 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U612 ( .A(KEYINPUT13), .B(n552), .Z(n553) );
  NOR2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n631), .A2(G43), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n1002) );
  INV_X1 U616 ( .A(G860), .ZN(n605) );
  OR2_X1 U617 ( .A1(n1002), .A2(n605), .ZN(G153) );
  INV_X1 U618 ( .A(G171), .ZN(G301) );
  NAND2_X1 U619 ( .A1(G868), .A2(G301), .ZN(n566) );
  NAND2_X1 U620 ( .A1(G66), .A2(n636), .ZN(n558) );
  NAND2_X1 U621 ( .A1(G92), .A2(n630), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U623 ( .A1(G79), .A2(n634), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G54), .A2(n631), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U627 ( .A(KEYINPUT69), .B(KEYINPUT15), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n564), .B(n563), .ZN(n989) );
  OR2_X1 U629 ( .A1(n989), .A2(G868), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(G284) );
  NAND2_X1 U631 ( .A1(G65), .A2(n636), .ZN(n568) );
  NAND2_X1 U632 ( .A1(G53), .A2(n631), .ZN(n567) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n630), .A2(G91), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT66), .ZN(n571) );
  NAND2_X1 U636 ( .A1(G78), .A2(n634), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT67), .B(n572), .Z(n573) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n1001) );
  XOR2_X1 U640 ( .A(n1001), .B(KEYINPUT68), .Z(G299) );
  NOR2_X1 U641 ( .A1(G868), .A2(G299), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n575), .B(KEYINPUT72), .ZN(n577) );
  INV_X1 U643 ( .A(G868), .ZN(n651) );
  NOR2_X1 U644 ( .A1(n651), .A2(G286), .ZN(n576) );
  NOR2_X1 U645 ( .A1(n577), .A2(n576), .ZN(G297) );
  NAND2_X1 U646 ( .A1(n605), .A2(G559), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n578), .A2(n989), .ZN(n579) );
  XNOR2_X1 U648 ( .A(n579), .B(KEYINPUT73), .ZN(n580) );
  XOR2_X1 U649 ( .A(KEYINPUT16), .B(n580), .Z(G148) );
  NOR2_X1 U650 ( .A1(G868), .A2(n1002), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G868), .A2(n989), .ZN(n581) );
  NOR2_X1 U652 ( .A1(G559), .A2(n581), .ZN(n582) );
  NOR2_X1 U653 ( .A1(n583), .A2(n582), .ZN(G282) );
  XOR2_X1 U654 ( .A(G2100), .B(KEYINPUT76), .Z(n594) );
  XOR2_X1 U655 ( .A(G2096), .B(KEYINPUT75), .Z(n592) );
  NAND2_X1 U656 ( .A1(G123), .A2(n880), .ZN(n584) );
  XNOR2_X1 U657 ( .A(n584), .B(KEYINPUT18), .ZN(n585) );
  XNOR2_X1 U658 ( .A(n585), .B(KEYINPUT74), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G111), .A2(n881), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G135), .A2(n876), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G99), .A2(n877), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n965) );
  XNOR2_X1 U665 ( .A(n592), .B(n965), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n594), .A2(n593), .ZN(G156) );
  NAND2_X1 U667 ( .A1(n630), .A2(G93), .ZN(n595) );
  XNOR2_X1 U668 ( .A(n595), .B(KEYINPUT78), .ZN(n597) );
  NAND2_X1 U669 ( .A1(G80), .A2(n634), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U671 ( .A(n598), .B(KEYINPUT79), .ZN(n600) );
  NAND2_X1 U672 ( .A1(G67), .A2(n636), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U674 ( .A1(n631), .A2(G55), .ZN(n601) );
  XOR2_X1 U675 ( .A(KEYINPUT80), .B(n601), .Z(n602) );
  OR2_X1 U676 ( .A1(n603), .A2(n602), .ZN(n652) );
  NAND2_X1 U677 ( .A1(G559), .A2(n989), .ZN(n604) );
  XOR2_X1 U678 ( .A(n1002), .B(n604), .Z(n648) );
  NAND2_X1 U679 ( .A1(n605), .A2(n648), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n606), .B(KEYINPUT77), .ZN(n607) );
  XOR2_X1 U681 ( .A(n652), .B(n607), .Z(G145) );
  NAND2_X1 U682 ( .A1(n630), .A2(G86), .ZN(n608) );
  XOR2_X1 U683 ( .A(KEYINPUT81), .B(n608), .Z(n610) );
  NAND2_X1 U684 ( .A1(n636), .A2(G61), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U686 ( .A(KEYINPUT82), .B(n611), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n634), .A2(G73), .ZN(n612) );
  XOR2_X1 U688 ( .A(KEYINPUT2), .B(n612), .Z(n613) );
  NOR2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U690 ( .A1(n631), .A2(G48), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U692 ( .A(KEYINPUT83), .B(n617), .Z(G305) );
  NAND2_X1 U693 ( .A1(G49), .A2(n631), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G74), .A2(G651), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U696 ( .A1(n636), .A2(n620), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n621), .A2(G87), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(G288) );
  AND2_X1 U699 ( .A1(n630), .A2(G85), .ZN(n627) );
  NAND2_X1 U700 ( .A1(G60), .A2(n636), .ZN(n625) );
  NAND2_X1 U701 ( .A1(G47), .A2(n631), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n629) );
  NAND2_X1 U704 ( .A1(n634), .A2(G72), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(G290) );
  NAND2_X1 U706 ( .A1(G88), .A2(n630), .ZN(n633) );
  NAND2_X1 U707 ( .A1(G50), .A2(n631), .ZN(n632) );
  NAND2_X1 U708 ( .A1(n633), .A2(n632), .ZN(n640) );
  NAND2_X1 U709 ( .A1(G75), .A2(n634), .ZN(n635) );
  XNOR2_X1 U710 ( .A(n635), .B(KEYINPUT84), .ZN(n638) );
  NAND2_X1 U711 ( .A1(n636), .A2(G62), .ZN(n637) );
  NAND2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U713 ( .A1(n640), .A2(n639), .ZN(G166) );
  XNOR2_X1 U714 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n642) );
  XNOR2_X1 U715 ( .A(G288), .B(KEYINPUT86), .ZN(n641) );
  XNOR2_X1 U716 ( .A(n642), .B(n641), .ZN(n643) );
  XOR2_X1 U717 ( .A(n652), .B(n643), .Z(n645) );
  XNOR2_X1 U718 ( .A(G290), .B(G166), .ZN(n644) );
  XNOR2_X1 U719 ( .A(n645), .B(n644), .ZN(n646) );
  XOR2_X1 U720 ( .A(G299), .B(n646), .Z(n647) );
  XNOR2_X1 U721 ( .A(G305), .B(n647), .ZN(n899) );
  XNOR2_X1 U722 ( .A(n899), .B(n648), .ZN(n649) );
  NAND2_X1 U723 ( .A1(n649), .A2(G868), .ZN(n650) );
  XOR2_X1 U724 ( .A(KEYINPUT87), .B(n650), .Z(n654) );
  NAND2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(G295) );
  NAND2_X1 U727 ( .A1(G2078), .A2(G2084), .ZN(n656) );
  XOR2_X1 U728 ( .A(KEYINPUT20), .B(KEYINPUT88), .Z(n655) );
  XNOR2_X1 U729 ( .A(n656), .B(n655), .ZN(n657) );
  NAND2_X1 U730 ( .A1(n657), .A2(G2090), .ZN(n658) );
  XOR2_X1 U731 ( .A(KEYINPUT21), .B(n658), .Z(n659) );
  XNOR2_X1 U732 ( .A(KEYINPUT89), .B(n659), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n660), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U734 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U735 ( .A1(G220), .A2(G219), .ZN(n661) );
  XOR2_X1 U736 ( .A(KEYINPUT22), .B(n661), .Z(n662) );
  NOR2_X1 U737 ( .A1(G218), .A2(n662), .ZN(n663) );
  NAND2_X1 U738 ( .A1(G96), .A2(n663), .ZN(n826) );
  NAND2_X1 U739 ( .A1(n826), .A2(G2106), .ZN(n667) );
  NAND2_X1 U740 ( .A1(G69), .A2(G120), .ZN(n664) );
  NOR2_X1 U741 ( .A1(G237), .A2(n664), .ZN(n665) );
  NAND2_X1 U742 ( .A1(G108), .A2(n665), .ZN(n825) );
  NAND2_X1 U743 ( .A1(n825), .A2(G567), .ZN(n666) );
  NAND2_X1 U744 ( .A1(n667), .A2(n666), .ZN(n909) );
  NAND2_X1 U745 ( .A1(G483), .A2(G661), .ZN(n668) );
  NOR2_X1 U746 ( .A1(n909), .A2(n668), .ZN(n824) );
  NAND2_X1 U747 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U748 ( .A1(G126), .A2(n880), .ZN(n670) );
  NAND2_X1 U749 ( .A1(G138), .A2(n876), .ZN(n669) );
  NAND2_X1 U750 ( .A1(n670), .A2(n669), .ZN(n674) );
  NAND2_X1 U751 ( .A1(G114), .A2(n881), .ZN(n672) );
  NAND2_X1 U752 ( .A1(G102), .A2(n877), .ZN(n671) );
  NAND2_X1 U753 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U754 ( .A1(n674), .A2(n673), .ZN(G164) );
  XOR2_X1 U755 ( .A(KEYINPUT90), .B(G166), .Z(G303) );
  NAND2_X1 U756 ( .A1(G160), .A2(G40), .ZN(n768) );
  INV_X1 U757 ( .A(n768), .ZN(n675) );
  NOR2_X1 U758 ( .A1(G164), .A2(G1384), .ZN(n769) );
  NAND2_X1 U759 ( .A1(n675), .A2(n769), .ZN(n676) );
  NAND2_X1 U760 ( .A1(G8), .A2(n720), .ZN(n762) );
  AND2_X1 U761 ( .A1(n704), .A2(G1996), .ZN(n677) );
  XNOR2_X1 U762 ( .A(n677), .B(KEYINPUT26), .ZN(n679) );
  AND2_X1 U763 ( .A1(n720), .A2(G1341), .ZN(n678) );
  OR2_X1 U764 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U765 ( .A1(n680), .A2(n1002), .ZN(n686) );
  NAND2_X1 U766 ( .A1(n686), .A2(n989), .ZN(n685) );
  AND2_X1 U767 ( .A1(n720), .A2(G1348), .ZN(n681) );
  XNOR2_X1 U768 ( .A(n681), .B(KEYINPUT103), .ZN(n683) );
  NAND2_X1 U769 ( .A1(n704), .A2(G2067), .ZN(n682) );
  NAND2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U771 ( .A1(n685), .A2(n684), .ZN(n688) );
  OR2_X1 U772 ( .A1(n989), .A2(n686), .ZN(n687) );
  NAND2_X1 U773 ( .A1(n688), .A2(n687), .ZN(n696) );
  NAND2_X1 U774 ( .A1(G2072), .A2(n704), .ZN(n689) );
  XNOR2_X1 U775 ( .A(KEYINPUT101), .B(n689), .ZN(n691) );
  INV_X1 U776 ( .A(KEYINPUT27), .ZN(n690) );
  XNOR2_X1 U777 ( .A(n691), .B(n690), .ZN(n694) );
  NAND2_X1 U778 ( .A1(G1956), .A2(n720), .ZN(n692) );
  XOR2_X1 U779 ( .A(KEYINPUT102), .B(n692), .Z(n693) );
  NOR2_X1 U780 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U781 ( .A1(n1001), .A2(n697), .ZN(n695) );
  NAND2_X1 U782 ( .A1(n696), .A2(n695), .ZN(n701) );
  NOR2_X1 U783 ( .A1(n697), .A2(n1001), .ZN(n699) );
  INV_X1 U784 ( .A(KEYINPUT28), .ZN(n698) );
  XNOR2_X1 U785 ( .A(n699), .B(n698), .ZN(n700) );
  NAND2_X1 U786 ( .A1(n701), .A2(n700), .ZN(n703) );
  OR2_X1 U787 ( .A1(n704), .A2(G1961), .ZN(n706) );
  XNOR2_X1 U788 ( .A(G2078), .B(KEYINPUT25), .ZN(n912) );
  NAND2_X1 U789 ( .A1(n704), .A2(n912), .ZN(n705) );
  NAND2_X1 U790 ( .A1(n706), .A2(n705), .ZN(n710) );
  AND2_X1 U791 ( .A1(n710), .A2(G171), .ZN(n707) );
  XOR2_X1 U792 ( .A(KEYINPUT100), .B(n707), .Z(n708) );
  NAND2_X1 U793 ( .A1(n709), .A2(n708), .ZN(n718) );
  NOR2_X1 U794 ( .A1(G171), .A2(n710), .ZN(n715) );
  NOR2_X1 U795 ( .A1(G1966), .A2(n762), .ZN(n730) );
  NOR2_X1 U796 ( .A1(G2084), .A2(n720), .ZN(n733) );
  NOR2_X1 U797 ( .A1(n730), .A2(n733), .ZN(n711) );
  NAND2_X1 U798 ( .A1(G8), .A2(n711), .ZN(n712) );
  XNOR2_X1 U799 ( .A(KEYINPUT30), .B(n712), .ZN(n713) );
  NOR2_X1 U800 ( .A1(G168), .A2(n713), .ZN(n714) );
  NOR2_X1 U801 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U802 ( .A(KEYINPUT31), .B(n716), .Z(n717) );
  NAND2_X1 U803 ( .A1(n718), .A2(n717), .ZN(n729) );
  NAND2_X1 U804 ( .A1(n729), .A2(G286), .ZN(n725) );
  NOR2_X1 U805 ( .A1(G1971), .A2(n762), .ZN(n719) );
  XOR2_X1 U806 ( .A(KEYINPUT105), .B(n719), .Z(n722) );
  NOR2_X1 U807 ( .A1(G2090), .A2(n720), .ZN(n721) );
  NOR2_X1 U808 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U809 ( .A1(G303), .A2(n723), .ZN(n724) );
  NAND2_X1 U810 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U811 ( .A1(n726), .A2(G8), .ZN(n727) );
  XNOR2_X1 U812 ( .A(n727), .B(KEYINPUT32), .ZN(n728) );
  XNOR2_X1 U813 ( .A(KEYINPUT106), .B(n728), .ZN(n747) );
  INV_X1 U814 ( .A(n729), .ZN(n731) );
  XNOR2_X1 U815 ( .A(n732), .B(KEYINPUT104), .ZN(n735) );
  NAND2_X1 U816 ( .A1(n733), .A2(G8), .ZN(n734) );
  NAND2_X1 U817 ( .A1(n735), .A2(n734), .ZN(n745) );
  NAND2_X1 U818 ( .A1(n747), .A2(n745), .ZN(n738) );
  NOR2_X1 U819 ( .A1(G2090), .A2(G303), .ZN(n736) );
  NAND2_X1 U820 ( .A1(G8), .A2(n736), .ZN(n737) );
  NAND2_X1 U821 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U822 ( .A1(n762), .A2(n739), .ZN(n766) );
  NAND2_X1 U823 ( .A1(G1976), .A2(G288), .ZN(n994) );
  XOR2_X1 U824 ( .A(G1981), .B(G305), .Z(n1005) );
  NOR2_X1 U825 ( .A1(G288), .A2(G1976), .ZN(n740) );
  XNOR2_X1 U826 ( .A(n740), .B(KEYINPUT107), .ZN(n748) );
  NOR2_X1 U827 ( .A1(n762), .A2(n748), .ZN(n741) );
  NAND2_X1 U828 ( .A1(KEYINPUT33), .A2(n741), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n1005), .A2(n742), .ZN(n755) );
  INV_X1 U830 ( .A(n755), .ZN(n743) );
  AND2_X1 U831 ( .A1(n994), .A2(n743), .ZN(n744) );
  AND2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n757) );
  INV_X1 U834 ( .A(n994), .ZN(n751) );
  INV_X1 U835 ( .A(n748), .ZN(n750) );
  NOR2_X1 U836 ( .A1(G303), .A2(G1971), .ZN(n749) );
  NOR2_X1 U837 ( .A1(n750), .A2(n749), .ZN(n995) );
  OR2_X1 U838 ( .A1(n751), .A2(n995), .ZN(n752) );
  NOR2_X1 U839 ( .A1(n762), .A2(n752), .ZN(n753) );
  NOR2_X1 U840 ( .A1(KEYINPUT33), .A2(n753), .ZN(n754) );
  OR2_X1 U841 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U842 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U843 ( .A(n758), .B(KEYINPUT108), .ZN(n764) );
  NOR2_X1 U844 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XNOR2_X1 U845 ( .A(n759), .B(KEYINPUT24), .ZN(n760) );
  XNOR2_X1 U846 ( .A(n760), .B(KEYINPUT99), .ZN(n761) );
  NOR2_X1 U847 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U848 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U849 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U850 ( .A(n767), .B(KEYINPUT109), .ZN(n802) );
  NOR2_X1 U851 ( .A1(n769), .A2(n768), .ZN(n816) );
  NAND2_X1 U852 ( .A1(G119), .A2(n880), .ZN(n771) );
  NAND2_X1 U853 ( .A1(G107), .A2(n881), .ZN(n770) );
  NAND2_X1 U854 ( .A1(n771), .A2(n770), .ZN(n776) );
  NAND2_X1 U855 ( .A1(G131), .A2(n876), .ZN(n773) );
  NAND2_X1 U856 ( .A1(G95), .A2(n877), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U858 ( .A(KEYINPUT93), .B(n774), .Z(n775) );
  NOR2_X1 U859 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U860 ( .A(KEYINPUT94), .B(n777), .Z(n890) );
  NAND2_X1 U861 ( .A1(G1991), .A2(n890), .ZN(n778) );
  XOR2_X1 U862 ( .A(KEYINPUT95), .B(n778), .Z(n788) );
  XOR2_X1 U863 ( .A(KEYINPUT38), .B(KEYINPUT96), .Z(n780) );
  NAND2_X1 U864 ( .A1(G105), .A2(n877), .ZN(n779) );
  XNOR2_X1 U865 ( .A(n780), .B(n779), .ZN(n784) );
  NAND2_X1 U866 ( .A1(G129), .A2(n880), .ZN(n782) );
  NAND2_X1 U867 ( .A1(G141), .A2(n876), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U869 ( .A1(n784), .A2(n783), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n881), .A2(G117), .ZN(n785) );
  NAND2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n874) );
  NAND2_X1 U872 ( .A1(G1996), .A2(n874), .ZN(n787) );
  NAND2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n974) );
  NAND2_X1 U874 ( .A1(n816), .A2(n974), .ZN(n789) );
  XNOR2_X1 U875 ( .A(KEYINPUT97), .B(n789), .ZN(n809) );
  XOR2_X1 U876 ( .A(KEYINPUT98), .B(n809), .Z(n800) );
  NAND2_X1 U877 ( .A1(G140), .A2(n876), .ZN(n791) );
  NAND2_X1 U878 ( .A1(G104), .A2(n877), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U880 ( .A(KEYINPUT34), .B(n792), .ZN(n798) );
  NAND2_X1 U881 ( .A1(n880), .A2(G128), .ZN(n793) );
  XNOR2_X1 U882 ( .A(n793), .B(KEYINPUT92), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G116), .A2(n881), .ZN(n794) );
  NAND2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U885 ( .A(KEYINPUT35), .B(n796), .Z(n797) );
  NOR2_X1 U886 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U887 ( .A(KEYINPUT36), .B(n799), .ZN(n895) );
  XNOR2_X1 U888 ( .A(KEYINPUT37), .B(G2067), .ZN(n814) );
  NOR2_X1 U889 ( .A1(n895), .A2(n814), .ZN(n961) );
  NAND2_X1 U890 ( .A1(n816), .A2(n961), .ZN(n812) );
  NAND2_X1 U891 ( .A1(n800), .A2(n812), .ZN(n801) );
  NOR2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n805) );
  XOR2_X1 U893 ( .A(G1986), .B(KEYINPUT91), .Z(n803) );
  XNOR2_X1 U894 ( .A(G290), .B(n803), .ZN(n993) );
  NAND2_X1 U895 ( .A1(n993), .A2(n816), .ZN(n804) );
  NAND2_X1 U896 ( .A1(n805), .A2(n804), .ZN(n819) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n874), .ZN(n967) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n890), .ZN(n970) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n806) );
  XNOR2_X1 U900 ( .A(KEYINPUT110), .B(n806), .ZN(n807) );
  NOR2_X1 U901 ( .A1(n970), .A2(n807), .ZN(n808) );
  NOR2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U903 ( .A1(n967), .A2(n810), .ZN(n811) );
  XNOR2_X1 U904 ( .A(n811), .B(KEYINPUT39), .ZN(n813) );
  NAND2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n815) );
  NAND2_X1 U906 ( .A1(n895), .A2(n814), .ZN(n960) );
  NAND2_X1 U907 ( .A1(n815), .A2(n960), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(n820), .ZN(G329) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U913 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(G188) );
  INV_X1 U917 ( .A(G120), .ZN(G236) );
  INV_X1 U918 ( .A(G96), .ZN(G221) );
  INV_X1 U919 ( .A(G69), .ZN(G235) );
  NOR2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U921 ( .A(n827), .B(KEYINPUT115), .ZN(G261) );
  INV_X1 U922 ( .A(G261), .ZN(G325) );
  XOR2_X1 U923 ( .A(G2438), .B(KEYINPUT112), .Z(n829) );
  XNOR2_X1 U924 ( .A(G2454), .B(G2435), .ZN(n828) );
  XNOR2_X1 U925 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U926 ( .A(n830), .B(G2430), .Z(n832) );
  XNOR2_X1 U927 ( .A(G1341), .B(G1348), .ZN(n831) );
  XNOR2_X1 U928 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U929 ( .A(G2427), .B(KEYINPUT113), .Z(n834) );
  XNOR2_X1 U930 ( .A(G2443), .B(G2446), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U932 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U933 ( .A(KEYINPUT111), .B(G2451), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(n839) );
  NAND2_X1 U935 ( .A1(G14), .A2(n839), .ZN(n840) );
  XOR2_X1 U936 ( .A(KEYINPUT114), .B(n840), .Z(G401) );
  XOR2_X1 U937 ( .A(KEYINPUT41), .B(G1961), .Z(n842) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U940 ( .A(n843), .B(KEYINPUT116), .Z(n845) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1976), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U943 ( .A(G1981), .B(G1966), .Z(n847) );
  XNOR2_X1 U944 ( .A(G1971), .B(G1956), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U946 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U947 ( .A(KEYINPUT117), .B(G2474), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(G229) );
  XOR2_X1 U949 ( .A(G2096), .B(G2100), .Z(n853) );
  XNOR2_X1 U950 ( .A(KEYINPUT42), .B(G2678), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U952 ( .A(KEYINPUT43), .B(G2072), .Z(n855) );
  XNOR2_X1 U953 ( .A(G2067), .B(G2090), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U956 ( .A(G2078), .B(G2084), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(G227) );
  NAND2_X1 U958 ( .A1(G136), .A2(n876), .ZN(n861) );
  NAND2_X1 U959 ( .A1(G112), .A2(n881), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n866) );
  NAND2_X1 U961 ( .A1(n880), .A2(G124), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G100), .A2(n877), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U965 ( .A1(n866), .A2(n865), .ZN(G162) );
  NAND2_X1 U966 ( .A1(G130), .A2(n880), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G118), .A2(n881), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n873) );
  NAND2_X1 U969 ( .A1(G142), .A2(n876), .ZN(n870) );
  NAND2_X1 U970 ( .A1(G106), .A2(n877), .ZN(n869) );
  NAND2_X1 U971 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U972 ( .A(n871), .B(KEYINPUT45), .Z(n872) );
  NOR2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(n894) );
  XOR2_X1 U975 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n888) );
  NAND2_X1 U976 ( .A1(G139), .A2(n876), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G103), .A2(n877), .ZN(n878) );
  NAND2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n886) );
  NAND2_X1 U979 ( .A1(G127), .A2(n880), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G115), .A2(n881), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n884), .Z(n885) );
  NOR2_X1 U983 ( .A1(n886), .A2(n885), .ZN(n977) );
  XNOR2_X1 U984 ( .A(G164), .B(n977), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U986 ( .A(n889), .B(G162), .Z(n892) );
  XNOR2_X1 U987 ( .A(G160), .B(n890), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n897) );
  XNOR2_X1 U990 ( .A(n895), .B(n965), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(G395) );
  XNOR2_X1 U993 ( .A(n1002), .B(n899), .ZN(n901) );
  XNOR2_X1 U994 ( .A(G286), .B(n989), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U996 ( .A(G171), .B(n902), .ZN(n903) );
  NOR2_X1 U997 ( .A1(G37), .A2(n903), .ZN(G397) );
  OR2_X1 U998 ( .A1(n909), .A2(G401), .ZN(n906) );
  NOR2_X1 U999 ( .A1(G229), .A2(G227), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(KEYINPUT49), .B(n904), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(n906), .A2(n905), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n907) );
  NAND2_X1 U1003 ( .A1(n908), .A2(n907), .ZN(G225) );
  INV_X1 U1004 ( .A(G225), .ZN(G308) );
  INV_X1 U1005 ( .A(n909), .ZN(G319) );
  INV_X1 U1006 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1007 ( .A(KEYINPUT119), .B(G1996), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(n910), .B(G32), .ZN(n920) );
  XOR2_X1 U1009 ( .A(G2072), .B(G33), .Z(n911) );
  NAND2_X1 U1010 ( .A1(n911), .A2(G28), .ZN(n918) );
  XNOR2_X1 U1011 ( .A(G27), .B(n912), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(G2067), .B(G26), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(G1991), .B(G25), .ZN(n913) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1015 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  XNOR2_X1 U1018 ( .A(n921), .B(KEYINPUT53), .ZN(n924) );
  XOR2_X1 U1019 ( .A(G2084), .B(G34), .Z(n922) );
  XNOR2_X1 U1020 ( .A(KEYINPUT54), .B(n922), .ZN(n923) );
  NAND2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(G35), .B(G2090), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(KEYINPUT55), .B(n927), .ZN(n929) );
  INV_X1 U1025 ( .A(G29), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n930), .A2(G11), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(n931), .B(KEYINPUT120), .ZN(n959) );
  XOR2_X1 U1029 ( .A(G1986), .B(G24), .Z(n933) );
  XOR2_X1 U1030 ( .A(G1971), .B(G22), .Z(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(G23), .B(G1976), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(KEYINPUT58), .B(n936), .ZN(n955) );
  XNOR2_X1 U1035 ( .A(G1961), .B(G5), .ZN(n952) );
  XNOR2_X1 U1036 ( .A(G1341), .B(G19), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(G6), .B(G1981), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1039 ( .A(KEYINPUT123), .B(n939), .Z(n943) );
  XNOR2_X1 U1040 ( .A(KEYINPUT59), .B(KEYINPUT124), .ZN(n940) );
  XNOR2_X1 U1041 ( .A(n940), .B(G4), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(G1348), .B(n941), .ZN(n942) );
  NAND2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(KEYINPUT122), .B(G1956), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(G20), .B(n944), .ZN(n945) );
  NOR2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1047 ( .A(KEYINPUT60), .B(n947), .Z(n949) );
  XNOR2_X1 U1048 ( .A(G1966), .B(G21), .ZN(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(KEYINPUT125), .B(n950), .ZN(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1052 ( .A(KEYINPUT126), .B(n953), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1054 ( .A(KEYINPUT61), .B(n956), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n957), .A2(G16), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n988) );
  INV_X1 U1057 ( .A(n960), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n976) );
  XOR2_X1 U1059 ( .A(G2084), .B(G160), .Z(n963) );
  XNOR2_X1 U1060 ( .A(KEYINPUT118), .B(n963), .ZN(n964) );
  NOR2_X1 U1061 ( .A1(n965), .A2(n964), .ZN(n972) );
  XOR2_X1 U1062 ( .A(G2090), .B(G162), .Z(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(n968), .B(KEYINPUT51), .ZN(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n982) );
  XOR2_X1 U1069 ( .A(G2072), .B(n977), .Z(n979) );
  XOR2_X1 U1070 ( .A(G164), .B(G2078), .Z(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1072 ( .A(KEYINPUT50), .B(n980), .Z(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(KEYINPUT52), .B(n983), .ZN(n985) );
  INV_X1 U1075 ( .A(KEYINPUT55), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n986), .A2(G29), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n1015) );
  XOR2_X1 U1079 ( .A(KEYINPUT56), .B(G16), .Z(n1013) );
  XNOR2_X1 U1080 ( .A(G171), .B(G1961), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(n989), .B(G1348), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n1000) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n997) );
  AND2_X1 U1085 ( .A1(G303), .A2(G1971), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1087 ( .A(KEYINPUT121), .B(n998), .Z(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1011) );
  XOR2_X1 U1089 ( .A(n1001), .B(G1956), .Z(n1004) );
  XNOR2_X1 U1090 ( .A(n1002), .B(G1341), .ZN(n1003) );
  NOR2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(G168), .B(G1966), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(n1007), .B(KEYINPUT57), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1097 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1098 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1099 ( .A(n1016), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1100 ( .A(G311), .ZN(G150) );
endmodule

