//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n586, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT70), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(KEYINPUT70), .A3(new_n464), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n469), .A2(new_n470), .B1(G113), .B2(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(KEYINPUT69), .A3(G125), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n460), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(new_n474), .ZN(G160));
  INV_X1    g050(.A(new_n461), .ZN(new_n476));
  INV_X1    g051(.A(new_n462), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n460), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(G136), .B2(new_n483), .ZN(G162));
  INV_X1    g059(.A(G138), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n486), .B1(new_n461), .B2(new_n462), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n486), .B(new_n489), .C1(new_n462), .C2(new_n461), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n491), .A2(new_n498), .A3(KEYINPUT71), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT71), .B1(new_n491), .B2(new_n498), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  OR2_X1    g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n503), .A2(new_n507), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  XOR2_X1   g093(.A(new_n518), .B(KEYINPUT73), .Z(new_n519));
  NAND2_X1  g094(.A1(new_n513), .A2(G62), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n516), .A2(new_n521), .ZN(G166));
  INV_X1    g097(.A(new_n514), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n525), .B(new_n527), .C1(new_n507), .C2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n524), .A2(new_n529), .ZN(G168));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n510), .A2(new_n512), .ZN(new_n532));
  INV_X1    g107(.A(G64), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n517), .B1(new_n534), .B2(KEYINPUT74), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n535), .B1(KEYINPUT74), .B2(new_n534), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n504), .A2(new_n505), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n508), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n523), .A2(G90), .B1(G52), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n523), .A2(G81), .B1(G43), .B2(new_n538), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n517), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(new_n547));
  XOR2_X1   g122(.A(new_n547), .B(KEYINPUT75), .Z(G153));
  NAND4_X1  g123(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  AOI22_X1  g127(.A1(new_n513), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n517), .ZN(new_n554));
  OAI211_X1 g129(.A(G53), .B(G543), .C1(new_n504), .C2(new_n505), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n523), .A2(G91), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(G299));
  INV_X1    g133(.A(G168), .ZN(G286));
  INV_X1    g134(.A(G166), .ZN(G303));
  AOI22_X1  g135(.A1(new_n523), .A2(G87), .B1(G49), .B2(new_n538), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(G288));
  INV_X1    g138(.A(G48), .ZN(new_n564));
  INV_X1    g139(.A(G86), .ZN(new_n565));
  OAI22_X1  g140(.A1(new_n564), .A2(new_n507), .B1(new_n514), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n517), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n566), .A2(new_n568), .ZN(G305));
  AOI22_X1  g144(.A1(new_n523), .A2(G85), .B1(G47), .B2(new_n538), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n517), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(G290));
  NAND3_X1  g148(.A1(new_n506), .A2(new_n513), .A3(G92), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT10), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G79), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G66), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n532), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(G54), .B2(new_n538), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G868), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(G171), .B2(new_n582), .ZN(G284));
  OAI21_X1  g159(.A(new_n583), .B1(G171), .B2(new_n582), .ZN(G321));
  NAND2_X1  g160(.A1(G299), .A2(new_n582), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n586), .B1(new_n582), .B2(G168), .ZN(G297));
  OAI21_X1  g162(.A(new_n586), .B1(new_n582), .B2(G168), .ZN(G280));
  AND2_X1   g163(.A1(new_n576), .A2(new_n580), .ZN(new_n589));
  XNOR2_X1  g164(.A(KEYINPUT76), .B(G559), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(G860), .B2(new_n590), .ZN(G148));
  NAND2_X1  g166(.A1(new_n545), .A2(new_n582), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n589), .A2(new_n590), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n592), .B1(new_n594), .B2(new_n582), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT77), .ZN(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XOR2_X1   g172(.A(KEYINPUT78), .B(KEYINPUT12), .Z(new_n598));
  NAND3_X1  g173(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT13), .ZN(new_n601));
  XNOR2_X1  g176(.A(KEYINPUT79), .B(G2100), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n478), .A2(G123), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT80), .ZN(new_n605));
  OR3_X1    g180(.A1(new_n460), .A2(KEYINPUT81), .A3(G111), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT81), .B1(new_n460), .B2(G111), .ZN(new_n607));
  OR2_X1    g182(.A1(G99), .A2(G2105), .ZN(new_n608));
  AND3_X1   g183(.A1(new_n607), .A2(G2104), .A3(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n606), .A2(new_n609), .B1(new_n483), .B2(G135), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(G2096), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n601), .A2(new_n602), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n611), .A2(G2096), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n603), .A2(new_n612), .A3(new_n613), .A4(new_n614), .ZN(G156));
  XNOR2_X1  g190(.A(G2427), .B(G2438), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2430), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT15), .B(G2435), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n619), .A2(KEYINPUT14), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT83), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2451), .B(G2454), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2443), .B(G2446), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n622), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(new_n631), .A3(G14), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(G401));
  INV_X1    g208(.A(KEYINPUT18), .ZN(new_n634));
  XOR2_X1   g209(.A(G2084), .B(G2090), .Z(new_n635));
  XNOR2_X1  g210(.A(G2067), .B(G2678), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT17), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n635), .A2(new_n636), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n637), .B2(KEYINPUT18), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2096), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(G227));
  XNOR2_X1  g220(.A(G1971), .B(G1976), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1956), .B(G2474), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1961), .B(G1966), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n649), .A2(new_n650), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n648), .A2(new_n657), .ZN(new_n658));
  OR3_X1    g233(.A1(new_n648), .A2(new_n651), .A3(new_n657), .ZN(new_n659));
  NAND4_X1  g234(.A1(new_n654), .A2(new_n655), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1991), .B(G1996), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G1981), .B(G1986), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G229));
  NOR2_X1   g241(.A1(G6), .A2(G16), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n566), .A2(new_n568), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n667), .B1(new_n668), .B2(G16), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT32), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1981), .ZN(new_n671));
  OR2_X1    g246(.A1(G16), .A2(G23), .ZN(new_n672));
  NAND2_X1  g247(.A1(G288), .A2(KEYINPUT89), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT89), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n561), .A2(new_n674), .A3(new_n562), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT33), .B(G1976), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT87), .B(G16), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n683), .A2(G22), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G166), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1971), .ZN(new_n686));
  NOR4_X1   g261(.A1(new_n671), .A2(new_n680), .A3(new_n681), .A4(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n683), .A2(G24), .ZN(new_n691));
  INV_X1    g266(.A(G290), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n683), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT88), .Z(new_n694));
  INV_X1    g269(.A(G1986), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n483), .A2(G131), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n478), .A2(G119), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n460), .A2(G107), .ZN(new_n700));
  OAI21_X1  g275(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n698), .B(new_n699), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G25), .B(new_n702), .S(G29), .Z(new_n703));
  XOR2_X1   g278(.A(KEYINPUT35), .B(G1991), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT86), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n696), .A2(new_n697), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n689), .A2(new_n690), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT36), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n683), .A2(G19), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n546), .B2(new_n683), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1341), .ZN(new_n712));
  NOR2_X1   g287(.A1(G4), .A2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT90), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n581), .B2(new_n677), .ZN(new_n715));
  INV_X1    g290(.A(G1348), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G29), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G26), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n483), .A2(G140), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n478), .A2(G128), .ZN(new_n722));
  OR2_X1    g297(.A1(G104), .A2(G2105), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n723), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n720), .B1(new_n726), .B2(new_n718), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G2067), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n712), .A2(new_n717), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  NOR2_X1   g305(.A1(G27), .A2(G29), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G164), .B2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2078), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n682), .A2(G20), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT23), .Z(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G299), .B2(G16), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1956), .ZN(new_n737));
  INV_X1    g312(.A(G1961), .ZN(new_n738));
  NOR2_X1   g313(.A1(G5), .A2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT94), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G301), .B2(new_n677), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n737), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  AOI211_X1 g317(.A(new_n733), .B(new_n742), .C1(new_n738), .C2(new_n741), .ZN(new_n743));
  NOR2_X1   g318(.A1(G29), .A2(G35), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G162), .B2(G29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT29), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2090), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n718), .A2(G32), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n483), .A2(G141), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT93), .ZN(new_n750));
  AND3_X1   g325(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT26), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n751), .B(new_n753), .C1(G129), .C2(new_n478), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n748), .B1(new_n755), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(G2072), .ZN(new_n759));
  OR2_X1    g334(.A1(G29), .A2(G33), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n483), .A2(G139), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT92), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT25), .Z(new_n764));
  AOI22_X1  g339(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n762), .B(new_n764), .C1(new_n460), .C2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n760), .B1(new_n766), .B2(new_n718), .ZN(new_n767));
  INV_X1    g342(.A(G1966), .ZN(new_n768));
  NOR2_X1   g343(.A1(G168), .A2(new_n677), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n677), .B2(G21), .ZN(new_n770));
  OAI221_X1 g345(.A(new_n758), .B1(new_n759), .B2(new_n767), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT31), .B(G11), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT30), .B(G28), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(new_n718), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n772), .B(new_n774), .C1(new_n611), .C2(new_n718), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n770), .B2(new_n768), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n767), .A2(new_n759), .B1(new_n756), .B2(new_n757), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AND2_X1   g353(.A1(KEYINPUT24), .A2(G34), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n718), .B1(KEYINPUT24), .B2(G34), .ZN(new_n780));
  OAI22_X1  g355(.A1(G160), .A2(new_n718), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2084), .ZN(new_n782));
  NOR4_X1   g357(.A1(new_n747), .A2(new_n771), .A3(new_n778), .A4(new_n782), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n730), .A2(new_n743), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n709), .A2(new_n784), .ZN(G150));
  INV_X1    g360(.A(G150), .ZN(G311));
  AOI22_X1  g361(.A1(new_n523), .A2(G93), .B1(G55), .B2(new_n538), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(new_n517), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G860), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n787), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n794), .B1(new_n787), .B2(new_n789), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n545), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n790), .A2(KEYINPUT95), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n799), .A2(new_n546), .A3(new_n795), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n589), .A2(G559), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT96), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(KEYINPUT38), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n803), .A2(KEYINPUT38), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n801), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n803), .A2(KEYINPUT38), .ZN(new_n808));
  INV_X1    g383(.A(new_n801), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n808), .A2(new_n809), .A3(new_n804), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT39), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(KEYINPUT97), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT97), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n811), .A2(new_n815), .A3(new_n812), .ZN(new_n816));
  AOI21_X1  g391(.A(G860), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n807), .A2(KEYINPUT39), .A3(new_n810), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT98), .Z(new_n819));
  AND3_X1   g394(.A1(new_n817), .A2(new_n819), .A3(KEYINPUT99), .ZN(new_n820));
  AOI21_X1  g395(.A(KEYINPUT99), .B1(new_n817), .B2(new_n819), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n793), .B1(new_n820), .B2(new_n821), .ZN(G145));
  NAND2_X1  g397(.A1(new_n766), .A2(KEYINPUT104), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n755), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n702), .B(new_n600), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT103), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n497), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n492), .A2(KEYINPUT103), .A3(new_n496), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n828), .A2(new_n829), .B1(new_n488), .B2(new_n490), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(new_n726), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n478), .A2(G130), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n460), .A2(G118), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G142), .B2(new_n483), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n831), .B(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n826), .B(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n611), .B(G162), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(G160), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT101), .B(KEYINPUT102), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(G37), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n842), .B2(new_n838), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g420(.A(KEYINPUT108), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n692), .A2(G303), .ZN(new_n847));
  NAND2_X1  g422(.A1(G290), .A2(G166), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n673), .A2(G305), .A3(new_n675), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(G305), .B1(new_n673), .B2(new_n675), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n676), .A2(new_n668), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n854), .A2(new_n850), .A3(new_n848), .A4(new_n847), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n846), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  AOI211_X1 g434(.A(KEYINPUT108), .B(new_n857), .C1(new_n853), .C2(new_n855), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n801), .A2(new_n594), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n798), .A2(new_n593), .A3(new_n800), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n581), .A2(new_n556), .A3(new_n554), .A4(new_n557), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n866));
  NAND3_X1  g441(.A1(G299), .A2(new_n576), .A3(new_n580), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n589), .A2(KEYINPUT105), .A3(G299), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n868), .A2(KEYINPUT106), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT106), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n864), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n868), .A2(KEYINPUT41), .A3(new_n869), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n865), .A2(new_n874), .A3(new_n867), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n876), .A2(new_n862), .A3(new_n863), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n861), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n877), .B(new_n872), .C1(new_n859), .C2(new_n860), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n879), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(G868), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n790), .A2(new_n582), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(G295));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n884), .A2(new_n887), .A3(new_n885), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n887), .B1(new_n884), .B2(new_n885), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(G331));
  INV_X1    g465(.A(new_n876), .ZN(new_n891));
  AOI21_X1  g466(.A(G168), .B1(new_n536), .B2(new_n539), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n536), .A2(G168), .A3(new_n539), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n796), .A2(new_n545), .A3(new_n797), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n546), .B1(new_n799), .B2(new_n795), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n893), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n894), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n798), .B(new_n800), .C1(new_n898), .C2(new_n892), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT110), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(KEYINPUT110), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n891), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n897), .A2(new_n899), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n868), .A2(new_n869), .ZN(new_n905));
  OR2_X1    g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n856), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n856), .B1(new_n903), .B2(new_n906), .ZN(new_n910));
  OR3_X1    g485(.A1(new_n909), .A2(KEYINPUT43), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  INV_X1    g487(.A(new_n856), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n870), .A2(new_n871), .ZN(new_n914));
  INV_X1    g489(.A(new_n904), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n914), .B(new_n901), .C1(new_n915), .C2(KEYINPUT110), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n905), .A2(new_n874), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n865), .A2(new_n867), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT41), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n904), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n904), .A2(KEYINPUT111), .A3(new_n917), .A4(new_n919), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n916), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n909), .B1(new_n913), .B2(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n911), .B(KEYINPUT44), .C1(new_n912), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n913), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n927), .A2(new_n912), .A3(new_n908), .A4(new_n907), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n909), .B2(new_n910), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT112), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT112), .ZN(new_n933));
  AOI211_X1 g508(.A(new_n933), .B(KEYINPUT44), .C1(new_n928), .C2(new_n929), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n926), .B1(new_n932), .B2(new_n934), .ZN(G397));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n830), .B2(G1384), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n471), .A2(new_n473), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(G2105), .ZN(new_n939));
  INV_X1    g514(.A(new_n467), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(new_n465), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n941), .A3(G40), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n937), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G1996), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT46), .ZN(new_n946));
  INV_X1    g521(.A(G2067), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n725), .B(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n943), .B1(new_n949), .B2(new_n755), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT47), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n755), .A2(G1996), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n750), .A2(new_n944), .A3(new_n754), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n954), .A3(new_n948), .ZN(new_n955));
  INV_X1    g530(.A(new_n704), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n702), .A2(new_n956), .ZN(new_n957));
  OAI22_X1  g532(.A1(new_n955), .A2(new_n957), .B1(G2067), .B2(new_n725), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n943), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n702), .B(new_n956), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n955), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n943), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT48), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n943), .A2(new_n695), .A3(new_n692), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n966), .B1(new_n964), .B2(new_n965), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n952), .A2(new_n959), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT118), .ZN(new_n969));
  INV_X1    g544(.A(G8), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT55), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n970), .B1(KEYINPUT114), .B2(new_n971), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n971), .A2(KEYINPUT114), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT115), .Z(new_n974));
  AND3_X1   g549(.A1(G303), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(G303), .B2(new_n972), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n828), .A2(new_n829), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n980), .B2(new_n491), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n942), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT71), .ZN(new_n983));
  INV_X1    g558(.A(new_n490), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n489), .B1(new_n472), .B2(new_n486), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n983), .B1(new_n986), .B2(new_n497), .ZN(new_n987));
  INV_X1    g562(.A(G1384), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n491), .A2(new_n498), .A3(KEYINPUT71), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT50), .ZN(new_n991));
  INV_X1    g566(.A(G2090), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n982), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n936), .A2(G1384), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n980), .B2(new_n491), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n996), .B(new_n942), .C1(new_n990), .C2(new_n936), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n993), .B(KEYINPUT113), .C1(new_n997), .C2(G1971), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(G8), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n996), .B1(new_n990), .B2(new_n936), .ZN(new_n1000));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n468), .A2(new_n474), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1971), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT113), .B1(new_n1005), .B2(new_n993), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n978), .B1(new_n999), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n987), .A2(new_n989), .A3(new_n994), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n937), .A2(new_n1008), .A3(new_n1002), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT117), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(new_n768), .ZN(new_n1011));
  INV_X1    g586(.A(G2084), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n982), .A2(new_n991), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1010), .B1(new_n1009), .B2(new_n768), .ZN(new_n1015));
  OAI211_X1 g590(.A(G8), .B(G168), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT63), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1007), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n982), .A2(new_n992), .A3(new_n991), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1971), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1023), .A2(G8), .A3(new_n977), .A4(new_n998), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G305), .A2(G1981), .ZN(new_n1025));
  INV_X1    g600(.A(G1981), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n668), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(KEYINPUT49), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n970), .B1(new_n1002), .B2(new_n981), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1025), .B(new_n1027), .C1(new_n1029), .C2(KEYINPUT49), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1976), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1032), .B1(new_n676), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT52), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(G288), .B2(new_n1035), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1032), .B(new_n1038), .C1(new_n676), .C2(new_n1035), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1034), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1024), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n969), .B1(new_n1019), .B2(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1024), .A2(new_n1040), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1043), .A2(KEYINPUT118), .A3(new_n1007), .A4(new_n1018), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT50), .B1(new_n830), .B2(G1384), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1045), .B(new_n1002), .C1(new_n990), .C2(KEYINPUT50), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(G2090), .ZN(new_n1047));
  OAI21_X1  g622(.A(G8), .B1(new_n1022), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n978), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1024), .A2(new_n1049), .A3(new_n1040), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1017), .B1(new_n1050), .B2(new_n1016), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1042), .A2(new_n1044), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G286), .A2(G8), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT124), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1053), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT51), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1009), .A2(new_n768), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT117), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1062), .A2(new_n1013), .A3(new_n1011), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1056), .B1(new_n1063), .B2(G8), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1058), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT62), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT126), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n942), .B1(new_n501), .B2(new_n994), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT125), .ZN(new_n1070));
  INV_X1    g645(.A(G2078), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .A4(new_n937), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n937), .A2(new_n1008), .A3(new_n1002), .A4(new_n1071), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT125), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(new_n1074), .A3(KEYINPUT53), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n982), .A2(new_n991), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n738), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1068), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1074), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT53), .B1(new_n1073), .B2(KEYINPUT125), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1068), .B(new_n1077), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1003), .B2(G2078), .ZN(new_n1085));
  AOI21_X1  g660(.A(G301), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1050), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1058), .B(KEYINPUT62), .C1(new_n1060), .C2(new_n1064), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1067), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1024), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1034), .A2(new_n1035), .A3(new_n562), .A4(new_n561), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1027), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1090), .A2(new_n1040), .B1(new_n1032), .B2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1052), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1076), .A2(new_n716), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1002), .A2(new_n981), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(G2067), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n581), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(G1348), .B1(new_n982), .B2(new_n991), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1101), .A2(new_n589), .A3(new_n1098), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT60), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AND2_X1   g678(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1104));
  NOR2_X1   g679(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT58), .B(G1341), .Z(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n1002), .B2(new_n981), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n942), .A2(G1996), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1000), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n546), .B1(new_n1111), .B2(KEYINPUT121), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n1113), .B(new_n1109), .C1(new_n1000), .C2(new_n1110), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1106), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1000), .A2(new_n1110), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1113), .B1(new_n1116), .B2(new_n1109), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1111), .A2(KEYINPUT121), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1117), .A2(new_n546), .A3(new_n1118), .A4(new_n1104), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1103), .A2(new_n1115), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G1956), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1046), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1123));
  XNOR2_X1  g698(.A(G299), .B(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n990), .A2(new_n936), .ZN(new_n1125));
  INV_X1    g700(.A(new_n996), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT56), .B(G2072), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1125), .A2(new_n1002), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1122), .A2(new_n1124), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1122), .A2(new_n1128), .A3(KEYINPUT120), .A4(new_n1124), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1122), .A2(new_n1128), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1124), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1101), .A2(new_n1098), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n581), .A2(KEYINPUT60), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1140), .A2(new_n1129), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1120), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1136), .B1(new_n581), .B2(new_n1141), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1133), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1095), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1065), .A2(new_n1050), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1085), .A2(G301), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1082), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(new_n1078), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n941), .A2(KEYINPUT127), .ZN(new_n1152));
  NOR4_X1   g727(.A1(new_n474), .A2(new_n1084), .A3(new_n1001), .A4(G2078), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n941), .A2(KEYINPUT127), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1155), .A2(new_n996), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n937), .A2(new_n1156), .B1(new_n1076), .B2(new_n738), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n1085), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(G171), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1151), .A2(KEYINPUT54), .A3(new_n1159), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1149), .A2(new_n1157), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1085), .B1(new_n1150), .B2(new_n1078), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1161), .B1(new_n1162), .B2(G171), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1148), .B(new_n1160), .C1(new_n1163), .C2(KEYINPUT54), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1147), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1144), .A2(new_n1095), .A3(new_n1146), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1094), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g742(.A(G290), .B(new_n695), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n962), .B1(new_n961), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n968), .B1(new_n1167), .B2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g745(.A1(G229), .A2(G401), .A3(new_n458), .A4(G227), .ZN(new_n1172));
  NAND3_X1  g746(.A1(new_n844), .A2(new_n930), .A3(new_n1172), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


