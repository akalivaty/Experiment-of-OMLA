//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT9), .ZN(new_n203));
  NAND2_X1  g002(.A1(G71gat), .A2(G78gat), .ZN(new_n204));
  OR2_X1    g003(.A1(G71gat), .A2(G78gat), .ZN(new_n205));
  NAND4_X1  g004(.A1(new_n203), .A2(KEYINPUT97), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT9), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(new_n202), .ZN(new_n209));
  XNOR2_X1  g008(.A(G57gat), .B(G64gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n204), .B(new_n205), .C1(new_n210), .C2(new_n207), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT97), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n206), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT21), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AND2_X1   g015(.A1(G15gat), .A2(G22gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(G15gat), .A2(G22gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT91), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G1gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(KEYINPUT91), .B(G1gat), .C1(new_n217), .C2(new_n218), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(new_n217), .B2(new_n218), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n223), .A2(KEYINPUT92), .A3(G8gat), .A4(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n221), .A2(new_n225), .A3(new_n222), .ZN(new_n227));
  NAND2_X1  g026(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n228));
  OR2_X1    g027(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT98), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT98), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n234), .A3(new_n231), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n214), .A2(new_n215), .ZN(new_n237));
  INV_X1    g036(.A(G127gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n241));
  XNOR2_X1  g040(.A(G155gat), .B(G183gat), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n241), .B(new_n242), .Z(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n239), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(new_n235), .A3(new_n233), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n240), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n244), .B1(new_n240), .B2(new_n246), .ZN(new_n248));
  NAND2_X1  g047(.A1(G231gat), .A2(G233gat), .ZN(new_n249));
  INV_X1    g048(.A(G211gat), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  OR3_X1    g051(.A1(new_n247), .A2(new_n248), .A3(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n247), .B2(new_n248), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G29gat), .ZN(new_n257));
  INV_X1    g056(.A(G36gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(G29gat), .A2(G36gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT14), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n259), .B1(new_n262), .B2(KEYINPUT88), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n260), .B(KEYINPUT14), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT88), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G50gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G43gat), .ZN(new_n269));
  INV_X1    g068(.A(G43gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G50gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n271), .A3(KEYINPUT15), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n259), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n262), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT89), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n270), .B2(G50gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n268), .A2(KEYINPUT89), .A3(G43gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(new_n271), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT15), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT90), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(KEYINPUT90), .A3(new_n282), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n277), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n274), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G85gat), .A2(G92gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT7), .ZN(new_n289));
  XNOR2_X1  g088(.A(G99gat), .B(G106gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(G99gat), .A2(G106gat), .ZN(new_n291));
  INV_X1    g090(.A(G85gat), .ZN(new_n292));
  INV_X1    g091(.A(G92gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(KEYINPUT8), .A2(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n289), .A2(new_n290), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n290), .B1(new_n289), .B2(new_n294), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n287), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G232gat), .ZN(new_n299));
  INV_X1    g098(.A(G233gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT41), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT17), .ZN(new_n304));
  INV_X1    g103(.A(new_n285), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n305), .A2(new_n276), .A3(new_n283), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n272), .B1(new_n263), .B2(new_n266), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n274), .A2(new_n286), .A3(KEYINPUT17), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n289), .A2(new_n294), .ZN(new_n310));
  INV_X1    g109(.A(new_n290), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n289), .A2(new_n290), .A3(new_n294), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n308), .A2(new_n309), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT99), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT99), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n308), .A2(new_n309), .A3(new_n317), .A4(new_n314), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n303), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(G190gat), .B(G218gat), .Z(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT100), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n320), .A2(KEYINPUT100), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n319), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n319), .A2(new_n322), .A3(new_n321), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n301), .A2(KEYINPUT41), .ZN(new_n328));
  XNOR2_X1  g127(.A(G134gat), .B(G162gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n326), .A2(new_n327), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n330), .ZN(new_n332));
  INV_X1    g131(.A(new_n327), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(new_n325), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT65), .ZN(new_n337));
  INV_X1    g136(.A(G190gat), .ZN(new_n338));
  AND2_X1   g137(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g142(.A(KEYINPUT28), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR3_X1   g147(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AND4_X1   g151(.A1(new_n337), .A2(new_n345), .A3(new_n346), .A4(new_n352), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n343), .A2(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n337), .B1(new_n354), .B2(new_n346), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT25), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n338), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G190gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n351), .B(new_n357), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NOR3_X1   g162(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n356), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT64), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n357), .A2(new_n351), .ZN(new_n368));
  INV_X1    g167(.A(new_n360), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(G190gat), .A3(new_n358), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n371));
  INV_X1    g170(.A(G169gat), .ZN(new_n372));
  INV_X1    g171(.A(G176gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n362), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT25), .A4(new_n375), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n366), .A2(new_n367), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n367), .B1(new_n366), .B2(new_n376), .ZN(new_n378));
  OAI22_X1  g177(.A1(new_n353), .A2(new_n355), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G113gat), .ZN(new_n380));
  INV_X1    g179(.A(G120gat), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT1), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(new_n380), .B2(new_n381), .ZN(new_n383));
  INV_X1    g182(.A(G134gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n238), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT66), .B(G127gat), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n383), .B(new_n385), .C1(new_n384), .C2(new_n386), .ZN(new_n387));
  OR2_X1    g186(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(KEYINPUT67), .A2(G113gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(G120gat), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G127gat), .B(G134gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n380), .A2(new_n381), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n387), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n378), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n366), .A2(new_n367), .A3(new_n376), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n345), .A2(new_n346), .A3(new_n352), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT65), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n354), .A2(new_n337), .A3(new_n346), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n402), .A2(new_n406), .A3(new_n395), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n397), .A2(new_n399), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT32), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(G15gat), .B(G43gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G71gat), .ZN(new_n413));
  INV_X1    g212(.A(G99gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n409), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n415), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n408), .B(KEYINPUT32), .C1(new_n410), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n397), .A2(new_n407), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n398), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n399), .B(new_n420), .C1(new_n397), .C2(new_n407), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT71), .B1(new_n419), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n419), .A2(new_n425), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n423), .A2(new_n424), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT71), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n428), .A2(new_n416), .A3(new_n429), .A4(new_n418), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(G22gat), .B(G50gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(KEYINPUT74), .B(KEYINPUT2), .Z(new_n434));
  XOR2_X1   g233(.A(G141gat), .B(G148gat), .Z(new_n435));
  INV_X1    g234(.A(G162gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(G155gat), .ZN(new_n437));
  INV_X1    g236(.A(G155gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(G162gat), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n434), .A2(new_n435), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT76), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n437), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n441), .B1(new_n437), .B2(new_n439), .ZN(new_n443));
  INV_X1    g242(.A(G148gat), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT75), .ZN(new_n445));
  INV_X1    g244(.A(G141gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n444), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n446), .A2(G148gat), .ZN(new_n450));
  OAI22_X1  g249(.A1(new_n442), .A2(new_n443), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT77), .B(G162gat), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n452), .B1(new_n453), .B2(G155gat), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT78), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n454), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n438), .A2(G162gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n436), .A2(G155gat), .ZN(new_n458));
  OAI21_X1  g257(.A(KEYINPUT76), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n437), .A2(new_n439), .A3(new_n441), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT78), .ZN(new_n462));
  INV_X1    g261(.A(new_n448), .ZN(new_n463));
  NOR2_X1   g262(.A1(KEYINPUT75), .A2(G141gat), .ZN(new_n464));
  OAI21_X1  g263(.A(G148gat), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n450), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n456), .A2(new_n461), .A3(new_n462), .A4(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n440), .B1(new_n455), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT3), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT29), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G211gat), .B(G218gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(G197gat), .B(G204gat), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT22), .ZN(new_n474));
  INV_X1    g273(.A(G218gat), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n474), .B1(new_n250), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n472), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n472), .B1(new_n476), .B2(new_n473), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT81), .B1(new_n471), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G228gat), .A2(G233gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT81), .ZN(new_n483));
  AOI211_X1 g282(.A(KEYINPUT3), .B(new_n440), .C1(new_n455), .C2(new_n468), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n483), .B(new_n479), .C1(new_n484), .C2(KEYINPUT29), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n455), .A2(new_n468), .ZN(new_n486));
  INV_X1    g285(.A(new_n440), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT29), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(new_n477), .B2(new_n478), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n488), .B1(KEYINPUT3), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n481), .A2(new_n482), .A3(new_n485), .A4(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT31), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n451), .A2(KEYINPUT78), .A3(new_n454), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n459), .A2(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n462), .B1(new_n496), .B2(new_n456), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n470), .B(new_n487), .C1(new_n495), .C2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n480), .B1(new_n498), .B2(new_n489), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n490), .A2(KEYINPUT82), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT3), .B1(new_n490), .B2(KEYINPUT82), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n469), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(G228gat), .B(G233gat), .C1(new_n499), .C2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n493), .A2(new_n494), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n494), .B1(new_n493), .B2(new_n503), .ZN(new_n505));
  XOR2_X1   g304(.A(G78gat), .B(G106gat), .Z(new_n506));
  NOR3_X1   g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n506), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n482), .B1(new_n499), .B2(new_n483), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n485), .A2(new_n492), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT31), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n493), .A2(new_n494), .A3(new_n503), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n433), .B1(new_n507), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n506), .B1(new_n504), .B2(new_n505), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n512), .A2(new_n513), .A3(new_n508), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(new_n432), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n431), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT35), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT86), .ZN(new_n521));
  XOR2_X1   g320(.A(G8gat), .B(G36gat), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G64gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(new_n293), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n366), .A2(new_n376), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n403), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT73), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n403), .A3(KEYINPUT73), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G226gat), .A2(G233gat), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n532), .B(KEYINPUT72), .Z(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(KEYINPUT29), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n379), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n480), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n402), .A2(new_n406), .A3(new_n533), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n529), .A2(new_n530), .A3(new_n535), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n538), .A2(new_n539), .A3(new_n480), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n525), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n535), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n542), .B1(new_n402), .B2(new_n406), .ZN(new_n543));
  INV_X1    g342(.A(new_n533), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(new_n529), .B2(new_n530), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n479), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n538), .A2(new_n539), .A3(new_n480), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n547), .A3(new_n524), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n541), .A2(KEYINPUT30), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n547), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n551), .A3(new_n525), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G1gat), .B(G29gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT0), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(G57gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G85gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n488), .A2(KEYINPUT3), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(new_n395), .A3(new_n498), .ZN(new_n559));
  NAND2_X1  g358(.A1(G225gat), .A2(G233gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(KEYINPUT5), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT4), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n563), .B1(new_n469), .B2(new_n396), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT80), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n469), .A2(new_n563), .A3(new_n396), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n486), .A2(new_n487), .A3(new_n396), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n565), .A3(KEYINPUT4), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n559), .B(new_n562), .C1(new_n567), .C2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n469), .A2(new_n396), .ZN(new_n573));
  AOI211_X1 g372(.A(new_n440), .B(new_n395), .C1(new_n455), .C2(new_n468), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n561), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT5), .ZN(new_n576));
  NOR3_X1   g375(.A1(new_n568), .A2(KEYINPUT79), .A3(KEYINPUT4), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n469), .A2(new_n470), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(new_n484), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n577), .B1(new_n579), .B2(new_n395), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT79), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(new_n568), .B2(KEYINPUT4), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n561), .B1(new_n582), .B2(new_n566), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n576), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n557), .B1(new_n572), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT6), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n568), .A2(KEYINPUT4), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(KEYINPUT79), .A3(new_n566), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n574), .A2(new_n581), .A3(new_n563), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n588), .A2(new_n559), .A3(new_n560), .A4(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n575), .A2(KEYINPUT5), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n557), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n571), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n585), .A2(new_n586), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g394(.A(KEYINPUT6), .B(new_n557), .C1(new_n572), .C2(new_n584), .ZN(new_n596));
  AOI211_X1 g395(.A(KEYINPUT35), .B(new_n553), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n519), .B(new_n521), .C1(new_n597), .C2(KEYINPUT86), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT70), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n419), .A2(new_n425), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n425), .B1(new_n419), .B2(new_n599), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n516), .A2(new_n432), .A3(new_n517), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n432), .B1(new_n516), .B2(new_n517), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n553), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n594), .A2(new_n586), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n593), .B1(new_n592), .B2(new_n571), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n596), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT35), .B1(new_n606), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n515), .A2(new_n518), .ZN(new_n615));
  OR3_X1    g414(.A1(new_n573), .A2(new_n574), .A3(new_n561), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n566), .A2(new_n565), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n587), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n618), .A2(new_n569), .B1(new_n395), .B2(new_n579), .ZN(new_n619));
  OAI211_X1 g418(.A(KEYINPUT39), .B(new_n616), .C1(new_n619), .C2(new_n560), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT84), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT40), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n557), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n559), .B1(new_n567), .B2(new_n570), .ZN(new_n624));
  XOR2_X1   g423(.A(KEYINPUT83), .B(KEYINPUT39), .Z(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n561), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n620), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n621), .A2(new_n622), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n620), .A2(new_n628), .A3(new_n623), .A4(new_n626), .ZN(new_n631));
  NAND4_X1  g430(.A1(new_n630), .A2(new_n585), .A3(new_n553), .A4(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT37), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n525), .B1(new_n550), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n546), .A2(KEYINPUT37), .A3(new_n547), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n636), .A2(KEYINPUT38), .B1(new_n550), .B2(new_n525), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n538), .A2(new_n539), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n479), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n534), .A2(new_n480), .A3(new_n536), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT37), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT85), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n642), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n634), .A4(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n595), .A2(new_n637), .A3(new_n596), .A4(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n615), .A2(new_n632), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n612), .A2(new_n518), .A3(new_n515), .ZN(new_n649));
  OAI21_X1  g448(.A(KEYINPUT36), .B1(new_n601), .B2(new_n602), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT36), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n426), .A2(new_n651), .A3(new_n427), .A4(new_n430), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  AOI211_X1 g453(.A(new_n256), .B(new_n336), .C1(new_n614), .C2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n231), .A2(new_n274), .A3(new_n286), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n230), .B(new_n226), .C1(new_n306), .C2(new_n307), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT95), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(G229gat), .A2(G233gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT94), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n661), .B(KEYINPUT13), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n287), .A2(KEYINPUT95), .A3(new_n230), .A4(new_n226), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n659), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(KEYINPUT96), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n659), .A2(new_n667), .A3(new_n663), .A4(new_n664), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT93), .ZN(new_n670));
  INV_X1    g469(.A(new_n230), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n228), .B1(new_n227), .B2(new_n229), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n226), .A2(new_n230), .A3(KEYINPUT93), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n673), .A2(new_n308), .A3(new_n309), .A4(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n661), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n676), .A3(new_n657), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT18), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT18), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n675), .A2(new_n679), .A3(new_n676), .A4(new_n657), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT87), .B(G197gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(G113gat), .B(G141gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT11), .B(G169gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT12), .Z(new_n687));
  AND3_X1   g486(.A1(new_n669), .A2(new_n681), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n669), .B2(new_n681), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n297), .A2(new_n209), .A3(new_n213), .A4(new_n206), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n214), .A2(new_n314), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT10), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  OR3_X1    g493(.A1(new_n214), .A2(new_n314), .A3(new_n693), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(G230gat), .A2(G233gat), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT101), .Z(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n691), .A2(new_n692), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n698), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(G120gat), .B(G148gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(new_n373), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G204gat), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n700), .A2(new_n702), .A3(new_n706), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n690), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n655), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n610), .A2(new_n611), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT102), .B(G1gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1324gat));
  AND2_X1   g515(.A1(new_n712), .A2(new_n553), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n718));
  OR3_X1    g517(.A1(new_n718), .A2(new_n224), .A3(KEYINPUT42), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n224), .B1(new_n718), .B2(KEYINPUT42), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n721), .A2(G8gat), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n717), .A2(KEYINPUT42), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(G8gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(G1325gat));
  AND3_X1   g524(.A1(new_n426), .A2(new_n427), .A3(new_n430), .ZN(new_n726));
  AOI21_X1  g525(.A(G15gat), .B1(new_n712), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n650), .A2(new_n652), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(G15gat), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(new_n712), .B2(new_n729), .ZN(G1326gat));
  INV_X1    g529(.A(new_n615), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n712), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT43), .B(G22gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1327gat));
  AOI21_X1  g533(.A(new_n335), .B1(new_n614), .B2(new_n654), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n256), .A2(new_n711), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n738), .A2(new_n257), .A3(new_n713), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT45), .ZN(new_n740));
  AOI211_X1 g539(.A(KEYINPUT44), .B(new_n335), .C1(new_n614), .C2(new_n654), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n553), .B1(new_n595), .B2(new_n596), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT86), .B1(new_n743), .B2(new_n520), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n726), .B(new_n521), .C1(new_n604), .C2(new_n605), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n419), .A2(new_n599), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n428), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n600), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n749), .B1(new_n518), .B2(new_n515), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n520), .B1(new_n750), .B2(new_n743), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n654), .B1(new_n746), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n742), .B1(new_n752), .B2(new_n336), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n741), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n737), .ZN(new_n755));
  INV_X1    g554(.A(new_n713), .ZN(new_n756));
  OAI21_X1  g555(.A(G29gat), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n757), .ZN(G1328gat));
  NAND3_X1  g557(.A1(new_n738), .A2(new_n258), .A3(new_n553), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT46), .Z(new_n760));
  OAI21_X1  g559(.A(G36gat), .B1(new_n755), .B2(new_n607), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1329gat));
  NAND2_X1  g561(.A1(new_n728), .A2(G43gat), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n738), .A2(new_n726), .ZN(new_n764));
  OAI22_X1  g563(.A1(new_n755), .A2(new_n763), .B1(G43gat), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g565(.A(G50gat), .B1(new_n755), .B2(new_n615), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n738), .A2(new_n268), .A3(new_n731), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT48), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n767), .B(new_n770), .C1(new_n768), .C2(KEYINPUT48), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(G1331gat));
  INV_X1    g574(.A(new_n690), .ZN(new_n776));
  INV_X1    g575(.A(new_n710), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n655), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT105), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT105), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n655), .A2(new_n781), .A3(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n713), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n553), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n788));
  XOR2_X1   g587(.A(KEYINPUT49), .B(G64gat), .Z(new_n789));
  OAI21_X1  g588(.A(new_n788), .B1(new_n787), .B2(new_n789), .ZN(G1333gat));
  INV_X1    g589(.A(G71gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n783), .B2(new_n431), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n780), .A2(G71gat), .A3(new_n728), .A4(new_n782), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT50), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n792), .A2(new_n796), .A3(new_n793), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(G1334gat));
  NAND2_X1  g597(.A1(new_n784), .A2(new_n731), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g599(.A1(new_n255), .A2(new_n776), .A3(new_n777), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n754), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G85gat), .B1(new_n802), .B2(new_n756), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n255), .A2(new_n776), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n735), .A2(new_n804), .ZN(new_n805));
  XOR2_X1   g604(.A(new_n805), .B(KEYINPUT51), .Z(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n710), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n713), .A2(new_n292), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(G1336gat));
  AND2_X1   g608(.A1(new_n754), .A2(new_n801), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n293), .B1(new_n810), .B2(new_n553), .ZN(new_n811));
  OR2_X1    g610(.A1(KEYINPUT106), .A2(KEYINPUT51), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n735), .B2(new_n804), .ZN(new_n813));
  AND4_X1   g612(.A1(new_n752), .A2(new_n336), .A3(new_n804), .A4(new_n812), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n607), .A2(G92gat), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n815), .A2(new_n777), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT52), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n807), .B2(new_n817), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n811), .B2(new_n821), .ZN(G1337gat));
  NAND3_X1  g621(.A1(new_n810), .A2(KEYINPUT107), .A3(new_n728), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT107), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n802), .B2(new_n653), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(G99gat), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n726), .A2(new_n414), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n807), .B2(new_n827), .ZN(G1338gat));
  NOR3_X1   g627(.A1(new_n615), .A2(G106gat), .A3(new_n777), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n806), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n731), .B(new_n801), .C1(new_n741), .C2(new_n753), .ZN(new_n832));
  XNOR2_X1  g631(.A(KEYINPUT108), .B(G106gat), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n830), .A2(new_n831), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n829), .B1(new_n813), .B2(new_n814), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT109), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT109), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n839), .B(new_n829), .C1(new_n813), .C2(new_n814), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n835), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n841), .A2(KEYINPUT110), .A3(KEYINPUT53), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT110), .B1(new_n841), .B2(KEYINPUT53), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n836), .B1(new_n842), .B2(new_n843), .ZN(G1339gat));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n694), .A2(new_n695), .A3(new_n698), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT54), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n698), .B1(new_n694), .B2(new_n695), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n696), .A2(new_n851), .A3(new_n699), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n707), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n846), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n700), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n706), .B1(new_n849), .B2(new_n851), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(KEYINPUT55), .A3(new_n856), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n854), .A2(new_n709), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n858), .B1(new_n689), .B2(new_n688), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n669), .A2(new_n681), .A3(new_n687), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n663), .B1(new_n659), .B2(new_n664), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n676), .B1(new_n675), .B2(new_n657), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n686), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n860), .A2(new_n710), .A3(new_n865), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n859), .A2(new_n866), .B1(new_n331), .B2(new_n334), .ZN(new_n867));
  AOI22_X1  g666(.A1(new_n666), .A2(new_n668), .B1(new_n678), .B2(new_n680), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n868), .A2(new_n687), .B1(new_n864), .B2(new_n863), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n869), .A2(new_n331), .A3(new_n858), .A4(new_n334), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n845), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n854), .A2(new_n709), .A3(new_n857), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n669), .A2(new_n681), .ZN(new_n874));
  INV_X1    g673(.A(new_n687), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n873), .B1(new_n876), .B2(new_n860), .ZN(new_n877));
  INV_X1    g676(.A(new_n866), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n335), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n879), .A2(KEYINPUT112), .A3(new_n870), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n872), .A2(new_n256), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n255), .A2(new_n777), .A3(new_n335), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(new_n776), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n756), .B(new_n553), .C1(new_n881), .C2(new_n884), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(new_n519), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n380), .B1(new_n886), .B2(new_n776), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n885), .A2(new_n750), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n690), .B1(new_n388), .B2(new_n389), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT113), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n890), .B(new_n891), .ZN(G1340gat));
  NAND3_X1  g691(.A1(new_n888), .A2(new_n381), .A3(new_n710), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n886), .A2(new_n710), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n381), .ZN(G1341gat));
  NAND2_X1  g694(.A1(new_n888), .A2(new_n255), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n256), .A2(new_n386), .ZN(new_n897));
  AOI22_X1  g696(.A1(new_n896), .A2(new_n386), .B1(new_n886), .B2(new_n897), .ZN(G1342gat));
  NOR2_X1   g697(.A1(new_n335), .A2(new_n553), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT114), .Z(new_n900));
  AOI211_X1 g699(.A(new_n756), .B(new_n900), .C1(new_n884), .C2(new_n881), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n384), .A3(new_n750), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT56), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n384), .B1(new_n886), .B2(new_n336), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n903), .A2(new_n904), .ZN(G1343gat));
  NOR2_X1   g704(.A1(new_n463), .A2(new_n464), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n881), .A2(new_n884), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n731), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(KEYINPUT115), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT116), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n877), .B2(new_n878), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT116), .B(new_n866), .C1(new_n690), .C2(new_n873), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n335), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n255), .B1(new_n914), .B2(new_n870), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n731), .B1(new_n915), .B2(new_n883), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n916), .A2(new_n909), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT115), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n615), .B1(new_n881), .B2(new_n884), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(KEYINPUT57), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n910), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n728), .A2(new_n756), .A3(new_n553), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n906), .B1(new_n923), .B2(new_n690), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n653), .A2(new_n731), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT117), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n885), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n776), .A2(new_n446), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT118), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT58), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT58), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n924), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1344gat));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n710), .A3(new_n922), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n444), .A2(KEYINPUT59), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n907), .A2(KEYINPUT57), .A3(new_n731), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n916), .A2(new_n909), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(new_n710), .A3(new_n922), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(G148gat), .ZN(new_n943));
  AOI22_X1  g742(.A1(new_n937), .A2(new_n938), .B1(new_n943), .B2(KEYINPUT59), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n444), .A3(new_n710), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n936), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n937), .A2(new_n938), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n943), .A2(KEYINPUT59), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(KEYINPUT119), .A3(new_n945), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n947), .A2(new_n951), .ZN(G1345gat));
  AOI21_X1  g751(.A(G155gat), .B1(new_n927), .B2(new_n255), .ZN(new_n953));
  INV_X1    g752(.A(new_n923), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n256), .A2(new_n438), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(G1346gat));
  NAND3_X1  g755(.A1(new_n954), .A2(KEYINPUT120), .A3(new_n336), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT120), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n958), .B1(new_n923), .B2(new_n335), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n957), .A2(new_n453), .A3(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(new_n453), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n901), .A2(new_n961), .A3(new_n926), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1347gat));
  AOI21_X1  g762(.A(new_n713), .B1(new_n881), .B2(new_n884), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n964), .A2(new_n553), .A3(new_n519), .ZN(new_n965));
  OAI21_X1  g764(.A(G169gat), .B1(new_n965), .B2(new_n690), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT121), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n964), .B(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n968), .A2(new_n553), .A3(new_n750), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n776), .A2(new_n372), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(G1348gat));
  NOR3_X1   g770(.A1(new_n965), .A2(new_n373), .A3(new_n777), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n969), .A2(new_n777), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n972), .B1(new_n973), .B2(new_n373), .ZN(G1349gat));
  INV_X1    g773(.A(KEYINPUT60), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n255), .B1(new_n340), .B2(new_n339), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n968), .A2(new_n553), .A3(new_n750), .A4(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT122), .ZN(new_n979));
  OAI21_X1  g778(.A(G183gat), .B1(new_n965), .B2(new_n256), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n979), .B1(new_n978), .B2(new_n980), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n975), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n978), .A2(new_n980), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT122), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n986), .A2(KEYINPUT60), .A3(new_n981), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n984), .A2(new_n987), .ZN(G1350gat));
  OAI21_X1  g787(.A(G190gat), .B1(new_n965), .B2(new_n335), .ZN(new_n989));
  XOR2_X1   g788(.A(KEYINPUT123), .B(KEYINPUT61), .Z(new_n990));
  XNOR2_X1  g789(.A(new_n989), .B(new_n990), .ZN(new_n991));
  OR2_X1    g790(.A1(new_n969), .A2(G190gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n991), .B1(new_n992), .B2(new_n335), .ZN(G1351gat));
  NOR2_X1   g792(.A1(new_n728), .A2(new_n607), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(new_n731), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n995), .B(KEYINPUT124), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n968), .A2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(G197gat), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n997), .A2(new_n998), .A3(new_n776), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n994), .A2(new_n756), .ZN(new_n1000));
  XOR2_X1   g799(.A(new_n1000), .B(KEYINPUT125), .Z(new_n1001));
  AOI21_X1  g800(.A(new_n1001), .B1(new_n940), .B2(new_n939), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n1002), .A2(new_n776), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n999), .B1(new_n998), .B2(new_n1003), .ZN(G1352gat));
  INV_X1    g803(.A(G204gat), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n997), .A2(new_n1005), .A3(new_n710), .ZN(new_n1006));
  OR2_X1    g805(.A1(new_n1006), .A2(KEYINPUT62), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n941), .A2(new_n710), .ZN(new_n1008));
  OAI21_X1  g807(.A(G204gat), .B1(new_n1008), .B2(new_n1001), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1006), .A2(KEYINPUT62), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(G1353gat));
  NAND2_X1  g810(.A1(new_n1002), .A2(new_n255), .ZN(new_n1012));
  AOI22_X1  g811(.A1(new_n1012), .A2(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n1013));
  OR2_X1    g812(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1014));
  OR2_X1    g813(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n997), .A2(new_n250), .A3(new_n255), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n1015), .A2(new_n1016), .A3(new_n1017), .ZN(G1354gat));
  AOI21_X1  g817(.A(G218gat), .B1(new_n997), .B2(new_n336), .ZN(new_n1019));
  NOR2_X1   g818(.A1(new_n335), .A2(new_n475), .ZN(new_n1020));
  XNOR2_X1  g819(.A(new_n1020), .B(KEYINPUT127), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1019), .B1(new_n1002), .B2(new_n1021), .ZN(G1355gat));
endmodule


