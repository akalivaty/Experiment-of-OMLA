//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n792, new_n793,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT86), .ZN(new_n206));
  AOI21_X1  g005(.A(G8gat), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(KEYINPUT86), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n204), .A2(KEYINPUT85), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT85), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n210), .B(G8gat), .C1(new_n211), .C2(new_n205), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT17), .ZN(new_n214));
  INV_X1    g013(.A(G50gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G43gat), .ZN(new_n216));
  INV_X1    g015(.A(G43gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G50gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT15), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT82), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n218), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT15), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G29gat), .A2(G36gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT14), .ZN(new_n227));
  INV_X1    g026(.A(G29gat), .ZN(new_n228));
  INV_X1    g027(.A(G36gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT83), .ZN(new_n231));
  NOR3_X1   g030(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT83), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n222), .A2(new_n220), .A3(new_n223), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n225), .A2(new_n226), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT84), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n235), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n241), .B1(KEYINPUT83), .B2(new_n230), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n242), .A2(new_n234), .B1(G29gat), .B2(G36gat), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n243), .A2(KEYINPUT84), .A3(new_n225), .A4(new_n237), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n241), .A2(new_n232), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n246), .A2(KEYINPUT81), .B1(G29gat), .B2(G36gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT81), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n241), .B2(new_n232), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n219), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n214), .B1(new_n245), .B2(new_n251), .ZN(new_n252));
  AOI211_X1 g051(.A(KEYINPUT17), .B(new_n250), .C1(new_n240), .C2(new_n244), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n213), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n245), .A2(new_n251), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n209), .A2(new_n212), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G229gat), .A2(G233gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n254), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n255), .B(new_n256), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n258), .B(KEYINPUT13), .Z(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n254), .A2(KEYINPUT18), .A3(new_n257), .A4(new_n258), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n261), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  XOR2_X1   g065(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n267));
  XNOR2_X1  g066(.A(G113gat), .B(G141gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G169gat), .B(G197gat), .Z(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT12), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n261), .A2(new_n264), .A3(new_n265), .A4(new_n272), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT24), .ZN(new_n278));
  INV_X1    g077(.A(G183gat), .ZN(new_n279));
  INV_X1    g078(.A(G190gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n281), .B(new_n282), .C1(G183gat), .C2(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  INV_X1    g083(.A(G169gat), .ZN(new_n285));
  INV_X1    g084(.A(G176gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n283), .B1(KEYINPUT65), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(KEYINPUT65), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n288), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT25), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(KEYINPUT64), .B(G169gat), .Z(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(KEYINPUT23), .A3(new_n286), .ZN(new_n296));
  INV_X1    g095(.A(new_n284), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(KEYINPUT25), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n296), .A2(new_n292), .A3(new_n283), .A4(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n287), .B(KEYINPUT26), .ZN(new_n300));
  OAI22_X1  g099(.A1(new_n300), .A2(new_n297), .B1(new_n279), .B2(new_n280), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT27), .B(G183gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n280), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT28), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n294), .B(new_n299), .C1(new_n301), .C2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G113gat), .B(G120gat), .ZN(new_n306));
  OR3_X1    g105(.A1(new_n306), .A2(KEYINPUT66), .A3(KEYINPUT1), .ZN(new_n307));
  OAI21_X1  g106(.A(KEYINPUT66), .B1(new_n306), .B2(KEYINPUT1), .ZN(new_n308));
  XOR2_X1   g107(.A(G127gat), .B(G134gat), .Z(new_n309));
  NAND3_X1  g108(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n308), .A2(new_n309), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n305), .B(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G227gat), .ZN(new_n314));
  INV_X1    g113(.A(G233gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n316), .B(KEYINPUT34), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G15gat), .B(G43gat), .Z(new_n319));
  XNOR2_X1  g118(.A(G71gat), .B(G99gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n322), .B2(KEYINPUT33), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT32), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n323), .A2(new_n325), .ZN(new_n327));
  OAI211_X1 g126(.A(KEYINPUT67), .B(new_n318), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  OR2_X1    g127(.A1(new_n323), .A2(new_n325), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n323), .A2(new_n325), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(new_n317), .A3(new_n330), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n328), .B(new_n331), .C1(KEYINPUT67), .C2(new_n318), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT36), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n318), .B1(new_n326), .B2(new_n327), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n331), .ZN(new_n335));
  OR2_X1    g134(.A1(new_n335), .A2(KEYINPUT36), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  XOR2_X1   g136(.A(KEYINPUT69), .B(G141gat), .Z(new_n338));
  INV_X1    g137(.A(G148gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT70), .B(G148gat), .ZN(new_n340));
  INV_X1    g139(.A(G141gat), .ZN(new_n341));
  OAI22_X1  g140(.A1(new_n338), .A2(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343));
  OR2_X1    g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(KEYINPUT2), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G141gat), .B(G148gat), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n343), .B(new_n344), .C1(new_n347), .C2(KEYINPUT2), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n346), .A2(new_n350), .A3(new_n348), .ZN(new_n352));
  OR3_X1    g151(.A1(new_n351), .A2(new_n312), .A3(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(KEYINPUT5), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n349), .A2(new_n312), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n356), .A2(KEYINPUT4), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n356), .A2(KEYINPUT4), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n353), .B(new_n355), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OR2_X1    g159(.A1(new_n356), .A2(KEYINPUT4), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT71), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n361), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  OR3_X1    g162(.A1(new_n356), .A2(new_n362), .A3(KEYINPUT4), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n354), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n353), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n349), .B(new_n312), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n354), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT5), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n360), .B1(new_n366), .B2(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(KEYINPUT72), .B(KEYINPUT0), .Z(new_n372));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  XOR2_X1   g173(.A(G57gat), .B(G85gat), .Z(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n351), .A2(new_n312), .A3(new_n352), .ZN(new_n379));
  AOI211_X1 g178(.A(new_n354), .B(new_n379), .C1(new_n363), .C2(new_n364), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n376), .B(new_n359), .C1(new_n380), .C2(new_n369), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT73), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n378), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT73), .B1(new_n371), .B2(new_n376), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n377), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OR3_X1    g184(.A1(new_n371), .A2(KEYINPUT6), .A3(new_n376), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT29), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n305), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(G197gat), .B(G204gat), .Z(new_n392));
  INV_X1    g191(.A(G211gat), .ZN(new_n393));
  INV_X1    g192(.A(G218gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT22), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n393), .A2(new_n394), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n392), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n400), .B(new_n395), .C1(new_n392), .C2(new_n396), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n305), .A2(new_n388), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n391), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G8gat), .B(G36gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(G64gat), .B(G92gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT68), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n390), .A2(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n305), .A2(new_n389), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n405), .B1(new_n413), .B2(new_n388), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n414), .B2(new_n411), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n406), .B(new_n410), .C1(new_n415), .C2(new_n404), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT30), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n406), .B1(new_n415), .B2(new_n404), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n409), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n416), .A2(new_n417), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n418), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT74), .B1(new_n387), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n404), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(new_n352), .B2(KEYINPUT29), .ZN(new_n425));
  AND2_X1   g224(.A1(G228gat), .A2(G233gat), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT3), .B1(new_n404), .B2(new_n389), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n425), .B(new_n426), .C1(new_n349), .C2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n403), .B(KEYINPUT75), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n389), .B1(new_n429), .B2(new_n401), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n349), .B1(new_n430), .B2(new_n350), .ZN(new_n431));
  INV_X1    g230(.A(new_n425), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n428), .B1(new_n433), .B2(new_n426), .ZN(new_n434));
  XNOR2_X1  g233(.A(G78gat), .B(G106gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(KEYINPUT31), .B(G50gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n435), .B(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT76), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n438), .A3(G22gat), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(G22gat), .B2(new_n437), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n434), .B(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n422), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT74), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n442), .A2(new_n385), .A3(new_n443), .A4(new_n386), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n423), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n422), .A2(KEYINPUT77), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT77), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n418), .A2(new_n448), .A3(new_n420), .A4(new_n421), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n358), .A2(new_n357), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n354), .B1(new_n451), .B2(new_n379), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n452), .A2(KEYINPUT39), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n452), .B(KEYINPUT39), .C1(new_n354), .C2(new_n367), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n454), .A3(new_n376), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT40), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(KEYINPUT78), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n455), .A2(new_n456), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n450), .A2(new_n377), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n419), .A2(KEYINPUT37), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT37), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n462), .B(new_n406), .C1(new_n415), .C2(new_n404), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n409), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT38), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n391), .A2(new_n424), .A3(new_n405), .ZN(new_n466));
  OAI211_X1 g265(.A(KEYINPUT37), .B(new_n466), .C1(new_n415), .C2(new_n424), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n463), .A2(new_n467), .A3(new_n468), .A4(new_n409), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT79), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n387), .A2(new_n416), .A3(new_n465), .A4(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n441), .B1(new_n460), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n337), .B1(new_n446), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n441), .B1(new_n334), .B2(new_n331), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(new_n447), .A3(new_n449), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n475), .A2(KEYINPUT35), .A3(new_n387), .ZN(new_n476));
  INV_X1    g275(.A(new_n441), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n332), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n423), .A2(new_n478), .A3(new_n444), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n476), .B1(new_n479), .B2(KEYINPUT35), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n277), .B1(new_n473), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G230gat), .A2(G233gat), .ZN(new_n483));
  INV_X1    g282(.A(G57gat), .ZN(new_n484));
  INV_X1    g283(.A(G64gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(G57gat), .A2(G64gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(G71gat), .A2(G78gat), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n486), .B(new_n487), .C1(new_n489), .C2(KEYINPUT9), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(KEYINPUT88), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT87), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n492), .B1(G71gat), .B2(G78gat), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT88), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(G71gat), .A3(G78gat), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n491), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n493), .B1(new_n491), .B2(new_n495), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n490), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OR3_X1    g297(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT89), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n485), .B1(new_n484), .B2(KEYINPUT89), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT9), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n501), .A2(G71gat), .A3(G78gat), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n499), .B(new_n500), .C1(new_n489), .C2(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G99gat), .ZN(new_n505));
  INV_X1    g304(.A(G106gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508));
  AND2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT96), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(KEYINPUT94), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT94), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n513), .A2(G99gat), .A3(G106gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT8), .ZN(new_n515));
  INV_X1    g314(.A(G92gat), .ZN(new_n516));
  AND2_X1   g315(.A1(KEYINPUT95), .A2(G85gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(KEYINPUT95), .A2(G85gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n507), .A2(new_n510), .A3(new_n508), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT93), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(G85gat), .A3(G92gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n526), .A3(KEYINPUT7), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT7), .B1(new_n524), .B2(new_n526), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n511), .B1(new_n522), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n526), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(new_n527), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n509), .A2(new_n510), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n535), .A2(new_n521), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n504), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n530), .A3(new_n511), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n536), .B1(new_n535), .B2(new_n521), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n498), .A2(new_n503), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n483), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT100), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G120gat), .B(G148gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT101), .ZN(new_n547));
  XNOR2_X1  g346(.A(G176gat), .B(G204gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n543), .B2(new_n544), .ZN(new_n550));
  INV_X1    g349(.A(new_n483), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT10), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n538), .A2(new_n552), .A3(new_n542), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n539), .A2(new_n540), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(KEYINPUT10), .A3(new_n504), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n545), .A2(new_n550), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n549), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n556), .B2(new_n543), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n504), .A2(KEYINPUT21), .ZN(new_n563));
  XOR2_X1   g362(.A(G183gat), .B(G211gat), .Z(new_n564));
  XOR2_X1   g363(.A(new_n563), .B(new_n564), .Z(new_n565));
  NAND2_X1  g364(.A1(new_n504), .A2(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n213), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT90), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT90), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n213), .A2(new_n569), .A3(new_n566), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n571), .B1(new_n568), .B2(new_n570), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n565), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n574), .ZN(new_n576));
  INV_X1    g375(.A(new_n565), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G127gat), .B(G155gat), .Z(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n575), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n575), .B2(new_n578), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n554), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(new_n252), .B2(new_n253), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT97), .ZN(new_n587));
  AND2_X1   g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n255), .A2(new_n554), .B1(KEYINPUT41), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT97), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n590), .B(new_n585), .C1(new_n252), .C2(new_n253), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n587), .A2(new_n589), .A3(new_n591), .A4(new_n593), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n595), .A2(KEYINPUT98), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT98), .B1(new_n595), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n588), .A2(KEYINPUT41), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n597), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n598), .A2(new_n603), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n584), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT99), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n595), .A2(new_n596), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT98), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n603), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n595), .A2(KEYINPUT98), .A3(new_n596), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n605), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(KEYINPUT99), .A3(new_n584), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n609), .A2(new_n617), .ZN(new_n618));
  AND3_X1   g417(.A1(new_n482), .A2(new_n562), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n387), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n450), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT42), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT16), .B(G8gat), .ZN(new_n624));
  OR3_X1    g423(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(G8gat), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n623), .B1(new_n622), .B2(new_n624), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(G1325gat));
  AOI21_X1  g427(.A(G15gat), .B1(new_n619), .B2(new_n335), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT102), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n333), .A2(new_n336), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n333), .B2(new_n336), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n633), .A2(G15gat), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n629), .B1(new_n619), .B2(new_n634), .ZN(G1326gat));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n441), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT43), .B(G22gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1327gat));
  INV_X1    g437(.A(new_n584), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n616), .A2(new_n561), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n482), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n228), .A3(new_n387), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT103), .B(KEYINPUT45), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n460), .A2(new_n471), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n477), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n445), .ZN(new_n648));
  INV_X1    g447(.A(new_n633), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n480), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n645), .B1(new_n650), .B2(new_n616), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n473), .A2(new_n481), .ZN(new_n652));
  INV_X1    g451(.A(new_n616), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(KEYINPUT44), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n584), .B(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n657), .A2(new_n561), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n651), .A2(new_n276), .A3(new_n654), .A4(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n385), .B2(new_n386), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n644), .B1(new_n660), .B2(new_n228), .ZN(G1328gat));
  NAND3_X1  g460(.A1(new_n641), .A2(new_n229), .A3(new_n450), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n662), .B(KEYINPUT46), .Z(new_n663));
  INV_X1    g462(.A(new_n450), .ZN(new_n664));
  OAI21_X1  g463(.A(G36gat), .B1(new_n659), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(G1329gat));
  OAI21_X1  g465(.A(G43gat), .B1(new_n659), .B2(new_n649), .ZN(new_n667));
  INV_X1    g466(.A(new_n335), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(G43gat), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n482), .A2(new_n639), .A3(new_n640), .A4(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n667), .A2(KEYINPUT47), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n670), .B(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(KEYINPUT47), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI211_X1 g475(.A(KEYINPUT106), .B(KEYINPUT47), .C1(new_n667), .C2(new_n673), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n671), .B1(new_n676), .B2(new_n677), .ZN(G1330gat));
  AOI21_X1  g477(.A(G50gat), .B1(new_n641), .B2(new_n441), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n659), .A2(new_n215), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(new_n441), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g481(.A1(new_n618), .A2(new_n561), .A3(new_n277), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT107), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n633), .B1(new_n647), .B2(new_n445), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(new_n480), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT108), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n387), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(G57gat), .ZN(G1332gat));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n686), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n691), .A2(new_n664), .ZN(new_n692));
  NOR2_X1   g491(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n693));
  AND2_X1   g492(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(new_n692), .B2(new_n693), .ZN(G1333gat));
  XNOR2_X1  g495(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n633), .A2(G71gat), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n691), .A2(new_n668), .ZN(new_n699));
  OAI221_X1 g498(.A(new_n697), .B1(new_n691), .B2(new_n698), .C1(new_n699), .C2(G71gat), .ZN(new_n700));
  INV_X1    g499(.A(new_n697), .ZN(new_n701));
  AOI21_X1  g500(.A(G71gat), .B1(new_n687), .B2(new_n335), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n691), .A2(new_n698), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n700), .A2(new_n704), .ZN(G1334gat));
  NAND2_X1  g504(.A1(new_n687), .A2(new_n441), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g506(.A1(new_n584), .A2(new_n276), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n651), .A2(new_n561), .A3(new_n654), .A4(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n385), .B2(new_n386), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n517), .A2(new_n518), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n653), .B(new_n708), .C1(new_n685), .C2(new_n480), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT51), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n387), .A2(new_n711), .A3(new_n561), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT110), .Z(new_n719));
  OAI22_X1  g518(.A1(new_n710), .A2(new_n711), .B1(new_n717), .B2(new_n719), .ZN(G1336gat));
  NAND4_X1  g519(.A1(new_n716), .A2(new_n516), .A3(new_n561), .A4(new_n450), .ZN(new_n721));
  OAI21_X1  g520(.A(G92gat), .B1(new_n709), .B2(new_n664), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1337gat));
  NOR3_X1   g524(.A1(new_n709), .A2(new_n505), .A3(new_n649), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n716), .A2(new_n561), .A3(new_n335), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(new_n505), .ZN(G1338gat));
  OAI21_X1  g527(.A(G106gat), .B1(new_n709), .B2(new_n477), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n716), .A2(new_n506), .A3(new_n561), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(new_n477), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT53), .ZN(new_n732));
  OR3_X1    g531(.A1(new_n709), .A2(KEYINPUT112), .A3(new_n477), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT112), .B1(new_n709), .B2(new_n477), .ZN(new_n734));
  AND3_X1   g533(.A1(new_n733), .A2(G106gat), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT53), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n730), .B2(new_n477), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n732), .B1(new_n735), .B2(new_n737), .ZN(G1339gat));
  NAND4_X1  g537(.A1(new_n609), .A2(new_n562), .A3(new_n277), .A4(new_n617), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n262), .A2(new_n263), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n258), .B1(new_n254), .B2(new_n257), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n271), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT115), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT115), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n744), .B(new_n271), .C1(new_n740), .C2(new_n741), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n743), .A2(new_n275), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n615), .A2(new_n605), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n553), .A2(new_n555), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n483), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n553), .A2(new_n555), .A3(new_n551), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n749), .A2(KEYINPUT54), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT113), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n749), .A2(new_n753), .A3(new_n750), .A4(KEYINPUT54), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT54), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n549), .B1(new_n556), .B2(new_n757), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n755), .A2(new_n756), .A3(KEYINPUT55), .A4(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n752), .A2(new_n758), .A3(new_n754), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n557), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT114), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n759), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n747), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n276), .A2(new_n759), .A3(new_n762), .A4(new_n763), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n743), .A2(new_n561), .A3(new_n275), .A4(new_n745), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n766), .A2(new_n767), .B1(new_n615), .B2(new_n605), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n656), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n739), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(new_n387), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n478), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(KEYINPUT116), .A3(new_n478), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n774), .A2(new_n664), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT117), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(G113gat), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n774), .A2(new_n664), .A3(new_n775), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT117), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n778), .A2(new_n779), .A3(new_n276), .A4(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n771), .A2(new_n664), .A3(new_n474), .ZN(new_n783));
  OAI21_X1  g582(.A(G113gat), .B1(new_n783), .B2(new_n277), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1340gat));
  INV_X1    g586(.A(G120gat), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n783), .A2(new_n788), .A3(new_n562), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n778), .A2(new_n561), .A3(new_n781), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n790), .B2(new_n788), .ZN(G1341gat));
  AOI21_X1  g590(.A(G127gat), .B1(new_n776), .B2(new_n584), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n783), .A2(new_n656), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(G127gat), .B2(new_n793), .ZN(G1342gat));
  NOR3_X1   g593(.A1(new_n780), .A2(G134gat), .A3(new_n616), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT56), .ZN(new_n796));
  OAI21_X1  g595(.A(G134gat), .B1(new_n783), .B2(new_n616), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(G1343gat));
  INV_X1    g597(.A(KEYINPUT122), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n387), .B(new_n664), .C1(new_n631), .C2(new_n632), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n801), .A2(new_n441), .A3(new_n770), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n802), .A2(G141gat), .A3(new_n277), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n770), .A2(new_n441), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n639), .B1(new_n765), .B2(new_n768), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n739), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n477), .A2(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n808), .A2(KEYINPUT119), .A3(new_n809), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n806), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(new_n276), .A3(new_n801), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n803), .B1(new_n815), .B2(new_n338), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT121), .ZN(new_n817));
  XNOR2_X1  g616(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(new_n817), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT121), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n338), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT119), .B1(new_n808), .B2(new_n809), .ZN(new_n824));
  INV_X1    g623(.A(new_n809), .ZN(new_n825));
  AOI211_X1 g624(.A(new_n811), .B(new_n825), .C1(new_n739), .C2(new_n807), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n800), .B1(new_n827), .B2(new_n806), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n823), .B1(new_n828), .B2(new_n276), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n829), .A2(new_n803), .A3(new_n818), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n799), .B(new_n820), .C1(new_n822), .C2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT58), .B1(new_n829), .B2(new_n803), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n338), .ZN(new_n834));
  INV_X1    g633(.A(new_n803), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n819), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n833), .A2(KEYINPUT121), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n799), .B1(new_n837), .B2(new_n820), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n832), .A2(new_n838), .ZN(G1344gat));
  INV_X1    g638(.A(new_n802), .ZN(new_n840));
  INV_X1    g639(.A(new_n340), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n841), .A3(new_n561), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n804), .A2(new_n805), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n808), .B(KEYINPUT123), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n441), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n846), .B2(new_n805), .ZN(new_n847));
  OR3_X1    g646(.A1(new_n847), .A2(new_n562), .A3(new_n800), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n843), .B1(new_n848), .B2(G148gat), .ZN(new_n849));
  AOI211_X1 g648(.A(KEYINPUT59), .B(new_n841), .C1(new_n828), .C2(new_n561), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n842), .B1(new_n849), .B2(new_n850), .ZN(G1345gat));
  AOI21_X1  g650(.A(G155gat), .B1(new_n840), .B2(new_n584), .ZN(new_n852));
  INV_X1    g651(.A(new_n828), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n656), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n852), .B1(new_n854), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g654(.A(G162gat), .B1(new_n840), .B2(new_n653), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n828), .A2(G162gat), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n653), .ZN(G1347gat));
  AOI211_X1 g657(.A(new_n387), .B(new_n664), .C1(new_n739), .C2(new_n769), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n478), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n295), .A3(new_n276), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT124), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n859), .A2(new_n474), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n285), .B1(new_n864), .B2(new_n276), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n863), .A2(new_n865), .ZN(G1348gat));
  NAND3_X1  g665(.A1(new_n864), .A2(G176gat), .A3(new_n561), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n286), .B1(new_n860), .B2(new_n562), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n867), .A2(new_n868), .ZN(G1349gat));
  AOI21_X1  g668(.A(new_n279), .B1(new_n864), .B2(new_n657), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n584), .A2(new_n302), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n861), .B2(new_n871), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g672(.A(new_n280), .B1(new_n864), .B2(new_n653), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT61), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n874), .B1(KEYINPUT125), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(KEYINPUT125), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n280), .A3(new_n653), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1351gat));
  NOR3_X1   g679(.A1(new_n633), .A2(new_n387), .A3(new_n664), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n847), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G197gat), .B1(new_n883), .B2(new_n277), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n882), .A2(new_n804), .ZN(new_n885));
  INV_X1    g684(.A(G197gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n886), .A3(new_n276), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(G1352gat));
  INV_X1    g687(.A(G204gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n885), .A2(new_n889), .A3(new_n561), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n890), .B(KEYINPUT62), .Z(new_n891));
  NOR3_X1   g690(.A1(new_n847), .A2(new_n562), .A3(new_n882), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n889), .ZN(G1353gat));
  OAI211_X1 g692(.A(KEYINPUT63), .B(G211gat), .C1(new_n883), .C2(new_n639), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT63), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n847), .A2(new_n639), .A3(new_n882), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n393), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(KEYINPUT126), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n885), .A2(new_n393), .A3(new_n584), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n900), .B(new_n895), .C1(new_n896), .C2(new_n393), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(G1354gat));
  NOR3_X1   g701(.A1(new_n847), .A2(new_n616), .A3(new_n882), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n394), .ZN(new_n904));
  OAI22_X1  g703(.A1(new_n903), .A2(new_n394), .B1(new_n616), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


