

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U567 ( .A1(n544), .A2(n543), .ZN(G160) );
  NOR2_X1 U568 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U569 ( .A1(G651), .A2(n588), .ZN(n809) );
  BUF_X1 U570 ( .A(n662), .Z(n675) );
  NAND2_X1 U571 ( .A1(n610), .A2(n725), .ZN(n662) );
  OR2_X1 U572 ( .A1(n687), .A2(n686), .ZN(n714) );
  XNOR2_X1 U573 ( .A(KEYINPUT13), .B(KEYINPUT70), .ZN(n618) );
  XNOR2_X1 U574 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X1 U575 ( .A1(n588), .A2(n553), .ZN(n801) );
  OR2_X1 U576 ( .A1(n760), .A2(n759), .ZN(n775) );
  NOR2_X1 U577 ( .A1(G651), .A2(G543), .ZN(n802) );
  INV_X1 U578 ( .A(G2104), .ZN(n540) );
  NOR2_X4 U579 ( .A1(G2105), .A2(n540), .ZN(n1010) );
  NAND2_X1 U580 ( .A1(G101), .A2(n1010), .ZN(n535) );
  XNOR2_X1 U581 ( .A(n535), .B(KEYINPUT23), .ZN(n536) );
  XNOR2_X1 U582 ( .A(n536), .B(KEYINPUT65), .ZN(n539) );
  NOR2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n537) );
  XOR2_X2 U584 ( .A(KEYINPUT17), .B(n537), .Z(n1012) );
  NAND2_X1 U585 ( .A1(G137), .A2(n1012), .ZN(n538) );
  NAND2_X1 U586 ( .A1(n539), .A2(n538), .ZN(n544) );
  AND2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n1005) );
  NAND2_X1 U588 ( .A1(G113), .A2(n1005), .ZN(n542) );
  AND2_X1 U589 ( .A1(n540), .A2(G2105), .ZN(n1006) );
  NAND2_X1 U590 ( .A1(G125), .A2(n1006), .ZN(n541) );
  NAND2_X1 U591 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U592 ( .A1(G138), .A2(n1012), .ZN(n545) );
  XNOR2_X1 U593 ( .A(n545), .B(KEYINPUT84), .ZN(n552) );
  NAND2_X1 U594 ( .A1(G114), .A2(n1005), .ZN(n546) );
  XNOR2_X1 U595 ( .A(KEYINPUT83), .B(n546), .ZN(n550) );
  NAND2_X1 U596 ( .A1(G102), .A2(n1010), .ZN(n548) );
  NAND2_X1 U597 ( .A1(G126), .A2(n1006), .ZN(n547) );
  NAND2_X1 U598 ( .A1(n548), .A2(n547), .ZN(n549) );
  NOR2_X1 U599 ( .A1(n550), .A2(n549), .ZN(n551) );
  AND2_X1 U600 ( .A1(n552), .A2(n551), .ZN(G164) );
  XOR2_X1 U601 ( .A(KEYINPUT0), .B(G543), .Z(n588) );
  INV_X1 U602 ( .A(G651), .ZN(n553) );
  NAND2_X1 U603 ( .A1(G78), .A2(n801), .ZN(n556) );
  NOR2_X1 U604 ( .A1(G543), .A2(n553), .ZN(n554) );
  XOR2_X1 U605 ( .A(KEYINPUT1), .B(n554), .Z(n805) );
  NAND2_X1 U606 ( .A1(G65), .A2(n805), .ZN(n555) );
  NAND2_X1 U607 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U608 ( .A1(G91), .A2(n802), .ZN(n558) );
  NAND2_X1 U609 ( .A1(G53), .A2(n809), .ZN(n557) );
  NAND2_X1 U610 ( .A1(n558), .A2(n557), .ZN(n559) );
  OR2_X1 U611 ( .A1(n560), .A2(n559), .ZN(G299) );
  NAND2_X1 U612 ( .A1(G64), .A2(n805), .ZN(n562) );
  NAND2_X1 U613 ( .A1(G52), .A2(n809), .ZN(n561) );
  NAND2_X1 U614 ( .A1(n562), .A2(n561), .ZN(n567) );
  NAND2_X1 U615 ( .A1(G77), .A2(n801), .ZN(n564) );
  NAND2_X1 U616 ( .A1(G90), .A2(n802), .ZN(n563) );
  NAND2_X1 U617 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U618 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  NOR2_X1 U619 ( .A1(n567), .A2(n566), .ZN(G171) );
  INV_X1 U620 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U621 ( .A(KEYINPUT6), .B(KEYINPUT72), .ZN(n571) );
  NAND2_X1 U622 ( .A1(G63), .A2(n805), .ZN(n569) );
  NAND2_X1 U623 ( .A1(G51), .A2(n809), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U625 ( .A(n571), .B(n570), .ZN(n577) );
  NAND2_X1 U626 ( .A1(n802), .A2(G89), .ZN(n572) );
  XNOR2_X1 U627 ( .A(n572), .B(KEYINPUT4), .ZN(n574) );
  NAND2_X1 U628 ( .A1(G76), .A2(n801), .ZN(n573) );
  NAND2_X1 U629 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U630 ( .A(KEYINPUT5), .B(n575), .Z(n576) );
  NOR2_X1 U631 ( .A1(n577), .A2(n576), .ZN(n580) );
  XNOR2_X1 U632 ( .A(KEYINPUT74), .B(KEYINPUT7), .ZN(n578) );
  XNOR2_X1 U633 ( .A(n578), .B(KEYINPUT73), .ZN(n579) );
  XNOR2_X1 U634 ( .A(n580), .B(n579), .ZN(G168) );
  XOR2_X1 U635 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U636 ( .A1(G88), .A2(n802), .ZN(n582) );
  NAND2_X1 U637 ( .A1(G50), .A2(n809), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U639 ( .A1(G75), .A2(n801), .ZN(n584) );
  NAND2_X1 U640 ( .A1(G62), .A2(n805), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U642 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U643 ( .A(n587), .B(KEYINPUT77), .ZN(G303) );
  NAND2_X1 U644 ( .A1(G49), .A2(n809), .ZN(n590) );
  NAND2_X1 U645 ( .A1(G87), .A2(n588), .ZN(n589) );
  NAND2_X1 U646 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U647 ( .A1(n805), .A2(n591), .ZN(n593) );
  NAND2_X1 U648 ( .A1(G651), .A2(G74), .ZN(n592) );
  NAND2_X1 U649 ( .A1(n593), .A2(n592), .ZN(G288) );
  NAND2_X1 U650 ( .A1(G73), .A2(n801), .ZN(n594) );
  XNOR2_X1 U651 ( .A(n594), .B(KEYINPUT2), .ZN(n601) );
  NAND2_X1 U652 ( .A1(G61), .A2(n805), .ZN(n596) );
  NAND2_X1 U653 ( .A1(G48), .A2(n809), .ZN(n595) );
  NAND2_X1 U654 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U655 ( .A1(n802), .A2(G86), .ZN(n597) );
  XOR2_X1 U656 ( .A(KEYINPUT76), .B(n597), .Z(n598) );
  NOR2_X1 U657 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U658 ( .A1(n601), .A2(n600), .ZN(G305) );
  INV_X1 U659 ( .A(G303), .ZN(G166) );
  NAND2_X1 U660 ( .A1(G60), .A2(n805), .ZN(n603) );
  NAND2_X1 U661 ( .A1(G47), .A2(n809), .ZN(n602) );
  NAND2_X1 U662 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U663 ( .A1(G72), .A2(n801), .ZN(n604) );
  XOR2_X1 U664 ( .A(KEYINPUT66), .B(n604), .Z(n605) );
  NOR2_X1 U665 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U666 ( .A1(n802), .A2(G85), .ZN(n607) );
  NAND2_X1 U667 ( .A1(n608), .A2(n607), .ZN(G290) );
  NAND2_X1 U668 ( .A1(G40), .A2(G160), .ZN(n609) );
  XNOR2_X1 U669 ( .A(n609), .B(KEYINPUT86), .ZN(n726) );
  INV_X1 U670 ( .A(n726), .ZN(n610) );
  NOR2_X1 U671 ( .A1(G164), .A2(G1384), .ZN(n725) );
  INV_X1 U672 ( .A(n662), .ZN(n611) );
  AND2_X1 U673 ( .A1(n611), .A2(G1996), .ZN(n612) );
  XOR2_X1 U674 ( .A(n612), .B(KEYINPUT26), .Z(n626) );
  AND2_X1 U675 ( .A1(n662), .A2(G1341), .ZN(n624) );
  NAND2_X1 U676 ( .A1(n805), .A2(G56), .ZN(n613) );
  XOR2_X1 U677 ( .A(KEYINPUT14), .B(n613), .Z(n621) );
  NAND2_X1 U678 ( .A1(n801), .A2(G68), .ZN(n614) );
  XNOR2_X1 U679 ( .A(KEYINPUT69), .B(n614), .ZN(n617) );
  NAND2_X1 U680 ( .A1(n802), .A2(G81), .ZN(n615) );
  XOR2_X1 U681 ( .A(n615), .B(KEYINPUT12), .Z(n616) );
  NOR2_X1 U682 ( .A1(n617), .A2(n616), .ZN(n619) );
  NOR2_X1 U683 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U684 ( .A1(n809), .A2(G43), .ZN(n622) );
  NAND2_X1 U685 ( .A1(n623), .A2(n622), .ZN(n1028) );
  NOR2_X1 U686 ( .A1(n624), .A2(n1028), .ZN(n625) );
  AND2_X1 U687 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U688 ( .A(n627), .B(KEYINPUT64), .ZN(n641) );
  NAND2_X1 U689 ( .A1(G92), .A2(n802), .ZN(n629) );
  NAND2_X1 U690 ( .A1(G54), .A2(n809), .ZN(n628) );
  NAND2_X1 U691 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U692 ( .A1(G79), .A2(n801), .ZN(n631) );
  NAND2_X1 U693 ( .A1(G66), .A2(n805), .ZN(n630) );
  NAND2_X1 U694 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U695 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U696 ( .A(n634), .B(KEYINPUT15), .ZN(n930) );
  INV_X1 U697 ( .A(n930), .ZN(n1025) );
  AND2_X1 U698 ( .A1(n641), .A2(n1025), .ZN(n640) );
  NAND2_X1 U699 ( .A1(G2067), .A2(n611), .ZN(n635) );
  XNOR2_X1 U700 ( .A(KEYINPUT97), .B(n635), .ZN(n638) );
  NAND2_X1 U701 ( .A1(G1348), .A2(n675), .ZN(n636) );
  XOR2_X1 U702 ( .A(KEYINPUT96), .B(n636), .Z(n637) );
  NOR2_X1 U703 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U704 ( .A1(n640), .A2(n639), .ZN(n643) );
  NOR2_X1 U705 ( .A1(n1025), .A2(n641), .ZN(n642) );
  NOR2_X1 U706 ( .A1(n643), .A2(n642), .ZN(n649) );
  INV_X1 U707 ( .A(G2072), .ZN(n894) );
  NOR2_X1 U708 ( .A1(n675), .A2(n894), .ZN(n645) );
  XOR2_X1 U709 ( .A(KEYINPUT27), .B(KEYINPUT95), .Z(n644) );
  XNOR2_X1 U710 ( .A(n645), .B(n644), .ZN(n647) );
  NAND2_X1 U711 ( .A1(n675), .A2(G1956), .ZN(n646) );
  NAND2_X1 U712 ( .A1(n647), .A2(n646), .ZN(n651) );
  NOR2_X1 U713 ( .A1(n651), .A2(G299), .ZN(n648) );
  NOR2_X1 U714 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U715 ( .A(KEYINPUT98), .B(n650), .ZN(n654) );
  NAND2_X1 U716 ( .A1(G299), .A2(n651), .ZN(n652) );
  XOR2_X1 U717 ( .A(KEYINPUT28), .B(n652), .Z(n653) );
  XNOR2_X1 U718 ( .A(n655), .B(KEYINPUT29), .ZN(n661) );
  XOR2_X1 U719 ( .A(G2078), .B(KEYINPUT25), .Z(n900) );
  NOR2_X1 U720 ( .A1(n900), .A2(n675), .ZN(n656) );
  XOR2_X1 U721 ( .A(KEYINPUT93), .B(n656), .Z(n658) );
  NOR2_X1 U722 ( .A1(n611), .A2(G1961), .ZN(n657) );
  NOR2_X1 U723 ( .A1(n658), .A2(n657), .ZN(n668) );
  NOR2_X1 U724 ( .A1(n668), .A2(G301), .ZN(n659) );
  XOR2_X1 U725 ( .A(KEYINPUT94), .B(n659), .Z(n660) );
  NAND2_X1 U726 ( .A1(n661), .A2(n660), .ZN(n674) );
  NAND2_X1 U727 ( .A1(G8), .A2(n662), .ZN(n663) );
  XNOR2_X1 U728 ( .A(KEYINPUT92), .B(n663), .ZN(n719) );
  NOR2_X1 U729 ( .A1(n719), .A2(G1966), .ZN(n687) );
  NOR2_X1 U730 ( .A1(G2084), .A2(n675), .ZN(n683) );
  NOR2_X1 U731 ( .A1(n687), .A2(n683), .ZN(n664) );
  NAND2_X1 U732 ( .A1(G8), .A2(n664), .ZN(n665) );
  XNOR2_X1 U733 ( .A(KEYINPUT30), .B(n665), .ZN(n666) );
  NOR2_X1 U734 ( .A1(G168), .A2(n666), .ZN(n667) );
  XNOR2_X1 U735 ( .A(KEYINPUT99), .B(n667), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n668), .A2(G301), .ZN(n669) );
  XNOR2_X1 U737 ( .A(KEYINPUT100), .B(n669), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n672), .B(KEYINPUT31), .ZN(n673) );
  NAND2_X1 U740 ( .A1(n674), .A2(n673), .ZN(n685) );
  NAND2_X1 U741 ( .A1(n685), .A2(G286), .ZN(n680) );
  NOR2_X1 U742 ( .A1(G2090), .A2(n675), .ZN(n677) );
  NOR2_X1 U743 ( .A1(n719), .A2(G1971), .ZN(n676) );
  NOR2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U745 ( .A1(n678), .A2(G303), .ZN(n679) );
  NAND2_X1 U746 ( .A1(n680), .A2(n679), .ZN(n681) );
  NAND2_X1 U747 ( .A1(n681), .A2(G8), .ZN(n682) );
  XNOR2_X1 U748 ( .A(KEYINPUT32), .B(n682), .ZN(n716) );
  NAND2_X1 U749 ( .A1(G8), .A2(n683), .ZN(n684) );
  NAND2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  AND2_X1 U751 ( .A1(n714), .A2(KEYINPUT102), .ZN(n688) );
  NAND2_X1 U752 ( .A1(n716), .A2(n688), .ZN(n706) );
  INV_X1 U753 ( .A(KEYINPUT102), .ZN(n692) );
  NOR2_X1 U754 ( .A1(G1976), .A2(G288), .ZN(n922) );
  NOR2_X1 U755 ( .A1(G1971), .A2(G303), .ZN(n689) );
  NOR2_X1 U756 ( .A1(n922), .A2(n689), .ZN(n690) );
  XOR2_X1 U757 ( .A(KEYINPUT101), .B(n690), .Z(n691) );
  OR2_X1 U758 ( .A1(n692), .A2(n691), .ZN(n704) );
  NAND2_X1 U759 ( .A1(n922), .A2(KEYINPUT33), .ZN(n693) );
  AND2_X1 U760 ( .A1(n693), .A2(KEYINPUT102), .ZN(n696) );
  INV_X1 U761 ( .A(n922), .ZN(n694) );
  NOR2_X1 U762 ( .A1(KEYINPUT102), .A2(n694), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n696), .A2(n695), .ZN(n697) );
  INV_X1 U764 ( .A(n719), .ZN(n707) );
  AND2_X1 U765 ( .A1(n697), .A2(n707), .ZN(n698) );
  XNOR2_X1 U766 ( .A(G1981), .B(G305), .ZN(n924) );
  OR2_X1 U767 ( .A1(n698), .A2(n924), .ZN(n708) );
  INV_X1 U768 ( .A(n708), .ZN(n699) );
  NAND2_X1 U769 ( .A1(n699), .A2(KEYINPUT33), .ZN(n703) );
  NOR2_X1 U770 ( .A1(G1981), .A2(G305), .ZN(n700) );
  XNOR2_X1 U771 ( .A(n700), .B(KEYINPUT24), .ZN(n701) );
  NAND2_X1 U772 ( .A1(n701), .A2(n707), .ZN(n702) );
  AND2_X1 U773 ( .A1(n703), .A2(n702), .ZN(n711) );
  AND2_X1 U774 ( .A1(n704), .A2(n711), .ZN(n705) );
  AND2_X1 U775 ( .A1(n706), .A2(n705), .ZN(n713) );
  NAND2_X1 U776 ( .A1(G1976), .A2(G288), .ZN(n919) );
  NAND2_X1 U777 ( .A1(n707), .A2(n919), .ZN(n709) );
  OR2_X1 U778 ( .A1(n709), .A2(n708), .ZN(n710) );
  AND2_X1 U779 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U780 ( .A1(n713), .A2(n712), .ZN(n723) );
  AND2_X1 U781 ( .A1(n714), .A2(n719), .ZN(n715) );
  AND2_X1 U782 ( .A1(n716), .A2(n715), .ZN(n721) );
  NAND2_X1 U783 ( .A1(G166), .A2(G8), .ZN(n717) );
  NOR2_X1 U784 ( .A1(G2090), .A2(n717), .ZN(n718) );
  AND2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n720) );
  OR2_X1 U786 ( .A1(n721), .A2(n720), .ZN(n722) );
  NOR2_X1 U787 ( .A1(n723), .A2(n722), .ZN(n760) );
  XOR2_X1 U788 ( .A(G1986), .B(KEYINPUT85), .Z(n724) );
  XNOR2_X1 U789 ( .A(G290), .B(n724), .ZN(n918) );
  NOR2_X1 U790 ( .A1(n726), .A2(n725), .ZN(n772) );
  AND2_X1 U791 ( .A1(n918), .A2(n772), .ZN(n758) );
  NAND2_X1 U792 ( .A1(n1012), .A2(G140), .ZN(n727) );
  XOR2_X1 U793 ( .A(KEYINPUT87), .B(n727), .Z(n729) );
  NAND2_X1 U794 ( .A1(n1010), .A2(G104), .ZN(n728) );
  NAND2_X1 U795 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U796 ( .A(KEYINPUT34), .B(n730), .ZN(n735) );
  NAND2_X1 U797 ( .A1(G116), .A2(n1005), .ZN(n732) );
  NAND2_X1 U798 ( .A1(G128), .A2(n1006), .ZN(n731) );
  NAND2_X1 U799 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U800 ( .A(KEYINPUT35), .B(n733), .Z(n734) );
  NOR2_X1 U801 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U802 ( .A(KEYINPUT36), .B(n736), .ZN(n1021) );
  XNOR2_X1 U803 ( .A(G2067), .B(KEYINPUT37), .ZN(n769) );
  NOR2_X1 U804 ( .A1(n1021), .A2(n769), .ZN(n860) );
  NAND2_X1 U805 ( .A1(n860), .A2(n772), .ZN(n737) );
  XNOR2_X1 U806 ( .A(n737), .B(KEYINPUT88), .ZN(n767) );
  NAND2_X1 U807 ( .A1(G131), .A2(n1012), .ZN(n739) );
  NAND2_X1 U808 ( .A1(G119), .A2(n1006), .ZN(n738) );
  NAND2_X1 U809 ( .A1(n739), .A2(n738), .ZN(n743) );
  NAND2_X1 U810 ( .A1(G95), .A2(n1010), .ZN(n741) );
  NAND2_X1 U811 ( .A1(G107), .A2(n1005), .ZN(n740) );
  NAND2_X1 U812 ( .A1(n741), .A2(n740), .ZN(n742) );
  OR2_X1 U813 ( .A1(n743), .A2(n742), .ZN(n993) );
  NAND2_X1 U814 ( .A1(G1991), .A2(n993), .ZN(n744) );
  XNOR2_X1 U815 ( .A(n744), .B(KEYINPUT89), .ZN(n755) );
  XOR2_X1 U816 ( .A(KEYINPUT91), .B(KEYINPUT38), .Z(n746) );
  NAND2_X1 U817 ( .A1(G105), .A2(n1010), .ZN(n745) );
  XNOR2_X1 U818 ( .A(n746), .B(n745), .ZN(n753) );
  NAND2_X1 U819 ( .A1(G141), .A2(n1012), .ZN(n748) );
  NAND2_X1 U820 ( .A1(G129), .A2(n1006), .ZN(n747) );
  NAND2_X1 U821 ( .A1(n748), .A2(n747), .ZN(n751) );
  NAND2_X1 U822 ( .A1(n1005), .A2(G117), .ZN(n749) );
  XOR2_X1 U823 ( .A(KEYINPUT90), .B(n749), .Z(n750) );
  NOR2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U825 ( .A1(n753), .A2(n752), .ZN(n1002) );
  AND2_X1 U826 ( .A1(G1996), .A2(n1002), .ZN(n754) );
  NOR2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n857) );
  INV_X1 U828 ( .A(n857), .ZN(n756) );
  NAND2_X1 U829 ( .A1(n756), .A2(n772), .ZN(n761) );
  NAND2_X1 U830 ( .A1(n767), .A2(n761), .ZN(n757) );
  OR2_X1 U831 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U832 ( .A1(G1996), .A2(n1002), .ZN(n877) );
  INV_X1 U833 ( .A(n761), .ZN(n764) );
  NOR2_X1 U834 ( .A1(G1991), .A2(n993), .ZN(n861) );
  NOR2_X1 U835 ( .A1(G1986), .A2(G290), .ZN(n762) );
  NOR2_X1 U836 ( .A1(n861), .A2(n762), .ZN(n763) );
  NOR2_X1 U837 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U838 ( .A1(n877), .A2(n765), .ZN(n766) );
  XNOR2_X1 U839 ( .A(n766), .B(KEYINPUT39), .ZN(n768) );
  NAND2_X1 U840 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U841 ( .A1(n1021), .A2(n769), .ZN(n884) );
  NAND2_X1 U842 ( .A1(n770), .A2(n884), .ZN(n771) );
  XOR2_X1 U843 ( .A(KEYINPUT103), .B(n771), .Z(n773) );
  NAND2_X1 U844 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U845 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U846 ( .A(n776), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U847 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U848 ( .A(G57), .ZN(G237) );
  INV_X1 U849 ( .A(G132), .ZN(G219) );
  INV_X1 U850 ( .A(G82), .ZN(G220) );
  XOR2_X1 U851 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n778) );
  NAND2_X1 U852 ( .A1(G7), .A2(G661), .ZN(n777) );
  XNOR2_X1 U853 ( .A(n778), .B(n777), .ZN(G223) );
  XOR2_X1 U854 ( .A(G223), .B(KEYINPUT68), .Z(n842) );
  NAND2_X1 U855 ( .A1(n842), .A2(G567), .ZN(n779) );
  XOR2_X1 U856 ( .A(KEYINPUT11), .B(n779), .Z(G234) );
  INV_X1 U857 ( .A(n1028), .ZN(n780) );
  XOR2_X1 U858 ( .A(G860), .B(KEYINPUT71), .Z(n786) );
  NAND2_X1 U859 ( .A1(n780), .A2(n786), .ZN(G153) );
  NAND2_X1 U860 ( .A1(G868), .A2(G301), .ZN(n782) );
  INV_X1 U861 ( .A(G868), .ZN(n823) );
  NAND2_X1 U862 ( .A1(n930), .A2(n823), .ZN(n781) );
  NAND2_X1 U863 ( .A1(n782), .A2(n781), .ZN(G284) );
  NAND2_X1 U864 ( .A1(G868), .A2(G286), .ZN(n784) );
  NAND2_X1 U865 ( .A1(G299), .A2(n823), .ZN(n783) );
  NAND2_X1 U866 ( .A1(n784), .A2(n783), .ZN(G297) );
  INV_X1 U867 ( .A(G559), .ZN(n785) );
  NOR2_X1 U868 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U869 ( .A1(n930), .A2(n787), .ZN(n788) );
  XOR2_X1 U870 ( .A(KEYINPUT16), .B(n788), .Z(G148) );
  NOR2_X1 U871 ( .A1(G868), .A2(n1028), .ZN(n791) );
  NAND2_X1 U872 ( .A1(G868), .A2(n1025), .ZN(n789) );
  NOR2_X1 U873 ( .A1(G559), .A2(n789), .ZN(n790) );
  NOR2_X1 U874 ( .A1(n791), .A2(n790), .ZN(G282) );
  NAND2_X1 U875 ( .A1(G123), .A2(n1006), .ZN(n792) );
  XNOR2_X1 U876 ( .A(n792), .B(KEYINPUT18), .ZN(n794) );
  NAND2_X1 U877 ( .A1(n1005), .A2(G111), .ZN(n793) );
  NAND2_X1 U878 ( .A1(n794), .A2(n793), .ZN(n798) );
  NAND2_X1 U879 ( .A1(G99), .A2(n1010), .ZN(n796) );
  NAND2_X1 U880 ( .A1(G135), .A2(n1012), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U882 ( .A1(n798), .A2(n797), .ZN(n998) );
  XNOR2_X1 U883 ( .A(n998), .B(G2096), .ZN(n800) );
  INV_X1 U884 ( .A(G2100), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n800), .A2(n799), .ZN(G156) );
  NAND2_X1 U886 ( .A1(G80), .A2(n801), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G93), .A2(n802), .ZN(n803) );
  NAND2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n808) );
  NAND2_X1 U889 ( .A1(G67), .A2(n805), .ZN(n806) );
  XNOR2_X1 U890 ( .A(KEYINPUT75), .B(n806), .ZN(n807) );
  NOR2_X1 U891 ( .A1(n808), .A2(n807), .ZN(n811) );
  NAND2_X1 U892 ( .A1(n809), .A2(G55), .ZN(n810) );
  NAND2_X1 U893 ( .A1(n811), .A2(n810), .ZN(n824) );
  NAND2_X1 U894 ( .A1(G559), .A2(n1025), .ZN(n812) );
  XNOR2_X1 U895 ( .A(n812), .B(n1028), .ZN(n820) );
  NOR2_X1 U896 ( .A1(G860), .A2(n820), .ZN(n813) );
  XOR2_X1 U897 ( .A(n824), .B(n813), .Z(G145) );
  XNOR2_X1 U898 ( .A(G166), .B(G290), .ZN(n814) );
  XNOR2_X1 U899 ( .A(n814), .B(n824), .ZN(n815) );
  XNOR2_X1 U900 ( .A(KEYINPUT78), .B(n815), .ZN(n817) );
  XNOR2_X1 U901 ( .A(G288), .B(KEYINPUT19), .ZN(n816) );
  XNOR2_X1 U902 ( .A(n817), .B(n816), .ZN(n818) );
  XNOR2_X1 U903 ( .A(n818), .B(G305), .ZN(n819) );
  XNOR2_X1 U904 ( .A(n819), .B(G299), .ZN(n1024) );
  XNOR2_X1 U905 ( .A(n1024), .B(n820), .ZN(n821) );
  NAND2_X1 U906 ( .A1(n821), .A2(G868), .ZN(n822) );
  XOR2_X1 U907 ( .A(KEYINPUT79), .B(n822), .Z(n826) );
  NAND2_X1 U908 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U909 ( .A1(n826), .A2(n825), .ZN(G295) );
  NAND2_X1 U910 ( .A1(G2078), .A2(G2084), .ZN(n828) );
  XOR2_X1 U911 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n827) );
  XNOR2_X1 U912 ( .A(n828), .B(n827), .ZN(n829) );
  NAND2_X1 U913 ( .A1(n829), .A2(G2090), .ZN(n830) );
  XOR2_X1 U914 ( .A(KEYINPUT81), .B(n830), .Z(n831) );
  XNOR2_X1 U915 ( .A(KEYINPUT21), .B(n831), .ZN(n832) );
  NAND2_X1 U916 ( .A1(n832), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U917 ( .A(KEYINPUT82), .B(G44), .ZN(n833) );
  XNOR2_X1 U918 ( .A(n833), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U919 ( .A1(G220), .A2(G219), .ZN(n834) );
  XOR2_X1 U920 ( .A(KEYINPUT22), .B(n834), .Z(n835) );
  NOR2_X1 U921 ( .A1(G218), .A2(n835), .ZN(n836) );
  NAND2_X1 U922 ( .A1(G96), .A2(n836), .ZN(n973) );
  NAND2_X1 U923 ( .A1(n973), .A2(G2106), .ZN(n840) );
  NAND2_X1 U924 ( .A1(G69), .A2(G120), .ZN(n837) );
  NOR2_X1 U925 ( .A1(G237), .A2(n837), .ZN(n838) );
  NAND2_X1 U926 ( .A1(G108), .A2(n838), .ZN(n974) );
  NAND2_X1 U927 ( .A1(n974), .A2(G567), .ZN(n839) );
  NAND2_X1 U928 ( .A1(n840), .A2(n839), .ZN(n975) );
  NAND2_X1 U929 ( .A1(G483), .A2(G661), .ZN(n841) );
  NOR2_X1 U930 ( .A1(n975), .A2(n841), .ZN(n846) );
  NAND2_X1 U931 ( .A1(n846), .A2(G36), .ZN(G176) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n842), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U934 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n844) );
  XOR2_X1 U936 ( .A(KEYINPUT105), .B(n844), .Z(n845) );
  NAND2_X1 U937 ( .A1(n846), .A2(n845), .ZN(n847) );
  XNOR2_X1 U938 ( .A(KEYINPUT106), .B(n847), .ZN(G188) );
  NAND2_X1 U940 ( .A1(G124), .A2(n1006), .ZN(n848) );
  XOR2_X1 U941 ( .A(KEYINPUT107), .B(n848), .Z(n849) );
  XNOR2_X1 U942 ( .A(n849), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U943 ( .A1(G136), .A2(n1012), .ZN(n850) );
  NAND2_X1 U944 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U945 ( .A(KEYINPUT108), .B(n852), .ZN(n856) );
  NAND2_X1 U946 ( .A1(G100), .A2(n1010), .ZN(n854) );
  NAND2_X1 U947 ( .A1(G112), .A2(n1005), .ZN(n853) );
  NAND2_X1 U948 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U949 ( .A1(n856), .A2(n855), .ZN(G162) );
  XNOR2_X1 U950 ( .A(G160), .B(G2084), .ZN(n858) );
  NAND2_X1 U951 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U952 ( .A1(n860), .A2(n859), .ZN(n863) );
  NOR2_X1 U953 ( .A1(n861), .A2(n998), .ZN(n862) );
  NAND2_X1 U954 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U955 ( .A(KEYINPUT114), .B(n864), .ZN(n882) );
  XOR2_X1 U956 ( .A(G164), .B(G2078), .Z(n874) );
  NAND2_X1 U957 ( .A1(G115), .A2(n1005), .ZN(n866) );
  NAND2_X1 U958 ( .A1(G127), .A2(n1006), .ZN(n865) );
  NAND2_X1 U959 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U960 ( .A(n867), .B(KEYINPUT47), .ZN(n869) );
  NAND2_X1 U961 ( .A1(G139), .A2(n1012), .ZN(n868) );
  NAND2_X1 U962 ( .A1(n869), .A2(n868), .ZN(n872) );
  NAND2_X1 U963 ( .A1(n1010), .A2(G103), .ZN(n870) );
  XOR2_X1 U964 ( .A(KEYINPUT112), .B(n870), .Z(n871) );
  NOR2_X1 U965 ( .A1(n872), .A2(n871), .ZN(n996) );
  XNOR2_X1 U966 ( .A(n894), .B(n996), .ZN(n873) );
  NOR2_X1 U967 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U968 ( .A(KEYINPUT50), .B(n875), .ZN(n880) );
  XOR2_X1 U969 ( .A(G2090), .B(G162), .Z(n876) );
  NOR2_X1 U970 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U971 ( .A(KEYINPUT51), .B(n878), .Z(n879) );
  NAND2_X1 U972 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U973 ( .A1(n882), .A2(n881), .ZN(n883) );
  NAND2_X1 U974 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U975 ( .A(n885), .B(KEYINPUT115), .ZN(n886) );
  XNOR2_X1 U976 ( .A(KEYINPUT52), .B(n886), .ZN(n887) );
  INV_X1 U977 ( .A(KEYINPUT55), .ZN(n909) );
  NAND2_X1 U978 ( .A1(n887), .A2(n909), .ZN(n888) );
  NAND2_X1 U979 ( .A1(n888), .A2(G29), .ZN(n971) );
  XNOR2_X1 U980 ( .A(KEYINPUT54), .B(G34), .ZN(n889) );
  XNOR2_X1 U981 ( .A(n889), .B(KEYINPUT117), .ZN(n890) );
  XNOR2_X1 U982 ( .A(G2084), .B(n890), .ZN(n907) );
  XNOR2_X1 U983 ( .A(G2090), .B(G35), .ZN(n905) );
  XNOR2_X1 U984 ( .A(G2067), .B(G26), .ZN(n892) );
  XNOR2_X1 U985 ( .A(G1996), .B(G32), .ZN(n891) );
  NOR2_X1 U986 ( .A1(n892), .A2(n891), .ZN(n899) );
  XOR2_X1 U987 ( .A(G1991), .B(G25), .Z(n893) );
  NAND2_X1 U988 ( .A1(n893), .A2(G28), .ZN(n897) );
  XOR2_X1 U989 ( .A(KEYINPUT116), .B(n894), .Z(n895) );
  XNOR2_X1 U990 ( .A(G33), .B(n895), .ZN(n896) );
  NOR2_X1 U991 ( .A1(n897), .A2(n896), .ZN(n898) );
  NAND2_X1 U992 ( .A1(n899), .A2(n898), .ZN(n902) );
  XNOR2_X1 U993 ( .A(G27), .B(n900), .ZN(n901) );
  NOR2_X1 U994 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U995 ( .A(KEYINPUT53), .B(n903), .ZN(n904) );
  NOR2_X1 U996 ( .A1(n905), .A2(n904), .ZN(n906) );
  NAND2_X1 U997 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U998 ( .A(n909), .B(n908), .ZN(n911) );
  INV_X1 U999 ( .A(G29), .ZN(n910) );
  NAND2_X1 U1000 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1001 ( .A1(G11), .A2(n912), .ZN(n969) );
  INV_X1 U1002 ( .A(G16), .ZN(n965) );
  XOR2_X1 U1003 ( .A(KEYINPUT56), .B(KEYINPUT118), .Z(n913) );
  XNOR2_X1 U1004 ( .A(n965), .B(n913), .ZN(n939) );
  XNOR2_X1 U1005 ( .A(G1341), .B(n1028), .ZN(n916) );
  XOR2_X1 U1006 ( .A(G1971), .B(G166), .Z(n914) );
  XNOR2_X1 U1007 ( .A(KEYINPUT122), .B(n914), .ZN(n915) );
  NOR2_X1 U1008 ( .A1(n916), .A2(n915), .ZN(n937) );
  XNOR2_X1 U1009 ( .A(G1956), .B(G299), .ZN(n917) );
  NOR2_X1 U1010 ( .A1(n918), .A2(n917), .ZN(n920) );
  NAND2_X1 U1011 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1012 ( .A1(n922), .A2(n921), .ZN(n929) );
  XNOR2_X1 U1013 ( .A(G1966), .B(KEYINPUT119), .ZN(n923) );
  XNOR2_X1 U1014 ( .A(n923), .B(G168), .ZN(n925) );
  NOR2_X1 U1015 ( .A1(n925), .A2(n924), .ZN(n927) );
  XOR2_X1 U1016 ( .A(KEYINPUT57), .B(KEYINPUT120), .Z(n926) );
  XNOR2_X1 U1017 ( .A(n927), .B(n926), .ZN(n928) );
  NAND2_X1 U1018 ( .A1(n929), .A2(n928), .ZN(n935) );
  XNOR2_X1 U1019 ( .A(n930), .B(G1348), .ZN(n932) );
  XNOR2_X1 U1020 ( .A(G301), .B(G1961), .ZN(n931) );
  NOR2_X1 U1021 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1022 ( .A(n933), .B(KEYINPUT121), .ZN(n934) );
  NOR2_X1 U1023 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1024 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1025 ( .A1(n939), .A2(n938), .ZN(n967) );
  XOR2_X1 U1026 ( .A(G1986), .B(G24), .Z(n941) );
  XOR2_X1 U1027 ( .A(G1971), .B(G22), .Z(n940) );
  NAND2_X1 U1028 ( .A1(n941), .A2(n940), .ZN(n943) );
  XNOR2_X1 U1029 ( .A(G23), .B(G1976), .ZN(n942) );
  NOR2_X1 U1030 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1031 ( .A(KEYINPUT58), .B(n944), .Z(n962) );
  XNOR2_X1 U1032 ( .A(G1961), .B(G5), .ZN(n959) );
  XNOR2_X1 U1033 ( .A(G1981), .B(G6), .ZN(n946) );
  XNOR2_X1 U1034 ( .A(G19), .B(G1341), .ZN(n945) );
  NOR2_X1 U1035 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1036 ( .A(KEYINPUT123), .B(n947), .Z(n951) );
  XNOR2_X1 U1037 ( .A(KEYINPUT59), .B(G4), .ZN(n948) );
  XNOR2_X1 U1038 ( .A(n948), .B(KEYINPUT124), .ZN(n949) );
  XNOR2_X1 U1039 ( .A(G1348), .B(n949), .ZN(n950) );
  NAND2_X1 U1040 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1041 ( .A(G20), .B(G1956), .ZN(n952) );
  NOR2_X1 U1042 ( .A1(n953), .A2(n952), .ZN(n954) );
  XOR2_X1 U1043 ( .A(KEYINPUT60), .B(n954), .Z(n956) );
  XNOR2_X1 U1044 ( .A(G1966), .B(G21), .ZN(n955) );
  NOR2_X1 U1045 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1046 ( .A(KEYINPUT125), .B(n957), .ZN(n958) );
  NOR2_X1 U1047 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1048 ( .A(KEYINPUT126), .B(n960), .Z(n961) );
  NOR2_X1 U1049 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1050 ( .A(KEYINPUT61), .B(n963), .ZN(n964) );
  NAND2_X1 U1051 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1052 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1053 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1054 ( .A1(n971), .A2(n970), .ZN(n972) );
  XOR2_X1 U1055 ( .A(KEYINPUT62), .B(n972), .Z(G311) );
  XNOR2_X1 U1056 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1057 ( .A(G120), .ZN(G236) );
  INV_X1 U1058 ( .A(G96), .ZN(G221) );
  INV_X1 U1059 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1060 ( .A1(n974), .A2(n973), .ZN(G325) );
  INV_X1 U1061 ( .A(G325), .ZN(G261) );
  INV_X1 U1062 ( .A(n975), .ZN(G319) );
  XOR2_X1 U1063 ( .A(G2100), .B(G2096), .Z(n977) );
  XNOR2_X1 U1064 ( .A(G2067), .B(G2090), .ZN(n976) );
  XNOR2_X1 U1065 ( .A(n977), .B(n976), .ZN(n981) );
  XOR2_X1 U1066 ( .A(G2678), .B(KEYINPUT42), .Z(n979) );
  XNOR2_X1 U1067 ( .A(G2072), .B(KEYINPUT43), .ZN(n978) );
  XNOR2_X1 U1068 ( .A(n979), .B(n978), .ZN(n980) );
  XOR2_X1 U1069 ( .A(n981), .B(n980), .Z(n983) );
  XNOR2_X1 U1070 ( .A(G2078), .B(G2084), .ZN(n982) );
  XNOR2_X1 U1071 ( .A(n983), .B(n982), .ZN(G227) );
  XOR2_X1 U1072 ( .A(G1971), .B(G1956), .Z(n985) );
  XNOR2_X1 U1073 ( .A(G1986), .B(G1966), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(n985), .B(n984), .ZN(n986) );
  XOR2_X1 U1075 ( .A(n986), .B(KEYINPUT41), .Z(n988) );
  XNOR2_X1 U1076 ( .A(G1991), .B(G1961), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(n988), .B(n987), .ZN(n992) );
  XOR2_X1 U1078 ( .A(G2474), .B(G1976), .Z(n990) );
  XNOR2_X1 U1079 ( .A(G1996), .B(G1981), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n990), .B(n989), .ZN(n991) );
  XNOR2_X1 U1081 ( .A(n992), .B(n991), .ZN(G229) );
  XNOR2_X1 U1082 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(n993), .B(KEYINPUT46), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(n995), .B(n994), .ZN(n997) );
  XOR2_X1 U1085 ( .A(n997), .B(n996), .Z(n1000) );
  XNOR2_X1 U1086 ( .A(G164), .B(n998), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(n1000), .B(n999), .ZN(n1001) );
  XOR2_X1 U1088 ( .A(n1001), .B(G162), .Z(n1004) );
  XOR2_X1 U1089 ( .A(G160), .B(n1002), .Z(n1003) );
  XNOR2_X1 U1090 ( .A(n1004), .B(n1003), .ZN(n1020) );
  NAND2_X1 U1091 ( .A1(G118), .A2(n1005), .ZN(n1008) );
  NAND2_X1 U1092 ( .A1(G130), .A2(n1006), .ZN(n1007) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1094 ( .A(KEYINPUT109), .B(n1009), .Z(n1018) );
  NAND2_X1 U1095 ( .A1(n1010), .A2(G106), .ZN(n1011) );
  XNOR2_X1 U1096 ( .A(KEYINPUT110), .B(n1011), .ZN(n1015) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(G142), .ZN(n1013) );
  XOR2_X1 U1098 ( .A(KEYINPUT111), .B(n1013), .Z(n1014) );
  NAND2_X1 U1099 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1100 ( .A(n1016), .B(KEYINPUT45), .Z(n1017) );
  NOR2_X1 U1101 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1102 ( .A(n1020), .B(n1019), .Z(n1022) );
  XOR2_X1 U1103 ( .A(n1022), .B(n1021), .Z(n1023) );
  NOR2_X1 U1104 ( .A1(G37), .A2(n1023), .ZN(G395) );
  XNOR2_X1 U1105 ( .A(G286), .B(n1024), .ZN(n1027) );
  XNOR2_X1 U1106 ( .A(n1025), .B(G171), .ZN(n1026) );
  XNOR2_X1 U1107 ( .A(n1027), .B(n1026), .ZN(n1029) );
  XOR2_X1 U1108 ( .A(n1029), .B(n1028), .Z(n1030) );
  NOR2_X1 U1109 ( .A1(G37), .A2(n1030), .ZN(G397) );
  XOR2_X1 U1110 ( .A(G2451), .B(G2443), .Z(n1032) );
  XNOR2_X1 U1111 ( .A(G1348), .B(G2454), .ZN(n1031) );
  XNOR2_X1 U1112 ( .A(n1032), .B(n1031), .ZN(n1033) );
  XOR2_X1 U1113 ( .A(n1033), .B(G2446), .Z(n1035) );
  XNOR2_X1 U1114 ( .A(G2430), .B(G2438), .ZN(n1034) );
  XNOR2_X1 U1115 ( .A(n1035), .B(n1034), .ZN(n1039) );
  XOR2_X1 U1116 ( .A(G2427), .B(G2435), .Z(n1037) );
  XNOR2_X1 U1117 ( .A(G1341), .B(KEYINPUT104), .ZN(n1036) );
  XNOR2_X1 U1118 ( .A(n1037), .B(n1036), .ZN(n1038) );
  XOR2_X1 U1119 ( .A(n1039), .B(n1038), .Z(n1040) );
  NAND2_X1 U1120 ( .A1(G14), .A2(n1040), .ZN(n1046) );
  NAND2_X1 U1121 ( .A1(G319), .A2(n1046), .ZN(n1043) );
  NOR2_X1 U1122 ( .A1(G227), .A2(G229), .ZN(n1041) );
  XNOR2_X1 U1123 ( .A(KEYINPUT49), .B(n1041), .ZN(n1042) );
  NOR2_X1 U1124 ( .A1(n1043), .A2(n1042), .ZN(n1045) );
  NOR2_X1 U1125 ( .A1(G395), .A2(G397), .ZN(n1044) );
  NAND2_X1 U1126 ( .A1(n1045), .A2(n1044), .ZN(G225) );
  INV_X1 U1127 ( .A(G225), .ZN(G308) );
  INV_X1 U1128 ( .A(G108), .ZN(G238) );
  INV_X1 U1129 ( .A(n1046), .ZN(G401) );
endmodule

