//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(KEYINPUT1), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n204), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(new_n207), .A3(new_n202), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT70), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(KEYINPUT70), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT27), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(G183gat), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT66), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT66), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G190gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n218), .A2(new_n222), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n218), .A2(KEYINPUT67), .A3(new_n222), .A4(new_n224), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n219), .A2(new_n220), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(new_n223), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  AND2_X1   g033(.A1(KEYINPUT68), .A2(KEYINPUT26), .ZN(new_n235));
  NOR2_X1   g034(.A1(KEYINPUT68), .A2(KEYINPUT26), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT69), .ZN(new_n238));
  INV_X1    g037(.A(G169gat), .ZN(new_n239));
  INV_X1    g038(.A(G176gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n234), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n241), .B1(KEYINPUT26), .B2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n233), .B1(new_n238), .B2(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n232), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT24), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n233), .A2(new_n246), .B1(G169gat), .B2(G176gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT23), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n248), .A2(new_n239), .A3(new_n240), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G183gat), .B(G190gat), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n247), .B(new_n251), .C1(new_n246), .C2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT64), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(KEYINPUT65), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT25), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n258), .B1(new_n253), .B2(new_n254), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n212), .B(new_n213), .C1(new_n245), .C2(new_n262), .ZN(new_n263));
  AOI211_X1 g062(.A(new_n258), .B(KEYINPUT25), .C1(new_n253), .C2(new_n254), .ZN(new_n264));
  INV_X1    g063(.A(new_n261), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n256), .B1(new_n253), .B2(new_n258), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n232), .A2(new_n244), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n267), .A2(new_n211), .A3(new_n210), .A4(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G227gat), .ZN(new_n270));
  INV_X1    g069(.A(G233gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n263), .A2(new_n269), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n263), .A2(new_n269), .A3(KEYINPUT71), .A4(new_n272), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT32), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT34), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n269), .ZN(new_n280));
  INV_X1    g079(.A(new_n272), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI211_X1 g081(.A(KEYINPUT34), .B(new_n272), .C1(new_n263), .C2(new_n269), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G15gat), .B(G43gat), .Z(new_n286));
  XNOR2_X1  g085(.A(G71gat), .B(G99gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT33), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n277), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n280), .A2(new_n281), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT34), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n280), .A2(new_n279), .A3(new_n281), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n296), .B1(new_n275), .B2(new_n276), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n285), .A2(new_n291), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n291), .B1(new_n285), .B2(new_n298), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G8gat), .B(G36gat), .Z(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(KEYINPUT76), .ZN(new_n303));
  XNOR2_X1  g102(.A(G64gat), .B(G92gat), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n303), .B(new_n304), .Z(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G211gat), .B(G218gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G218gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT73), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G218gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT22), .B1(new_n313), .B2(G211gat), .ZN(new_n314));
  XOR2_X1   g113(.A(G197gat), .B(G204gat), .Z(new_n315));
  OAI21_X1  g114(.A(new_n308), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT22), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT73), .B(G218gat), .ZN(new_n318));
  INV_X1    g117(.A(G211gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n315), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n307), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n245), .A2(new_n262), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT74), .B1(new_n267), .B2(new_n268), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n267), .A2(new_n268), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n326), .A2(KEYINPUT29), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n324), .B1(new_n330), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n327), .B1(new_n245), .B2(new_n262), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n267), .A2(KEYINPUT74), .A3(new_n268), .ZN(new_n336));
  XOR2_X1   g135(.A(KEYINPUT75), .B(KEYINPUT29), .Z(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(new_n326), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n335), .A2(new_n336), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n267), .A2(new_n326), .A3(new_n268), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n340), .A2(new_n324), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n306), .B1(new_n334), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT77), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n325), .B1(new_n335), .B2(new_n336), .ZN(new_n345));
  INV_X1    g144(.A(new_n333), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n323), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n340), .A2(new_n324), .A3(new_n341), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n347), .A2(KEYINPUT30), .A3(new_n348), .A4(new_n305), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n350), .B(new_n306), .C1(new_n334), .C2(new_n342), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n348), .A3(new_n305), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT30), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n344), .A2(new_n349), .A3(new_n351), .A4(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n357));
  XNOR2_X1  g156(.A(G78gat), .B(G106gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT31), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(G50gat), .ZN(new_n360));
  OR3_X1    g159(.A1(KEYINPUT80), .A2(G155gat), .A3(G162gat), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n363), .B1(G155gat), .B2(G162gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(KEYINPUT79), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n361), .B(new_n362), .C1(new_n364), .C2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n365), .B(KEYINPUT79), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n370), .A2(KEYINPUT81), .A3(new_n362), .A4(new_n361), .ZN(new_n371));
  INV_X1    g170(.A(G141gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G148gat), .ZN(new_n373));
  INV_X1    g172(.A(G148gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G141gat), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n373), .A2(new_n375), .B1(KEYINPUT2), .B2(new_n365), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n369), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  OR2_X1    g177(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(KEYINPUT82), .A2(G148gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(G141gat), .A3(new_n380), .ZN(new_n381));
  OR3_X1    g180(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n381), .A2(new_n373), .B1(new_n382), .B2(new_n365), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n316), .B2(new_n322), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI211_X1 g188(.A(KEYINPUT84), .B(KEYINPUT29), .C1(new_n316), .C2(new_n322), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n376), .B1(new_n367), .B2(new_n368), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n383), .B1(new_n393), .B2(new_n371), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n338), .B1(new_n394), .B2(new_n386), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n392), .B1(new_n395), .B2(new_n323), .ZN(new_n396));
  INV_X1    g195(.A(G228gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(new_n271), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n378), .A2(new_n386), .A3(new_n384), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n337), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(KEYINPUT85), .A3(new_n324), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n391), .A2(new_n396), .A3(new_n398), .A4(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G22gat), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n395), .A2(new_n323), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n323), .A2(new_n337), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n394), .B1(new_n405), .B2(new_n386), .ZN(new_n406));
  OAI22_X1  g205(.A1(new_n404), .A2(new_n406), .B1(new_n397), .B2(new_n271), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n402), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n403), .B1(new_n402), .B2(new_n407), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n357), .B(new_n360), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n402), .A2(new_n407), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(G22gat), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n402), .A2(new_n403), .A3(new_n407), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n360), .B1(new_n415), .B2(new_n357), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(KEYINPUT86), .A3(new_n414), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n411), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G1gat), .B(G29gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT0), .ZN(new_n420));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n385), .A2(new_n210), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n378), .A2(new_n209), .A3(new_n384), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n424), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n394), .A2(KEYINPUT4), .A3(new_n209), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n385), .A2(KEYINPUT83), .A3(KEYINPUT3), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(new_n394), .B2(new_n386), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n399), .A2(new_n210), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n434), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n430), .B1(new_n441), .B2(new_n428), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n439), .B1(new_n437), .B2(new_n435), .ZN(new_n443));
  NOR4_X1   g242(.A1(new_n443), .A2(new_n434), .A3(new_n424), .A4(new_n429), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n423), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n438), .A2(new_n440), .ZN(new_n447));
  INV_X1    g246(.A(new_n434), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n447), .A2(KEYINPUT5), .A3(new_n448), .A4(new_n428), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n422), .B(KEYINPUT87), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n443), .A2(new_n429), .A3(new_n434), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n449), .B(new_n451), .C1(new_n452), .C2(new_n430), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n445), .A2(new_n446), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n442), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n455), .A2(KEYINPUT6), .A3(new_n422), .A4(new_n449), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT35), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n301), .A2(new_n356), .A3(new_n418), .A4(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT78), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n351), .A2(new_n349), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n347), .A2(new_n348), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n350), .B1(new_n461), .B2(new_n306), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n459), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n344), .A2(KEYINPUT78), .A3(new_n349), .A4(new_n351), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n449), .B(new_n422), .C1(new_n452), .C2(new_n430), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n445), .A2(new_n446), .A3(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n466), .A2(new_n456), .B1(new_n353), .B2(new_n352), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n291), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n278), .A2(new_n284), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n295), .A2(new_n297), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n415), .A2(new_n357), .ZN(new_n473));
  INV_X1    g272(.A(new_n360), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n417), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n285), .A2(new_n291), .A3(new_n298), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n472), .A2(new_n410), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT92), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n418), .A2(KEYINPUT92), .A3(new_n476), .A4(new_n472), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n468), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT35), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n458), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n418), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT72), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(KEYINPUT36), .C1(new_n299), .C2(new_n300), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(KEYINPUT36), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n486), .A2(KEYINPUT36), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n472), .A2(new_n488), .A3(new_n489), .A4(new_n476), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT40), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n447), .A2(new_n448), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT39), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(new_n429), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n450), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT39), .B1(new_n427), .B2(new_n429), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n497), .B1(new_n493), .B2(new_n429), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n492), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n498), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n500), .A2(KEYINPUT40), .A3(new_n450), .A4(new_n495), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n499), .A2(new_n501), .A3(new_n453), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n355), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT88), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n355), .A2(new_n502), .A3(KEYINPUT88), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n506), .A3(new_n418), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT91), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT38), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n340), .A2(new_n323), .A3(new_n341), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n510), .A2(KEYINPUT37), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n324), .B1(new_n345), .B2(new_n346), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT89), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g312(.A1(new_n512), .A2(KEYINPUT89), .A3(KEYINPUT37), .A4(new_n510), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n509), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n347), .A2(new_n517), .A3(new_n348), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n305), .B1(new_n518), .B2(KEYINPUT90), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT90), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n347), .A2(new_n520), .A3(new_n517), .A4(new_n348), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n508), .B1(new_n516), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n454), .A2(new_n456), .A3(new_n352), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(KEYINPUT90), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n461), .A2(KEYINPUT37), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n525), .A2(new_n526), .A3(new_n521), .A4(new_n306), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n524), .B1(new_n527), .B2(KEYINPUT38), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n512), .A2(KEYINPUT37), .A3(new_n510), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT89), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(KEYINPUT38), .B1(new_n531), .B2(new_n514), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n532), .A2(KEYINPUT91), .A3(new_n521), .A4(new_n519), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n523), .A2(new_n528), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n485), .B(new_n491), .C1(new_n507), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n483), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G183gat), .B(G211gat), .Z(new_n537));
  AOI21_X1  g336(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n538), .A2(KEYINPUT98), .ZN(new_n539));
  XOR2_X1   g338(.A(G57gat), .B(G64gat), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(KEYINPUT98), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G71gat), .B(G78gat), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n539), .A2(new_n540), .A3(new_n543), .A4(new_n541), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT21), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G127gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n550), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n549), .B(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(G127gat), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n537), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(G127gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n551), .A2(new_n552), .ZN(new_n559));
  INV_X1    g358(.A(new_n537), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n563));
  INV_X1    g362(.A(G155gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G8gat), .ZN(new_n566));
  INV_X1    g365(.A(G15gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n403), .ZN(new_n568));
  NAND2_X1  g367(.A1(G15gat), .A2(G22gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G1gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(KEYINPUT16), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(G1gat), .A3(new_n569), .ZN(new_n573));
  AOI211_X1 g372(.A(KEYINPUT94), .B(new_n566), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n566), .A2(KEYINPUT94), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n566), .A2(KEYINPUT94), .ZN(new_n576));
  AND4_X1   g375(.A1(new_n575), .A2(new_n572), .A3(new_n576), .A4(new_n573), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n579), .B1(new_n548), .B2(new_n547), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT99), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n580), .A2(KEYINPUT99), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n565), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n580), .A2(KEYINPUT99), .ZN(new_n585));
  INV_X1    g384(.A(new_n565), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n585), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n562), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n557), .A2(new_n584), .A3(new_n561), .A4(new_n587), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G99gat), .B(G106gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(KEYINPUT103), .A2(KEYINPUT7), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G99gat), .ZN(new_n598));
  INV_X1    g397(.A(G106gat), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT8), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(G85gat), .B(G92gat), .C1(KEYINPUT103), .C2(KEYINPUT7), .ZN(new_n602));
  AND2_X1   g401(.A1(KEYINPUT103), .A2(KEYINPUT7), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n593), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n606), .A2(new_n597), .A3(new_n592), .A4(new_n600), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(G29gat), .A2(G36gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT14), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT14), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n611), .B1(G29gat), .B2(G36gat), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OR2_X1    g412(.A1(KEYINPUT93), .A2(G29gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(KEYINPUT93), .A2(G29gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(G36gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n617), .A3(KEYINPUT15), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT15), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n610), .A2(new_n612), .ZN(new_n620));
  INV_X1    g419(.A(G36gat), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n621), .B1(new_n614), .B2(new_n615), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n619), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G43gat), .B(G50gat), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT17), .ZN(new_n626));
  INV_X1    g425(.A(new_n624), .ZN(new_n627));
  NAND4_X1  g426(.A1(new_n613), .A2(new_n617), .A3(KEYINPUT15), .A4(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n626), .B1(new_n625), .B2(new_n628), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n608), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT100), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT41), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n625), .A2(new_n628), .ZN(new_n636));
  INV_X1    g435(.A(new_n608), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n635), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n631), .A2(new_n229), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n229), .B1(new_n631), .B2(new_n638), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n309), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n641), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(G218gat), .A3(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n633), .A2(new_n634), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT101), .ZN(new_n646));
  INV_X1    g445(.A(G134gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G162gat), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n642), .A2(new_n644), .A3(KEYINPUT102), .A4(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n644), .A3(KEYINPUT102), .ZN(new_n651));
  INV_X1    g450(.A(new_n649), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n591), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n579), .B1(new_n629), .B2(new_n630), .ZN(new_n656));
  NAND2_X1  g455(.A1(G229gat), .A2(G233gat), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT95), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n578), .A2(new_n658), .A3(new_n636), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n578), .B2(new_n636), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n656), .B(new_n657), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT18), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n664), .A2(KEYINPUT18), .A3(new_n657), .A4(new_n656), .ZN(new_n665));
  OAI22_X1  g464(.A1(new_n659), .A2(new_n660), .B1(new_n578), .B2(new_n636), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n657), .B(KEYINPUT13), .Z(new_n667));
  AND3_X1   g466(.A1(new_n666), .A2(KEYINPUT96), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT96), .B1(new_n666), .B2(new_n667), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n663), .B(new_n665), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(G113gat), .B(G141gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G197gat), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT11), .B(G169gat), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(KEYINPUT12), .Z(new_n675));
  NAND2_X1  g474(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n666), .A2(new_n667), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT96), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n666), .A2(KEYINPUT96), .A3(new_n667), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n675), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n663), .A4(new_n665), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n676), .A2(new_n683), .A3(KEYINPUT97), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT97), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n685), .A3(new_n675), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n547), .A2(new_n608), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n545), .A2(new_n605), .A3(new_n546), .A4(new_n607), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT104), .B(KEYINPUT10), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n637), .A2(KEYINPUT10), .A3(new_n545), .A4(new_n546), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n688), .A2(KEYINPUT105), .A3(new_n689), .A4(new_n690), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(G230gat), .A2(G233gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n688), .A2(new_n689), .ZN(new_n699));
  INV_X1    g498(.A(new_n697), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(G120gat), .B(G148gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(G176gat), .B(G204gat), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n703), .B(new_n704), .Z(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n698), .A2(new_n701), .A3(new_n705), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n655), .A2(new_n687), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n536), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n466), .A2(new_n456), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(new_n571), .ZN(G1324gat));
  AND2_X1   g513(.A1(new_n536), .A2(new_n710), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT16), .B(G8gat), .Z(new_n716));
  NAND3_X1  g515(.A1(new_n715), .A2(new_n355), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G8gat), .B1(new_n711), .B2(new_n356), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n718), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT106), .Z(G1325gat));
  NAND3_X1  g522(.A1(new_n715), .A2(new_n567), .A3(new_n301), .ZN(new_n724));
  OAI21_X1  g523(.A(G15gat), .B1(new_n711), .B2(new_n491), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(G1326gat));
  NAND2_X1  g525(.A1(new_n715), .A2(new_n484), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT107), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT43), .B(G22gat), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1327gat));
  NAND2_X1  g529(.A1(new_n653), .A2(new_n650), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n483), .B2(new_n535), .ZN(new_n732));
  INV_X1    g531(.A(new_n591), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n687), .A2(new_n733), .A3(new_n709), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n735), .A2(new_n712), .A3(new_n616), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT45), .Z(new_n737));
  INV_X1    g536(.A(new_n731), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT44), .B1(new_n536), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n740));
  AOI211_X1 g539(.A(new_n740), .B(new_n731), .C1(new_n483), .C2(new_n535), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n734), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n616), .B1(new_n743), .B2(new_n712), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n737), .A2(new_n744), .ZN(G1328gat));
  OAI21_X1  g544(.A(G36gat), .B1(new_n743), .B2(new_n356), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n747));
  AOI21_X1  g546(.A(G36gat), .B1(new_n747), .B2(KEYINPUT46), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n355), .A3(new_n734), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n747), .A2(KEYINPUT46), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n746), .A2(new_n751), .ZN(G1329gat));
  INV_X1    g551(.A(new_n491), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G43gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n472), .A2(new_n476), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n735), .A2(new_n755), .ZN(new_n756));
  OAI22_X1  g555(.A1(new_n743), .A2(new_n754), .B1(G43gat), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g557(.A(G50gat), .B1(new_n743), .B2(new_n418), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n735), .A2(G50gat), .A3(new_n418), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT48), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n761), .B(new_n763), .ZN(G1331gat));
  NAND3_X1  g563(.A1(new_n687), .A2(new_n654), .A3(new_n709), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT110), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n483), .B2(new_n535), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n712), .B(KEYINPUT111), .Z(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g569(.A(new_n356), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(KEYINPUT112), .ZN(new_n773));
  NOR2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1333gat));
  NAND2_X1  g574(.A1(new_n767), .A2(new_n753), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n755), .A2(G71gat), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n776), .A2(G71gat), .B1(new_n767), .B2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g578(.A1(new_n767), .A2(new_n484), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g580(.A1(new_n687), .A2(new_n591), .ZN(new_n782));
  INV_X1    g581(.A(new_n709), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n739), .A2(new_n741), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n712), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G85gat), .ZN(new_n789));
  INV_X1    g588(.A(new_n782), .ZN(new_n790));
  XNOR2_X1  g589(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n536), .A2(new_n738), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n731), .B(new_n782), .C1(new_n483), .C2(new_n535), .ZN(new_n793));
  AND2_X1   g592(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OR3_X1    g595(.A1(new_n712), .A2(G85gat), .A3(new_n783), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n789), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n789), .B(KEYINPUT114), .C1(new_n796), .C2(new_n797), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(G1336gat));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n355), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G92gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n803), .B1(new_n805), .B2(KEYINPUT115), .ZN(new_n806));
  OR3_X1    g605(.A1(new_n356), .A2(G92gat), .A3(new_n783), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n796), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OAI221_X1 g608(.A(new_n805), .B1(KEYINPUT115), .B2(new_n803), .C1(new_n796), .C2(new_n807), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(G1337gat));
  NAND2_X1  g610(.A1(new_n786), .A2(new_n753), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n598), .B1(new_n812), .B2(KEYINPUT116), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(KEYINPUT116), .B2(new_n812), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n301), .A2(new_n598), .A3(new_n709), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n796), .B2(new_n815), .ZN(G1338gat));
  AOI21_X1  g615(.A(new_n599), .B1(new_n786), .B2(new_n484), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n418), .A2(G106gat), .A3(new_n783), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n795), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g618(.A(KEYINPUT117), .B(KEYINPUT53), .C1(new_n817), .C2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821));
  INV_X1    g620(.A(new_n458), .ZN(new_n822));
  INV_X1    g621(.A(new_n468), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT92), .B1(new_n301), .B2(new_n418), .ZN(new_n824));
  AND4_X1   g623(.A1(KEYINPUT92), .A2(new_n418), .A3(new_n476), .A4(new_n472), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n822), .B1(new_n826), .B2(KEYINPUT35), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n485), .A2(new_n487), .A3(new_n490), .ZN(new_n828));
  INV_X1    g627(.A(new_n534), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n505), .A2(new_n506), .A3(new_n418), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n738), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n740), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n732), .A2(KEYINPUT44), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n833), .A2(new_n484), .A3(new_n834), .A4(new_n784), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n835), .A2(G106gat), .B1(new_n795), .B2(new_n818), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n821), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n742), .A2(KEYINPUT118), .A3(new_n484), .A4(new_n784), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n842), .A3(G106gat), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT53), .B1(new_n795), .B2(new_n818), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n843), .A2(KEYINPUT119), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT119), .B1(new_n843), .B2(new_n844), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n839), .B1(new_n845), .B2(new_n846), .ZN(G1339gat));
  NAND3_X1  g646(.A1(new_n687), .A2(new_n654), .A3(new_n783), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT120), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n687), .A2(new_n654), .A3(new_n850), .A4(new_n783), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n693), .A2(new_n700), .A3(new_n694), .A4(new_n695), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n698), .A2(KEYINPUT54), .A3(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n696), .A2(new_n855), .A3(new_n697), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n854), .A2(KEYINPUT55), .A3(new_n706), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n708), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT121), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n857), .A2(new_n860), .A3(new_n708), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n854), .A2(new_n706), .A3(new_n856), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n859), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n666), .A2(new_n667), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n657), .B1(new_n664), .B2(new_n656), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n674), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n653), .A2(new_n683), .A3(new_n650), .A4(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n683), .A2(new_n709), .A3(new_n869), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n872), .B1(new_n865), .B2(new_n687), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n871), .B1(new_n873), .B2(new_n731), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n852), .B1(new_n874), .B2(new_n733), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n768), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n824), .A2(new_n825), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n355), .A3(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n687), .ZN(new_n879));
  AOI21_X1  g678(.A(G113gat), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n875), .A2(new_n418), .A3(new_n301), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n355), .A2(new_n712), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n879), .A2(G113gat), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(G1340gat));
  AOI21_X1  g684(.A(G120gat), .B1(new_n878), .B2(new_n709), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n709), .A2(G120gat), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n883), .B2(new_n887), .ZN(G1341gat));
  NAND3_X1  g687(.A1(new_n878), .A2(new_n552), .A3(new_n733), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n883), .A2(new_n733), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n552), .ZN(G1342gat));
  AND2_X1   g690(.A1(new_n883), .A2(new_n738), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n647), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n647), .A3(new_n738), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n893), .B1(KEYINPUT56), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(KEYINPUT56), .B2(new_n894), .ZN(G1343gat));
  INV_X1    g695(.A(new_n876), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n753), .A2(new_n355), .A3(new_n418), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n372), .B1(new_n899), .B2(new_n687), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n491), .A2(new_n882), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n875), .A2(new_n484), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n418), .A2(new_n903), .ZN(new_n905));
  INV_X1    g704(.A(new_n858), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n684), .A2(new_n906), .A3(new_n686), .A4(new_n864), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n738), .B1(new_n907), .B2(new_n872), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n591), .B1(new_n908), .B2(new_n871), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n852), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n905), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n901), .B1(new_n904), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n879), .A2(G141gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n900), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT58), .Z(G1344gat));
  NAND2_X1  g717(.A1(new_n379), .A2(new_n380), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n914), .B2(new_n709), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n875), .A2(new_n923), .A3(new_n905), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(new_n875), .B2(new_n905), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n848), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n926), .B2(new_n484), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n491), .A2(new_n709), .A3(new_n882), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT124), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n931));
  INV_X1    g730(.A(new_n929), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n875), .A2(new_n905), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT123), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n926), .A2(new_n484), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n903), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n931), .B(new_n932), .C1(new_n937), .C2(new_n924), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n930), .A2(G148gat), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n922), .B1(new_n939), .B2(KEYINPUT59), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n899), .A2(new_n919), .A3(new_n783), .ZN(new_n941));
  OAI21_X1  g740(.A(KEYINPUT125), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  INV_X1    g742(.A(new_n941), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n925), .A2(new_n927), .ZN(new_n945));
  INV_X1    g744(.A(new_n924), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n929), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n374), .B1(new_n947), .B2(new_n931), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n920), .B1(new_n948), .B2(new_n930), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n943), .B(new_n944), .C1(new_n949), .C2(new_n922), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n942), .A2(new_n950), .ZN(G1345gat));
  INV_X1    g750(.A(new_n899), .ZN(new_n952));
  AOI21_X1  g751(.A(G155gat), .B1(new_n952), .B2(new_n733), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n733), .A2(G155gat), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(KEYINPUT126), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n953), .B1(new_n914), .B2(new_n955), .ZN(G1346gat));
  OAI21_X1  g755(.A(G162gat), .B1(new_n915), .B2(new_n731), .ZN(new_n957));
  OR3_X1    g756(.A1(new_n899), .A2(G162gat), .A3(new_n731), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1347gat));
  NAND3_X1  g758(.A1(new_n875), .A2(new_n712), .A3(new_n355), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n960), .A2(new_n877), .ZN(new_n961));
  AOI21_X1  g760(.A(G169gat), .B1(new_n961), .B2(new_n879), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n768), .A2(new_n356), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n881), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n687), .A2(new_n239), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1348gat));
  NAND3_X1  g765(.A1(new_n961), .A2(new_n240), .A3(new_n709), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n964), .A2(new_n709), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(new_n240), .ZN(G1349gat));
  NAND4_X1  g768(.A1(new_n961), .A2(new_n218), .A3(new_n222), .A4(new_n733), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n964), .A2(new_n733), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n971), .B2(new_n216), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g772(.A(new_n229), .B1(new_n964), .B2(new_n738), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT61), .Z(new_n975));
  NAND3_X1  g774(.A1(new_n961), .A2(new_n229), .A3(new_n738), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(G1351gat));
  NOR3_X1   g776(.A1(new_n960), .A2(new_n418), .A3(new_n753), .ZN(new_n978));
  AOI21_X1  g777(.A(G197gat), .B1(new_n978), .B2(new_n879), .ZN(new_n979));
  INV_X1    g778(.A(new_n963), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n928), .A2(new_n753), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n879), .A2(G197gat), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(G1352gat));
  INV_X1    g782(.A(G204gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n978), .A2(new_n984), .A3(new_n709), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT62), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n984), .B1(new_n981), .B2(new_n709), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n986), .A2(new_n987), .ZN(G1353gat));
  NAND3_X1  g787(.A1(new_n978), .A2(new_n319), .A3(new_n733), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n981), .A2(new_n733), .ZN(new_n991));
  AND4_X1   g790(.A1(new_n990), .A2(new_n991), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT63), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n319), .B1(KEYINPUT127), .B2(new_n993), .ZN(new_n994));
  AOI22_X1  g793(.A1(new_n991), .A2(new_n994), .B1(new_n990), .B2(KEYINPUT63), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n989), .B1(new_n992), .B2(new_n995), .ZN(G1354gat));
  AOI21_X1  g795(.A(G218gat), .B1(new_n978), .B2(new_n738), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n731), .A2(new_n318), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n997), .B1(new_n981), .B2(new_n998), .ZN(G1355gat));
endmodule


