//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G140), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(KEYINPUT78), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT78), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(new_n187), .A3(G125), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(KEYINPUT16), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT16), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n188), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT24), .B(G110), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G119), .ZN(new_n201));
  INV_X1    g015(.A(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G128), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT76), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n201), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(new_n201), .B2(new_n203), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n199), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT23), .B1(new_n200), .B2(G119), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n200), .A2(G119), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G110), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n200), .B(G119), .C1(KEYINPUT77), .C2(KEYINPUT23), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT65), .A2(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT65), .A2(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G125), .B(G140), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT80), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AND3_X1   g034(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT80), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n198), .B(new_n215), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n205), .A2(new_n206), .A3(new_n199), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n212), .B1(new_n211), .B2(new_n213), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT79), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n194), .A2(new_n227), .A3(new_n196), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n227), .B1(new_n194), .B2(new_n196), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n225), .B(new_n226), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n194), .A2(new_n227), .A3(new_n196), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n198), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n226), .B1(new_n233), .B2(new_n225), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n222), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(KEYINPUT81), .ZN(new_n236));
  AND2_X1   g050(.A1(KEYINPUT69), .A2(G953), .ZN(new_n237));
  NOR2_X1   g051(.A1(KEYINPUT69), .A2(G953), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n239), .A2(G221), .A3(G234), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G137), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n240), .B(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT81), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n244), .B(new_n222), .C1(new_n231), .C2(new_n234), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n236), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G902), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n242), .B(new_n222), .C1(new_n231), .C2(new_n234), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT82), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n233), .A2(new_n225), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(KEYINPUT79), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n230), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT82), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n252), .A2(new_n253), .A3(new_n242), .A4(new_n222), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n246), .A2(new_n247), .A3(new_n249), .A4(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n249), .A2(new_n254), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n258), .A2(KEYINPUT25), .A3(new_n247), .A4(new_n246), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G234), .ZN(new_n261));
  OAI21_X1  g075(.A(G217), .B1(new_n261), .B2(G902), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n262), .B(KEYINPUT75), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT83), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n260), .A2(KEYINPUT83), .A3(new_n263), .ZN(new_n267));
  INV_X1    g081(.A(new_n263), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n258), .A2(new_n247), .A3(new_n268), .A4(new_n246), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(KEYINPUT84), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n266), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT85), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT73), .ZN(new_n273));
  OR2_X1    g087(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n274));
  INV_X1    g088(.A(G137), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G134), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(KEYINPUT67), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G137), .ZN(new_n281));
  AND2_X1   g095(.A1(KEYINPUT11), .A2(G134), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n275), .A2(G134), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n278), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G131), .ZN(new_n287));
  INV_X1    g101(.A(G131), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n278), .A2(new_n283), .A3(new_n288), .A4(new_n285), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n227), .A2(G143), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n218), .B2(G143), .ZN(new_n292));
  AND2_X1   g106(.A1(KEYINPUT0), .A2(G128), .ZN(new_n293));
  NOR2_X1   g107(.A1(KEYINPUT0), .A2(G128), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n227), .A2(G143), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n296), .B1(new_n218), .B2(G143), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n292), .A2(new_n295), .B1(new_n297), .B2(new_n293), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  OR2_X1    g113(.A1(KEYINPUT65), .A2(G146), .ZN(new_n300));
  NAND2_X1  g114(.A1(KEYINPUT65), .A2(G146), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(G143), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n296), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n200), .B1(new_n302), .B2(KEYINPUT1), .ZN(new_n306));
  INV_X1    g120(.A(new_n291), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n300), .A2(new_n301), .ZN(new_n308));
  INV_X1    g122(.A(G143), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n305), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(G134), .B1(new_n279), .B2(new_n281), .ZN(new_n312));
  INV_X1    g126(.A(new_n276), .ZN(new_n313));
  OAI21_X1  g127(.A(G131), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n289), .A3(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(G116), .B(G119), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT2), .B(G113), .ZN(new_n317));
  XOR2_X1   g131(.A(new_n316), .B(new_n317), .Z(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n299), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n216), .A2(new_n217), .A3(new_n309), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n323));
  OAI21_X1  g137(.A(G128), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n324), .A2(new_n292), .B1(new_n297), .B2(new_n304), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n314), .A2(new_n289), .ZN(new_n326));
  OAI21_X1  g140(.A(KEYINPUT68), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n314), .A2(new_n289), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(new_n311), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n299), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n290), .A2(new_n298), .B1(new_n328), .B2(new_n311), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n331), .A2(new_n332), .B1(KEYINPUT30), .B2(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n321), .B1(new_n334), .B2(new_n318), .ZN(new_n335));
  XOR2_X1   g149(.A(KEYINPUT26), .B(G101), .Z(new_n336));
  OR2_X1    g150(.A1(KEYINPUT69), .A2(G953), .ZN(new_n337));
  INV_X1    g151(.A(G237), .ZN(new_n338));
  NAND2_X1  g152(.A1(KEYINPUT69), .A2(G953), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n337), .A2(G210), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT27), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n239), .A2(new_n342), .A3(G210), .A4(new_n338), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT70), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n344), .B1(new_n341), .B2(new_n343), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n336), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n343), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT70), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n350));
  INV_X1    g164(.A(new_n336), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n273), .B1(new_n335), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n353), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n331), .A2(new_n332), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n333), .A2(KEYINPUT30), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n356), .A2(new_n318), .A3(new_n357), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n355), .B(KEYINPUT73), .C1(new_n358), .C2(new_n321), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n315), .A2(KEYINPUT68), .B1(new_n290), .B2(new_n298), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n319), .B1(new_n361), .B2(new_n330), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT28), .B1(new_n362), .B2(new_n321), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT72), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n299), .A2(new_n315), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n299), .B2(new_n315), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n319), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT28), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n363), .A2(new_n369), .A3(new_n353), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n354), .A2(new_n359), .A3(new_n360), .A4(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n333), .A2(new_n319), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT28), .B1(new_n372), .B2(new_n321), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n355), .A2(new_n360), .ZN(new_n376));
  AOI21_X1  g190(.A(G902), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n371), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G472), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT32), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT31), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n353), .A2(new_n320), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT71), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n353), .A2(new_n320), .A3(KEYINPUT71), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n381), .B1(new_n358), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n334), .A2(new_n318), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n388), .A2(KEYINPUT31), .A3(new_n384), .A4(new_n385), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n353), .B1(new_n363), .B2(new_n369), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(G902), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G472), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n380), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(new_n387), .B2(new_n389), .ZN(new_n396));
  NOR4_X1   g210(.A1(new_n396), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n379), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT74), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT74), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n400), .B(new_n379), .C1(new_n395), .C2(new_n397), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT85), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n266), .A2(new_n402), .A3(new_n267), .A4(new_n270), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n272), .A2(new_n399), .A3(new_n401), .A4(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G478), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(KEYINPUT15), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n200), .A2(G143), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n309), .A2(G128), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(G134), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT101), .ZN(new_n412));
  INV_X1    g226(.A(G116), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n413), .A2(G122), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(G122), .ZN(new_n415));
  INV_X1    g229(.A(G107), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(KEYINPUT102), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n415), .A2(KEYINPUT14), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n419), .B1(new_n421), .B2(new_n415), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n412), .B(new_n418), .C1(new_n416), .C2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G134), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n410), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n414), .A2(new_n415), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(G107), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n417), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT13), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n409), .A2(new_n429), .ZN(new_n430));
  MUX2_X1   g244(.A(new_n430), .B(new_n429), .S(new_n408), .Z(new_n431));
  OAI211_X1 g245(.A(new_n425), .B(new_n428), .C1(new_n431), .C2(new_n424), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n423), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT9), .B(G234), .ZN(new_n434));
  INV_X1    g248(.A(G217), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n434), .A2(new_n435), .A3(G953), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n423), .A2(new_n432), .A3(new_n436), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n407), .B1(new_n440), .B2(new_n247), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n247), .A3(new_n407), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(G952), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(G953), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n261), .B2(new_n338), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(G898), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT103), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI211_X1 g265(.A(new_n247), .B(new_n239), .C1(G234), .C2(G237), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n444), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n337), .A2(G214), .A3(new_n338), .A4(new_n339), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n309), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n239), .A2(G143), .A3(G214), .A4(new_n338), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(KEYINPUT96), .A2(KEYINPUT18), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(G131), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n191), .A2(new_n193), .ZN(new_n462));
  OAI22_X1  g276(.A1(new_n221), .A2(new_n220), .B1(new_n462), .B2(new_n227), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n456), .B(new_n457), .C1(new_n288), .C2(new_n459), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n466));
  AOI211_X1 g280(.A(new_n466), .B(new_n288), .C1(new_n456), .C2(new_n457), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n456), .A2(new_n457), .A3(new_n288), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n288), .B1(new_n456), .B2(new_n457), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n467), .B1(new_n470), .B2(new_n466), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT99), .B1(new_n228), .B2(new_n229), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT99), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n198), .A2(new_n473), .A3(new_n232), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n465), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G113), .B(G122), .ZN(new_n477));
  XNOR2_X1  g291(.A(KEYINPUT98), .B(G104), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  AOI211_X1 g295(.A(new_n479), .B(new_n465), .C1(new_n471), .C2(new_n475), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n247), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G475), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT20), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT19), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n219), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n218), .B(new_n487), .C1(new_n462), .C2(new_n486), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n198), .B(new_n488), .C1(new_n468), .C2(new_n469), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT97), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT97), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n489), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n479), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n471), .A2(new_n475), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n480), .A3(new_n490), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(G475), .A2(G902), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n485), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n499), .ZN(new_n501));
  AOI211_X1 g315(.A(KEYINPUT20), .B(new_n501), .C1(new_n495), .C2(new_n497), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n484), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT100), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT100), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n484), .B(new_n505), .C1(new_n500), .C2(new_n502), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n454), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(G214), .B1(G237), .B2(G902), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n509), .B(KEYINPUT91), .Z(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n298), .A2(G125), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n311), .A2(new_n189), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G224), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(G953), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(KEYINPUT7), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT87), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT3), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n416), .A4(G104), .ZN(new_n521));
  INV_X1    g335(.A(G104), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n522), .A2(KEYINPUT87), .A3(G107), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT3), .B1(new_n522), .B2(G107), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G101), .ZN(new_n526));
  INV_X1    g340(.A(G101), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(new_n521), .C1(new_n523), .C2(new_n524), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(KEYINPUT4), .A3(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n529), .B(new_n318), .C1(KEYINPUT4), .C2(new_n526), .ZN(new_n530));
  INV_X1    g344(.A(new_n316), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n317), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT5), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n533), .A2(new_n202), .A3(KEYINPUT92), .A4(G116), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G113), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n533), .A2(new_n202), .A3(G116), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n316), .A2(KEYINPUT5), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT88), .B1(new_n416), .B2(G104), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT88), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n522), .A3(G107), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n541), .B(new_n543), .C1(new_n522), .C2(G107), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G101), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n528), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G110), .B(G122), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n530), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n517), .A2(KEYINPUT7), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n512), .A2(new_n513), .A3(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n518), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT93), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n539), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n316), .A2(KEYINPUT93), .A3(KEYINPUT5), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n532), .B1(new_n557), .B2(new_n538), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT94), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n547), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI211_X1 g374(.A(KEYINPUT94), .B(new_n532), .C1(new_n557), .C2(new_n538), .ZN(new_n561));
  OAI22_X1  g375(.A1(new_n560), .A2(new_n561), .B1(new_n547), .B2(new_n540), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n549), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(G902), .B1(new_n553), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G210), .B1(G237), .B2(G902), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n530), .A2(new_n548), .ZN(new_n567));
  INV_X1    g381(.A(new_n549), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(KEYINPUT6), .A3(new_n550), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n514), .B(new_n517), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT6), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n567), .A2(new_n572), .A3(new_n568), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n565), .A2(new_n566), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n566), .B1(new_n565), .B2(new_n574), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n511), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT95), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n553), .A2(new_n564), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n580), .A2(new_n574), .A3(new_n247), .ZN(new_n581));
  INV_X1    g395(.A(new_n566), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n510), .B1(new_n583), .B2(new_n575), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT95), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G469), .ZN(new_n588));
  OAI21_X1  g402(.A(G128), .B1(new_n307), .B2(new_n323), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n322), .B2(new_n296), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n305), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n547), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT10), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n546), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n592), .A2(new_n593), .B1(new_n594), .B2(new_n311), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n290), .B(KEYINPUT89), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n298), .B(new_n529), .C1(KEYINPUT4), .C2(new_n526), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(G110), .B(G140), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT86), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n239), .A2(G227), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n547), .A2(new_n311), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n546), .B1(new_n305), .B2(new_n590), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n290), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT12), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n592), .B1(new_n311), .B2(new_n547), .ZN(new_n608));
  AOI21_X1  g422(.A(KEYINPUT12), .B1(new_n608), .B2(new_n290), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n598), .B(new_n602), .C1(new_n607), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n594), .A2(new_n311), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n611), .B(new_n597), .C1(KEYINPUT10), .C2(new_n604), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n290), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n602), .B1(new_n613), .B2(new_n598), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT90), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n610), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI211_X1 g430(.A(KEYINPUT90), .B(new_n602), .C1(new_n613), .C2(new_n598), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n588), .B(new_n247), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n619));
  INV_X1    g433(.A(new_n602), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n598), .B1(new_n607), .B2(new_n609), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n621), .A2(new_n613), .B1(new_n622), .B2(new_n620), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(G469), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n588), .A2(new_n247), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n618), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(G221), .B1(new_n434), .B2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n508), .A2(new_n587), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n404), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n527), .ZN(G3));
  NAND2_X1  g447(.A1(new_n272), .A2(new_n403), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n390), .A2(new_n392), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n247), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(G472), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n393), .A2(new_n394), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n634), .A2(new_n629), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n440), .A2(new_n405), .A3(new_n247), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n440), .A2(KEYINPUT33), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT33), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n438), .B2(new_n439), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n247), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n643), .B1(new_n647), .B2(G478), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n648), .A2(new_n504), .A3(new_n506), .ZN(new_n649));
  INV_X1    g463(.A(new_n453), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n584), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n641), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  INV_X1    g469(.A(new_n503), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n444), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n658));
  OR3_X1    g472(.A1(new_n657), .A2(new_n651), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n658), .B1(new_n657), .B2(new_n651), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n641), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT35), .B(G107), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  AOI21_X1  g479(.A(KEYINPUT83), .B1(new_n260), .B2(new_n263), .ZN(new_n666));
  AOI211_X1 g480(.A(new_n265), .B(new_n268), .C1(new_n257), .C2(new_n259), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n236), .A2(new_n245), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n243), .A2(KEYINPUT36), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n669), .B(new_n670), .Z(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n247), .A3(new_n268), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n630), .A2(new_n639), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT105), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  INV_X1    g491(.A(new_n629), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n399), .A2(new_n401), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(G900), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n448), .B1(new_n452), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n657), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n673), .A2(new_n584), .A3(new_n682), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XNOR2_X1  g499(.A(KEYINPUT107), .B(KEYINPUT39), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n681), .B(new_n686), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n678), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT40), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n388), .A2(new_n384), .A3(new_n385), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n355), .B1(new_n372), .B2(new_n321), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(G472), .B1(new_n692), .B2(G902), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n395), .B2(new_n397), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n583), .A2(new_n575), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n696), .B(KEYINPUT38), .Z(new_n697));
  NOR3_X1   g511(.A1(new_n689), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n266), .A2(new_n267), .A3(new_n672), .ZN(new_n699));
  INV_X1    g513(.A(new_n506), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n494), .A2(new_n479), .ZN(new_n701));
  AOI22_X1  g515(.A1(new_n701), .A2(new_n492), .B1(new_n476), .B2(new_n480), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT20), .B1(new_n702), .B2(new_n501), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n498), .A2(new_n485), .A3(new_n499), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n505), .B1(new_n705), .B2(new_n484), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n699), .A2(new_n511), .A3(new_n707), .A4(new_n444), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  OR2_X1    g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n698), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G143), .ZN(G45));
  NOR2_X1   g527(.A1(new_n649), .A2(new_n681), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n673), .A2(new_n584), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n679), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n227), .ZN(G48));
  NAND2_X1  g531(.A1(new_n613), .A2(new_n598), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n620), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT90), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n614), .A2(new_n615), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n721), .A3(new_n610), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n588), .B1(new_n722), .B2(new_n247), .ZN(new_n723));
  INV_X1    g537(.A(new_n618), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n628), .ZN(new_n726));
  NOR4_X1   g540(.A1(new_n404), .A2(new_n649), .A3(new_n651), .A4(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT41), .B(G113), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n399), .A2(new_n401), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n726), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n272), .A3(new_n403), .A4(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n730), .B1(new_n734), .B2(new_n661), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n634), .A2(new_n731), .A3(new_n726), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n736), .A2(KEYINPUT108), .A3(new_n662), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G116), .ZN(G18));
  AOI21_X1  g553(.A(new_n508), .B1(new_n668), .B2(new_n672), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT109), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n725), .A2(new_n741), .A3(new_n584), .A4(new_n628), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n247), .B1(new_n616), .B2(new_n617), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(G469), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n744), .A2(new_n584), .A3(new_n628), .A4(new_n618), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT109), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n740), .A2(new_n399), .A3(new_n401), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G119), .ZN(G21));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n707), .A2(new_n750), .A3(new_n584), .A4(new_n444), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n504), .A2(new_n444), .A3(new_n584), .A4(new_n506), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT112), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n266), .A2(new_n267), .A3(new_n270), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n636), .A2(KEYINPUT111), .A3(G472), .ZN(new_n756));
  INV_X1    g570(.A(new_n390), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n374), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n369), .A2(KEYINPUT110), .A3(new_n373), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n353), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n394), .B(new_n247), .C1(new_n757), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n756), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n638), .A2(KEYINPUT111), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n726), .A2(new_n453), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n754), .A2(new_n755), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G122), .ZN(G24));
  NAND4_X1  g582(.A1(new_n747), .A2(new_n765), .A3(new_n673), .A4(new_n714), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G125), .ZN(G27));
  AND2_X1   g584(.A1(new_n755), .A2(new_n398), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n624), .B(KEYINPUT113), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n618), .A2(new_n626), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n696), .A2(new_n510), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n628), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n771), .A2(KEYINPUT42), .A3(new_n714), .A4(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n714), .ZN(new_n779));
  INV_X1    g593(.A(new_n777), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n404), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n778), .B1(new_n781), .B2(KEYINPUT42), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G131), .ZN(G33));
  NOR2_X1   g597(.A1(new_n404), .A2(new_n780), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n682), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  OAI21_X1  g600(.A(G469), .B1(new_n623), .B2(KEYINPUT45), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n621), .A2(new_n613), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n622), .A2(new_n620), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n788), .A2(KEYINPUT45), .A3(new_n789), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT114), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(KEYINPUT114), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n625), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n724), .B1(new_n794), .B2(KEYINPUT46), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n794), .A2(KEYINPUT46), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n628), .B(new_n687), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n775), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n507), .A2(new_n648), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT43), .Z(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n640), .A3(new_n673), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n800), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G137), .ZN(G39));
  OAI21_X1  g622(.A(new_n628), .B1(new_n796), .B2(new_n797), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g625(.A(KEYINPUT47), .B(new_n628), .C1(new_n796), .C2(new_n797), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n731), .A2(new_n714), .A3(new_n775), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n272), .B2(new_n403), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  NAND3_X1  g631(.A1(new_n748), .A2(new_n767), .A3(new_n674), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n579), .A2(new_n586), .A3(new_n650), .ZN(new_n819));
  INV_X1    g633(.A(new_n443), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT115), .B1(new_n820), .B2(new_n441), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n442), .A2(new_n822), .A3(new_n443), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n507), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n819), .B1(new_n825), .B2(new_n649), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n637), .A2(new_n629), .A3(new_n638), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n272), .A2(new_n826), .A3(new_n403), .A4(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n828), .B1(new_n404), .B2(new_n631), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n727), .A2(new_n818), .A3(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n824), .A2(new_n503), .A3(new_n681), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n673), .A2(new_n775), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n777), .A2(new_n714), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n765), .A2(new_n673), .ZN(new_n834));
  OAI22_X1  g648(.A1(new_n679), .A2(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n682), .B2(new_n784), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n830), .A2(new_n738), .A3(new_n782), .A4(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n769), .B1(new_n679), .B2(new_n683), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n716), .ZN(new_n839));
  INV_X1    g653(.A(new_n628), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n681), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n772), .ZN(new_n842));
  INV_X1    g656(.A(new_n773), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n699), .A2(new_n844), .A3(new_n694), .ZN(new_n845));
  INV_X1    g659(.A(new_n754), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT52), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n838), .A2(new_n716), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(KEYINPUT53), .B1(new_n837), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n736), .A2(new_n652), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n829), .A2(new_n818), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT108), .B1(new_n736), .B2(new_n662), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n404), .A2(new_n661), .A3(new_n730), .A4(new_n726), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n782), .A2(new_n836), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n838), .A2(new_n716), .A3(new_n849), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n679), .A2(new_n715), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n684), .A2(new_n863), .A3(new_n847), .A4(new_n769), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(new_n850), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n861), .A2(KEYINPUT52), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n860), .A2(new_n862), .A3(new_n868), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n853), .B(KEYINPUT54), .C1(new_n869), .C2(KEYINPUT53), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n860), .A2(KEYINPUT53), .A3(new_n862), .A4(new_n868), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n837), .B2(new_n852), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n725), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n776), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n695), .A2(new_n878), .A3(new_n448), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n634), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n707), .A3(new_n648), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n802), .A2(new_n448), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n755), .A2(new_n765), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n747), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n446), .B(new_n881), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n882), .A2(new_n878), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n771), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n889), .A2(KEYINPUT48), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(KEYINPUT48), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n885), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n877), .A2(new_n628), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n893), .B(new_n775), .C1(new_n813), .C2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n697), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n896), .A2(new_n511), .A3(new_n726), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT50), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  AND4_X1   g712(.A1(KEYINPUT50), .A2(new_n882), .A3(new_n884), .A4(new_n897), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n895), .B(KEYINPUT51), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n888), .A2(KEYINPUT118), .A3(new_n673), .A4(new_n765), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n882), .A2(new_n878), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n902), .B1(new_n903), .B2(new_n834), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n648), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n880), .A2(new_n507), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n892), .B1(new_n900), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n908), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT117), .B1(new_n898), .B2(new_n899), .ZN(new_n911));
  OR3_X1    g725(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT117), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n910), .A2(new_n895), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT51), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n909), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n876), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(G952), .B2(G953), .ZN(new_n917));
  NOR4_X1   g731(.A1(new_n896), .A2(new_n510), .A3(new_n840), .A4(new_n801), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n725), .B(KEYINPUT49), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n755), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n917), .B1(new_n694), .B2(new_n920), .ZN(G75));
  NOR2_X1   g735(.A1(new_n239), .A2(G952), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT119), .Z(new_n923));
  AOI21_X1  g737(.A(new_n247), .B1(new_n871), .B2(new_n873), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT56), .B1(new_n924), .B2(G210), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n570), .A2(new_n573), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(new_n571), .Z(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT55), .Z(new_n928));
  OAI21_X1  g742(.A(new_n923), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(G210), .ZN(new_n930));
  AOI211_X1 g744(.A(new_n930), .B(new_n247), .C1(new_n871), .C2(new_n873), .ZN(new_n931));
  INV_X1    g745(.A(new_n928), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n931), .A2(KEYINPUT56), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT120), .B1(new_n929), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n925), .A2(new_n928), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n932), .B1(new_n931), .B2(KEYINPUT56), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n935), .A2(new_n936), .A3(new_n937), .A4(new_n923), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n934), .A2(new_n938), .ZN(G51));
  NAND2_X1  g753(.A1(new_n871), .A2(new_n873), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT54), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n875), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n625), .B(KEYINPUT57), .Z(new_n944));
  OAI21_X1  g758(.A(new_n722), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n924), .A2(new_n793), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n922), .B1(new_n945), .B2(new_n946), .ZN(G54));
  NAND3_X1  g761(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n948), .A2(new_n702), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n702), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n922), .ZN(G60));
  NOR2_X1   g765(.A1(new_n644), .A2(new_n646), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT121), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(G478), .A2(G902), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT59), .Z(new_n956));
  OAI211_X1 g770(.A(KEYINPUT122), .B(new_n954), .C1(new_n876), .C2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT122), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n870), .B2(new_n875), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n953), .ZN(new_n960));
  INV_X1    g774(.A(new_n923), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n954), .A2(new_n956), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n961), .B1(new_n942), .B2(new_n962), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n957), .A2(new_n960), .A3(new_n963), .ZN(G63));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT60), .Z(new_n966));
  NAND3_X1  g780(.A1(new_n940), .A2(new_n671), .A3(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n940), .A2(new_n966), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n258), .A2(new_n246), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n923), .B(new_n967), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G66));
  OAI21_X1  g786(.A(G953), .B1(new_n451), .B2(new_n515), .ZN(new_n973));
  INV_X1    g787(.A(new_n858), .ZN(new_n974));
  INV_X1    g788(.A(new_n239), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n926), .B1(G898), .B2(new_n239), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G69));
  AND2_X1   g792(.A1(new_n807), .A2(new_n785), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n771), .A2(new_n754), .ZN(new_n980));
  OR3_X1    g794(.A1(new_n798), .A2(KEYINPUT124), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT124), .B1(new_n798), .B2(new_n980), .ZN(new_n982));
  AOI22_X1  g796(.A1(new_n981), .A2(new_n982), .B1(new_n813), .B2(new_n815), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n984), .A2(KEYINPUT125), .A3(new_n782), .A4(new_n839), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n979), .A2(new_n983), .A3(new_n782), .A4(new_n839), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n985), .A2(new_n988), .A3(new_n239), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n334), .B(KEYINPUT123), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n487), .B1(new_n462), .B2(new_n486), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n990), .B(new_n991), .Z(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(G900), .B2(new_n975), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n989), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n712), .A2(new_n839), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT62), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n799), .B(new_n688), .C1(new_n649), .C2(new_n825), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n997), .A2(new_n732), .A3(new_n272), .A4(new_n403), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n816), .A2(new_n807), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n239), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n239), .B1(G227), .B2(G900), .ZN(new_n1001));
  AOI22_X1  g815(.A1(new_n1000), .A2(new_n992), .B1(KEYINPUT126), .B2(new_n1001), .ZN(new_n1002));
  OR2_X1    g816(.A1(new_n1001), .A2(KEYINPUT126), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n994), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n994), .B2(new_n1002), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1004), .A2(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(new_n335), .A2(new_n355), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n985), .A2(new_n988), .A3(new_n974), .ZN(new_n1008));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT63), .Z(new_n1010));
  AOI21_X1  g824(.A(new_n1007), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1010), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n996), .A2(new_n999), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n1013), .B2(new_n974), .ZN(new_n1014));
  NOR3_X1   g828(.A1(new_n1014), .A2(new_n355), .A3(new_n335), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n853), .B1(new_n869), .B2(KEYINPUT53), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n354), .A2(new_n359), .A3(new_n690), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n1010), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT127), .Z(new_n1019));
  NOR2_X1   g833(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  NOR4_X1   g834(.A1(new_n1011), .A2(new_n1015), .A3(new_n922), .A4(new_n1020), .ZN(G57));
endmodule


