

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768;

  AND2_X1 U375 ( .A1(n371), .A2(n368), .ZN(n444) );
  OR2_X1 U376 ( .A1(n536), .A2(n374), .ZN(n370) );
  XNOR2_X1 U377 ( .A(n444), .B(n443), .ZN(n516) );
  XNOR2_X2 U378 ( .A(n482), .B(G134), .ZN(n468) );
  NOR2_X2 U379 ( .A1(n679), .A2(KEYINPUT44), .ZN(n605) );
  XNOR2_X2 U380 ( .A(n595), .B(KEYINPUT35), .ZN(n679) );
  INV_X1 U381 ( .A(n649), .ZN(n354) );
  AND2_X1 U382 ( .A1(n623), .A2(n622), .ZN(n629) );
  XNOR2_X1 U383 ( .A(n602), .B(KEYINPUT107), .ZN(n678) );
  AND2_X1 U384 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U385 ( .A1(n356), .A2(n376), .ZN(n601) );
  XNOR2_X1 U386 ( .A(n497), .B(n360), .ZN(n554) );
  OR2_X1 U387 ( .A1(n661), .A2(n646), .ZN(n493) );
  XNOR2_X1 U388 ( .A(G101), .B(KEYINPUT71), .ZN(n391) );
  XNOR2_X1 U389 ( .A(n651), .B(KEYINPUT85), .ZN(n641) );
  NOR2_X2 U390 ( .A1(n572), .A2(n571), .ZN(n573) );
  INV_X1 U391 ( .A(n379), .ZN(n355) );
  XNOR2_X1 U392 ( .A(n505), .B(KEYINPUT0), .ZN(n589) );
  BUF_X2 U393 ( .A(n508), .Z(n710) );
  XNOR2_X2 U394 ( .A(n433), .B(n432), .ZN(n532) );
  XNOR2_X2 U395 ( .A(n468), .B(n396), .ZN(n433) );
  XNOR2_X1 U396 ( .A(n479), .B(n424), .ZN(n531) );
  XNOR2_X1 U397 ( .A(G113), .B(G143), .ZN(n447) );
  AND2_X1 U398 ( .A1(n718), .A2(n374), .ZN(n373) );
  AND2_X1 U399 ( .A1(n370), .A2(n369), .ZN(n368) );
  NAND2_X1 U400 ( .A1(n523), .A2(KEYINPUT30), .ZN(n369) );
  XNOR2_X1 U401 ( .A(G119), .B(G128), .ZN(n414) );
  XNOR2_X1 U402 ( .A(n423), .B(G125), .ZN(n479) );
  INV_X1 U403 ( .A(KEYINPUT39), .ZN(n517) );
  NAND2_X1 U404 ( .A1(n359), .A2(n363), .ZN(n362) );
  INV_X1 U405 ( .A(G237), .ZN(n399) );
  XNOR2_X1 U406 ( .A(G116), .B(G113), .ZN(n392) );
  NOR2_X2 U407 ( .A1(G953), .A2(G237), .ZN(n451) );
  NAND2_X1 U408 ( .A1(G234), .A2(G237), .ZN(n403) );
  OR2_X1 U409 ( .A1(n689), .A2(G902), .ZN(n440) );
  BUF_X1 U410 ( .A(n641), .Z(n647) );
  NAND2_X1 U411 ( .A1(n354), .A2(n646), .ZN(n363) );
  INV_X1 U412 ( .A(G140), .ZN(n446) );
  XNOR2_X1 U413 ( .A(G110), .B(G107), .ZN(n437) );
  XNOR2_X1 U414 ( .A(KEYINPUT18), .B(KEYINPUT89), .ZN(n481) );
  XNOR2_X1 U415 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n483) );
  NOR2_X1 U416 ( .A1(n442), .A2(n372), .ZN(n371) );
  BUF_X1 U417 ( .A(n507), .Z(n614) );
  NAND2_X1 U418 ( .A1(n379), .A2(n377), .ZN(n376) );
  AND2_X1 U419 ( .A1(n717), .A2(n378), .ZN(n377) );
  XNOR2_X1 U420 ( .A(n710), .B(KEYINPUT6), .ZN(n587) );
  AND2_X1 U421 ( .A1(n697), .A2(G472), .ZN(n383) );
  XNOR2_X1 U422 ( .A(n426), .B(n425), .ZN(n680) );
  XNOR2_X1 U423 ( .A(n422), .B(n421), .ZN(n426) );
  AND2_X1 U424 ( .A1(n697), .A2(G210), .ZN(n382) );
  XOR2_X1 U425 ( .A(KEYINPUT91), .B(n658), .Z(n692) );
  OR2_X1 U426 ( .A1(n592), .A2(n519), .ZN(n759) );
  AND2_X1 U427 ( .A1(n381), .A2(n380), .ZN(n356) );
  AND2_X1 U428 ( .A1(n697), .A2(G478), .ZN(n357) );
  OR2_X1 U429 ( .A1(n355), .A2(n584), .ZN(n358) );
  AND2_X1 U430 ( .A1(n647), .A2(KEYINPUT83), .ZN(n359) );
  XOR2_X1 U431 ( .A(KEYINPUT76), .B(KEYINPUT19), .Z(n360) );
  OR2_X1 U432 ( .A1(n646), .A2(n645), .ZN(n361) );
  NAND2_X2 U433 ( .A1(n364), .A2(n362), .ZN(n653) );
  NAND2_X1 U434 ( .A1(n365), .A2(n361), .ZN(n364) );
  NAND2_X1 U435 ( .A1(n366), .A2(n385), .ZN(n365) );
  NAND2_X1 U436 ( .A1(n643), .A2(n642), .ZN(n366) );
  NOR2_X1 U437 ( .A1(n367), .A2(n768), .ZN(n545) );
  XNOR2_X1 U438 ( .A(n367), .B(n676), .ZN(G33) );
  XNOR2_X1 U439 ( .A(n543), .B(KEYINPUT40), .ZN(n367) );
  AND2_X1 U440 ( .A1(n536), .A2(n373), .ZN(n372) );
  INV_X1 U441 ( .A(KEYINPUT30), .ZN(n374) );
  XNOR2_X1 U442 ( .A(n508), .B(KEYINPUT106), .ZN(n536) );
  NAND2_X1 U443 ( .A1(n375), .A2(n506), .ZN(n380) );
  NAND2_X1 U444 ( .A1(n717), .A2(n700), .ZN(n375) );
  NAND2_X1 U445 ( .A1(n589), .A2(n506), .ZN(n381) );
  NOR2_X1 U446 ( .A1(n584), .A2(n506), .ZN(n378) );
  INV_X1 U447 ( .A(n589), .ZN(n379) );
  NAND2_X1 U448 ( .A1(n653), .A2(n382), .ZN(n665) );
  AND2_X1 U449 ( .A1(n653), .A2(n697), .ZN(n687) );
  NAND2_X1 U450 ( .A1(n653), .A2(n357), .ZN(n684) );
  NAND2_X1 U451 ( .A1(n653), .A2(n383), .ZN(n672) );
  NAND2_X1 U452 ( .A1(n653), .A2(n384), .ZN(n656) );
  AND2_X1 U453 ( .A1(n697), .A2(G475), .ZN(n384) );
  AND2_X1 U454 ( .A1(n646), .A2(n644), .ZN(n385) );
  XOR2_X1 U455 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n386) );
  NOR2_X1 U456 ( .A1(n568), .A2(n567), .ZN(n569) );
  INV_X1 U457 ( .A(KEYINPUT83), .ZN(n642) );
  XNOR2_X1 U458 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U459 ( .A(n586), .B(KEYINPUT74), .ZN(n607) );
  BUF_X1 U460 ( .A(n607), .Z(n711) );
  INV_X1 U461 ( .A(KEYINPUT75), .ZN(n443) );
  NAND2_X1 U462 ( .A1(n451), .A2(G210), .ZN(n388) );
  INV_X1 U463 ( .A(G137), .ZN(n387) );
  XNOR2_X1 U464 ( .A(n388), .B(n387), .ZN(n390) );
  XNOR2_X1 U465 ( .A(G146), .B(KEYINPUT5), .ZN(n389) );
  XNOR2_X1 U466 ( .A(n390), .B(n389), .ZN(n395) );
  XNOR2_X1 U467 ( .A(n392), .B(n391), .ZN(n394) );
  XNOR2_X1 U468 ( .A(KEYINPUT3), .B(G119), .ZN(n393) );
  XNOR2_X1 U469 ( .A(n394), .B(n393), .ZN(n477) );
  XNOR2_X1 U470 ( .A(n395), .B(n477), .ZN(n397) );
  XNOR2_X2 U471 ( .A(G143), .B(G128), .ZN(n482) );
  XNOR2_X1 U472 ( .A(KEYINPUT4), .B(G131), .ZN(n396) );
  XNOR2_X1 U473 ( .A(n397), .B(n433), .ZN(n668) );
  OR2_X1 U474 ( .A1(n668), .A2(G902), .ZN(n398) );
  XNOR2_X1 U475 ( .A(n398), .B(G472), .ZN(n508) );
  INV_X1 U476 ( .A(G902), .ZN(n472) );
  NAND2_X1 U477 ( .A1(n472), .A2(n399), .ZN(n489) );
  AND2_X1 U478 ( .A1(n489), .A2(G214), .ZN(n523) );
  INV_X1 U479 ( .A(n523), .ZN(n718) );
  XNOR2_X1 U480 ( .A(G902), .B(KEYINPUT92), .ZN(n400) );
  XNOR2_X1 U481 ( .A(n400), .B(KEYINPUT15), .ZN(n648) );
  NAND2_X1 U482 ( .A1(n648), .A2(G234), .ZN(n401) );
  XNOR2_X1 U483 ( .A(KEYINPUT20), .B(n401), .ZN(n427) );
  AND2_X1 U484 ( .A1(n427), .A2(G221), .ZN(n402) );
  XNOR2_X1 U485 ( .A(n402), .B(KEYINPUT21), .ZN(n700) );
  XNOR2_X1 U486 ( .A(n403), .B(KEYINPUT14), .ZN(n411) );
  NAND2_X1 U487 ( .A1(n411), .A2(G902), .ZN(n404) );
  XOR2_X1 U488 ( .A(KEYINPUT94), .B(n404), .Z(n499) );
  INV_X1 U489 ( .A(KEYINPUT64), .ZN(n405) );
  XNOR2_X2 U490 ( .A(n405), .B(G953), .ZN(n657) );
  INV_X1 U491 ( .A(n657), .ZN(n406) );
  NAND2_X1 U492 ( .A1(n499), .A2(n406), .ZN(n408) );
  INV_X1 U493 ( .A(KEYINPUT108), .ZN(n407) );
  XNOR2_X1 U494 ( .A(n408), .B(n407), .ZN(n410) );
  INV_X1 U495 ( .A(G900), .ZN(n409) );
  NAND2_X1 U496 ( .A1(n410), .A2(n409), .ZN(n412) );
  NAND2_X1 U497 ( .A1(G952), .A2(n411), .ZN(n734) );
  OR2_X1 U498 ( .A1(G953), .A2(n734), .ZN(n500) );
  NAND2_X1 U499 ( .A1(n412), .A2(n500), .ZN(n413) );
  AND2_X1 U500 ( .A1(n700), .A2(n413), .ZN(n520) );
  INV_X1 U501 ( .A(n520), .ZN(n431) );
  XOR2_X1 U502 ( .A(KEYINPUT23), .B(G110), .Z(n415) );
  XNOR2_X1 U503 ( .A(n415), .B(n414), .ZN(n417) );
  XNOR2_X1 U504 ( .A(G137), .B(G140), .ZN(n432) );
  INV_X1 U505 ( .A(n432), .ZN(n416) );
  XOR2_X1 U506 ( .A(n417), .B(n416), .Z(n422) );
  XNOR2_X1 U507 ( .A(KEYINPUT8), .B(KEYINPUT68), .ZN(n418) );
  XNOR2_X1 U508 ( .A(n418), .B(KEYINPUT69), .ZN(n420) );
  NAND2_X1 U509 ( .A1(n657), .A2(G234), .ZN(n419) );
  XNOR2_X1 U510 ( .A(n420), .B(n419), .ZN(n469) );
  NAND2_X1 U511 ( .A1(n469), .A2(G221), .ZN(n421) );
  INV_X1 U512 ( .A(G146), .ZN(n423) );
  INV_X1 U513 ( .A(KEYINPUT10), .ZN(n424) );
  XNOR2_X1 U514 ( .A(n531), .B(KEYINPUT24), .ZN(n425) );
  NAND2_X1 U515 ( .A1(n680), .A2(n472), .ZN(n430) );
  NAND2_X1 U516 ( .A1(G217), .A2(n427), .ZN(n428) );
  XNOR2_X1 U517 ( .A(KEYINPUT25), .B(n428), .ZN(n429) );
  XNOR2_X2 U518 ( .A(n430), .B(n429), .ZN(n613) );
  NOR2_X1 U519 ( .A1(n431), .A2(n613), .ZN(n441) );
  NAND2_X1 U520 ( .A1(n657), .A2(G227), .ZN(n436) );
  XNOR2_X1 U521 ( .A(G101), .B(G146), .ZN(n434) );
  XNOR2_X1 U522 ( .A(KEYINPUT77), .B(n434), .ZN(n435) );
  XNOR2_X1 U523 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U524 ( .A(n437), .B(G104), .ZN(n476) );
  XNOR2_X1 U525 ( .A(n438), .B(n476), .ZN(n439) );
  XNOR2_X1 U526 ( .A(n532), .B(n439), .ZN(n689) );
  XNOR2_X2 U527 ( .A(n440), .B(G469), .ZN(n507) );
  NAND2_X1 U528 ( .A1(n441), .A2(n614), .ZN(n442) );
  XNOR2_X1 U529 ( .A(G131), .B(KEYINPUT99), .ZN(n445) );
  XNOR2_X1 U530 ( .A(n386), .B(n445), .ZN(n449) );
  XNOR2_X1 U531 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U532 ( .A(n531), .B(n450), .Z(n457) );
  NAND2_X1 U533 ( .A1(n451), .A2(G214), .ZN(n453) );
  XNOR2_X1 U534 ( .A(G122), .B(G104), .ZN(n452) );
  XNOR2_X1 U535 ( .A(n453), .B(n452), .ZN(n455) );
  XOR2_X1 U536 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n454) );
  XNOR2_X1 U537 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U538 ( .A(n457), .B(n456), .ZN(n654) );
  NOR2_X1 U539 ( .A1(n654), .A2(G902), .ZN(n459) );
  XNOR2_X1 U540 ( .A(KEYINPUT13), .B(KEYINPUT101), .ZN(n458) );
  XNOR2_X1 U541 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X2 U542 ( .A(n460), .B(G475), .ZN(n592) );
  XOR2_X1 U543 ( .A(KEYINPUT7), .B(G107), .Z(n462) );
  XNOR2_X1 U544 ( .A(G116), .B(G122), .ZN(n461) );
  XNOR2_X1 U545 ( .A(n462), .B(n461), .ZN(n466) );
  XOR2_X1 U546 ( .A(KEYINPUT102), .B(KEYINPUT9), .Z(n464) );
  XNOR2_X1 U547 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n463) );
  XNOR2_X1 U548 ( .A(n464), .B(n463), .ZN(n465) );
  XOR2_X1 U549 ( .A(n466), .B(n465), .Z(n467) );
  XNOR2_X1 U550 ( .A(n468), .B(n467), .ZN(n471) );
  AND2_X1 U551 ( .A1(n469), .A2(G217), .ZN(n470) );
  XNOR2_X1 U552 ( .A(n471), .B(n470), .ZN(n685) );
  NAND2_X1 U553 ( .A1(n685), .A2(n472), .ZN(n474) );
  INV_X1 U554 ( .A(G478), .ZN(n473) );
  XNOR2_X1 U555 ( .A(n474), .B(n473), .ZN(n591) );
  INV_X1 U556 ( .A(n591), .ZN(n519) );
  XNOR2_X1 U557 ( .A(KEYINPUT16), .B(G122), .ZN(n475) );
  XNOR2_X1 U558 ( .A(n476), .B(n475), .ZN(n478) );
  XNOR2_X1 U559 ( .A(n478), .B(n477), .ZN(n638) );
  NAND2_X1 U560 ( .A1(n657), .A2(G224), .ZN(n480) );
  XNOR2_X1 U561 ( .A(n480), .B(n479), .ZN(n487) );
  XNOR2_X1 U562 ( .A(n482), .B(n481), .ZN(n485) );
  XNOR2_X1 U563 ( .A(n483), .B(KEYINPUT93), .ZN(n484) );
  XNOR2_X1 U564 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U565 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U566 ( .A(n638), .B(n488), .ZN(n661) );
  INV_X1 U567 ( .A(n648), .ZN(n646) );
  NAND2_X1 U568 ( .A1(n489), .A2(G210), .ZN(n491) );
  INV_X1 U569 ( .A(KEYINPUT79), .ZN(n490) );
  XNOR2_X1 U570 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X2 U571 ( .A(n493), .B(n492), .ZN(n496) );
  INV_X1 U572 ( .A(n496), .ZN(n546) );
  NAND2_X1 U573 ( .A1(n519), .A2(n546), .ZN(n494) );
  NOR2_X1 U574 ( .A1(n592), .A2(n494), .ZN(n495) );
  AND2_X1 U575 ( .A1(n516), .A2(n495), .ZN(n567) );
  XOR2_X1 U576 ( .A(G143), .B(n567), .Z(G45) );
  NOR2_X2 U577 ( .A1(n496), .A2(n523), .ZN(n497) );
  INV_X1 U578 ( .A(G898), .ZN(n498) );
  AND2_X1 U579 ( .A1(n498), .A2(G953), .ZN(n636) );
  NAND2_X1 U580 ( .A1(n499), .A2(n636), .ZN(n501) );
  NAND2_X1 U581 ( .A1(n501), .A2(n500), .ZN(n503) );
  INV_X1 U582 ( .A(KEYINPUT95), .ZN(n502) );
  XNOR2_X1 U583 ( .A(n503), .B(n502), .ZN(n504) );
  NAND2_X1 U584 ( .A1(n554), .A2(n504), .ZN(n505) );
  INV_X1 U585 ( .A(n700), .ZN(n584) );
  AND2_X1 U586 ( .A1(n592), .A2(n591), .ZN(n717) );
  XNOR2_X1 U587 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n506) );
  XNOR2_X2 U588 ( .A(n507), .B(KEYINPUT1), .ZN(n585) );
  XNOR2_X1 U589 ( .A(n585), .B(KEYINPUT90), .ZN(n551) );
  INV_X1 U590 ( .A(n587), .ZN(n509) );
  INV_X1 U591 ( .A(n613), .ZN(n699) );
  NOR2_X1 U592 ( .A1(n509), .A2(n699), .ZN(n510) );
  NAND2_X1 U593 ( .A1(n551), .A2(n510), .ZN(n511) );
  XOR2_X1 U594 ( .A(KEYINPUT78), .B(n511), .Z(n512) );
  NAND2_X1 U595 ( .A1(n601), .A2(n512), .ZN(n514) );
  XNOR2_X1 U596 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n513) );
  XNOR2_X1 U597 ( .A(n514), .B(n513), .ZN(n603) );
  XNOR2_X1 U598 ( .A(G119), .B(KEYINPUT126), .ZN(n515) );
  XNOR2_X1 U599 ( .A(n603), .B(n515), .ZN(G21) );
  XNOR2_X1 U600 ( .A(n496), .B(KEYINPUT38), .ZN(n719) );
  NAND2_X1 U601 ( .A1(n516), .A2(n719), .ZN(n518) );
  XNOR2_X2 U602 ( .A(n518), .B(n517), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n592), .A2(n519), .ZN(n761) );
  NOR2_X1 U604 ( .A1(n542), .A2(n761), .ZN(n575) );
  XOR2_X1 U605 ( .A(G134), .B(n575), .Z(G36) );
  XNOR2_X1 U606 ( .A(n520), .B(KEYINPUT70), .ZN(n521) );
  AND2_X1 U607 ( .A1(n613), .A2(n521), .ZN(n537) );
  INV_X1 U608 ( .A(n537), .ZN(n522) );
  NOR2_X1 U609 ( .A1(n759), .A2(n522), .ZN(n547) );
  OR2_X1 U610 ( .A1(n587), .A2(n523), .ZN(n548) );
  INV_X1 U611 ( .A(n548), .ZN(n524) );
  NAND2_X1 U612 ( .A1(n547), .A2(n524), .ZN(n525) );
  INV_X1 U613 ( .A(n585), .ZN(n599) );
  INV_X1 U614 ( .A(n599), .ZN(n702) );
  NOR2_X1 U615 ( .A1(n525), .A2(n702), .ZN(n526) );
  XNOR2_X1 U616 ( .A(n526), .B(KEYINPUT43), .ZN(n527) );
  NOR2_X1 U617 ( .A1(n527), .A2(n546), .ZN(n574) );
  XOR2_X1 U618 ( .A(G140), .B(n574), .Z(G42) );
  NAND2_X1 U619 ( .A1(n601), .A2(n599), .ZN(n529) );
  NAND2_X1 U620 ( .A1(n699), .A2(n587), .ZN(n528) );
  NOR2_X1 U621 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U622 ( .A(KEYINPUT105), .B(n530), .Z(n620) );
  XOR2_X1 U623 ( .A(G101), .B(n620), .Z(G3) );
  XOR2_X1 U624 ( .A(n532), .B(n531), .Z(n579) );
  XOR2_X1 U625 ( .A(KEYINPUT110), .B(KEYINPUT41), .Z(n535) );
  NAND2_X1 U626 ( .A1(n719), .A2(n718), .ZN(n533) );
  XNOR2_X1 U627 ( .A(n533), .B(KEYINPUT109), .ZN(n723) );
  NAND2_X1 U628 ( .A1(n723), .A2(n717), .ZN(n534) );
  XNOR2_X1 U629 ( .A(n535), .B(n534), .ZN(n736) );
  BUF_X1 U630 ( .A(n536), .Z(n596) );
  NAND2_X1 U631 ( .A1(n537), .A2(n596), .ZN(n538) );
  XNOR2_X1 U632 ( .A(n538), .B(KEYINPUT28), .ZN(n540) );
  INV_X1 U633 ( .A(n614), .ZN(n539) );
  OR2_X1 U634 ( .A1(n540), .A2(n539), .ZN(n553) );
  NOR2_X1 U635 ( .A1(n736), .A2(n553), .ZN(n541) );
  XNOR2_X1 U636 ( .A(n541), .B(KEYINPUT42), .ZN(n768) );
  NOR2_X2 U637 ( .A1(n542), .A2(n759), .ZN(n543) );
  XOR2_X1 U638 ( .A(KEYINPUT86), .B(KEYINPUT46), .Z(n544) );
  XNOR2_X1 U639 ( .A(n545), .B(n544), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n547), .A2(n546), .ZN(n549) );
  NOR2_X1 U641 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U642 ( .A(n550), .B(KEYINPUT36), .ZN(n552) );
  NAND2_X1 U643 ( .A1(n552), .A2(n551), .ZN(n767) );
  INV_X1 U644 ( .A(n553), .ZN(n555) );
  NAND2_X1 U645 ( .A1(n555), .A2(n554), .ZN(n557) );
  NAND2_X1 U646 ( .A1(n557), .A2(KEYINPUT47), .ZN(n556) );
  NAND2_X1 U647 ( .A1(n767), .A2(n556), .ZN(n563) );
  INV_X1 U648 ( .A(n557), .ZN(n757) );
  NOR2_X1 U649 ( .A1(KEYINPUT47), .A2(KEYINPUT67), .ZN(n558) );
  NAND2_X1 U650 ( .A1(n757), .A2(n558), .ZN(n560) );
  NAND2_X1 U651 ( .A1(KEYINPUT67), .A2(KEYINPUT47), .ZN(n559) );
  NAND2_X1 U652 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U653 ( .A1(n759), .A2(n761), .ZN(n722) );
  AND2_X1 U654 ( .A1(n561), .A2(n722), .ZN(n562) );
  NOR2_X1 U655 ( .A1(n563), .A2(n562), .ZN(n564) );
  INV_X1 U656 ( .A(n722), .ZN(n565) );
  NAND2_X1 U657 ( .A1(KEYINPUT47), .A2(n565), .ZN(n566) );
  XOR2_X1 U658 ( .A(KEYINPUT82), .B(n566), .Z(n568) );
  XOR2_X1 U659 ( .A(KEYINPUT81), .B(n569), .Z(n570) );
  NAND2_X1 U660 ( .A1(n564), .A2(n570), .ZN(n571) );
  XNOR2_X1 U661 ( .A(n573), .B(KEYINPUT48), .ZN(n577) );
  NOR2_X1 U662 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U663 ( .A1(n577), .A2(n576), .ZN(n651) );
  XOR2_X1 U664 ( .A(n579), .B(n647), .Z(n578) );
  NAND2_X1 U665 ( .A1(n578), .A2(n657), .ZN(n583) );
  XNOR2_X1 U666 ( .A(G227), .B(n579), .ZN(n580) );
  NAND2_X1 U667 ( .A1(n580), .A2(G900), .ZN(n581) );
  NAND2_X1 U668 ( .A1(n581), .A2(G953), .ZN(n582) );
  NAND2_X1 U669 ( .A1(n583), .A2(n582), .ZN(G72) );
  NOR2_X1 U670 ( .A1(n584), .A2(n613), .ZN(n703) );
  NAND2_X1 U671 ( .A1(n703), .A2(n585), .ZN(n586) );
  NOR2_X1 U672 ( .A1(n607), .A2(n587), .ZN(n588) );
  XNOR2_X1 U673 ( .A(n588), .B(KEYINPUT33), .ZN(n727) );
  NOR2_X1 U674 ( .A1(n727), .A2(n355), .ZN(n590) );
  XNOR2_X1 U675 ( .A(n590), .B(KEYINPUT34), .ZN(n594) );
  NOR2_X1 U676 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U677 ( .A1(n594), .A2(n593), .ZN(n595) );
  INV_X1 U678 ( .A(n596), .ZN(n597) );
  AND2_X1 U679 ( .A1(n597), .A2(n613), .ZN(n598) );
  AND2_X1 U680 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U681 ( .A1(n678), .A2(n603), .ZN(n604) );
  XNOR2_X2 U682 ( .A(n604), .B(KEYINPUT87), .ZN(n624) );
  NAND2_X1 U683 ( .A1(n605), .A2(n624), .ZN(n606) );
  XNOR2_X1 U684 ( .A(n606), .B(KEYINPUT72), .ZN(n623) );
  NAND2_X1 U685 ( .A1(n679), .A2(KEYINPUT44), .ZN(n619) );
  INV_X1 U686 ( .A(n711), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n608), .A2(n710), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n609), .A2(n355), .ZN(n612) );
  XOR2_X1 U689 ( .A(KEYINPUT31), .B(KEYINPUT96), .Z(n610) );
  XNOR2_X1 U690 ( .A(n610), .B(KEYINPUT97), .ZN(n611) );
  XNOR2_X1 U691 ( .A(n612), .B(n611), .ZN(n762) );
  NOR2_X1 U692 ( .A1(n613), .A2(n710), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n616) );
  OR2_X1 U694 ( .A1(n358), .A2(n616), .ZN(n747) );
  NAND2_X1 U695 ( .A1(n762), .A2(n747), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n617), .A2(n722), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(n621) );
  NOR2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n622) );
  INV_X1 U699 ( .A(KEYINPUT65), .ZN(n627) );
  INV_X1 U700 ( .A(n624), .ZN(n625) );
  NAND2_X1 U701 ( .A1(n625), .A2(KEYINPUT44), .ZN(n626) );
  XNOR2_X1 U702 ( .A(n627), .B(n626), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X2 U704 ( .A(n630), .B(KEYINPUT45), .ZN(n650) );
  INV_X1 U705 ( .A(n650), .ZN(n649) );
  NOR2_X1 U706 ( .A1(n649), .A2(G953), .ZN(n635) );
  NAND2_X1 U707 ( .A1(G953), .A2(G224), .ZN(n631) );
  XNOR2_X1 U708 ( .A(KEYINPUT61), .B(n631), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n632), .A2(G898), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n633), .B(KEYINPUT125), .ZN(n634) );
  NOR2_X1 U711 ( .A1(n635), .A2(n634), .ZN(n640) );
  INV_X1 U712 ( .A(n636), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U714 ( .A(n640), .B(n639), .ZN(G69) );
  NAND2_X1 U715 ( .A1(n650), .A2(n641), .ZN(n694) );
  INV_X1 U716 ( .A(n694), .ZN(n643) );
  NAND2_X1 U717 ( .A1(KEYINPUT2), .A2(KEYINPUT84), .ZN(n644) );
  INV_X1 U718 ( .A(KEYINPUT2), .ZN(n695) );
  NOR2_X1 U719 ( .A1(n695), .A2(KEYINPUT84), .ZN(n645) );
  NOR2_X1 U720 ( .A1(n651), .A2(n695), .ZN(n652) );
  NAND2_X1 U721 ( .A1(n354), .A2(n652), .ZN(n697) );
  XOR2_X1 U722 ( .A(KEYINPUT59), .B(n654), .Z(n655) );
  XNOR2_X1 U723 ( .A(n656), .B(n655), .ZN(n659) );
  NOR2_X1 U724 ( .A1(n657), .A2(G952), .ZN(n658) );
  NOR2_X2 U725 ( .A1(n659), .A2(n692), .ZN(n660) );
  XNOR2_X1 U726 ( .A(n660), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U727 ( .A(KEYINPUT88), .B(KEYINPUT54), .ZN(n662) );
  XOR2_X1 U728 ( .A(n662), .B(KEYINPUT55), .Z(n663) );
  XNOR2_X1 U729 ( .A(n661), .B(n663), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n665), .B(n664), .ZN(n666) );
  NOR2_X2 U731 ( .A1(n666), .A2(n692), .ZN(n667) );
  XNOR2_X1 U732 ( .A(n667), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U733 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n669) );
  XNOR2_X1 U734 ( .A(n669), .B(KEYINPUT62), .ZN(n670) );
  XNOR2_X1 U735 ( .A(n668), .B(n670), .ZN(n671) );
  XNOR2_X1 U736 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X2 U737 ( .A1(n673), .A2(n692), .ZN(n675) );
  INV_X1 U738 ( .A(KEYINPUT63), .ZN(n674) );
  XNOR2_X1 U739 ( .A(n675), .B(n674), .ZN(G57) );
  XNOR2_X1 U740 ( .A(G131), .B(KEYINPUT127), .ZN(n676) );
  XNOR2_X1 U741 ( .A(G110), .B(KEYINPUT114), .ZN(n677) );
  XNOR2_X1 U742 ( .A(n678), .B(n677), .ZN(G12) );
  XOR2_X1 U743 ( .A(n679), .B(G122), .Z(G24) );
  NAND2_X1 U744 ( .A1(n687), .A2(G217), .ZN(n682) );
  XOR2_X1 U745 ( .A(KEYINPUT124), .B(n680), .Z(n681) );
  XNOR2_X1 U746 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U747 ( .A1(n683), .A2(n692), .ZN(G66) );
  XOR2_X1 U748 ( .A(n685), .B(n684), .Z(n686) );
  NOR2_X1 U749 ( .A1(n686), .A2(n692), .ZN(G63) );
  NAND2_X1 U750 ( .A1(n687), .A2(G469), .ZN(n691) );
  XOR2_X1 U751 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n688) );
  XNOR2_X1 U752 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U753 ( .A(n691), .B(n690), .ZN(n693) );
  NOR2_X1 U754 ( .A1(n693), .A2(n692), .ZN(G54) );
  NAND2_X1 U755 ( .A1(n694), .A2(n695), .ZN(n696) );
  XNOR2_X1 U756 ( .A(n696), .B(KEYINPUT80), .ZN(n698) );
  NAND2_X1 U757 ( .A1(n698), .A2(n697), .ZN(n743) );
  NOR2_X1 U758 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U759 ( .A(KEYINPUT49), .B(n701), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U761 ( .A(KEYINPUT50), .B(n704), .Z(n705) );
  XNOR2_X1 U762 ( .A(KEYINPUT118), .B(n705), .ZN(n706) );
  NAND2_X1 U763 ( .A1(n707), .A2(n706), .ZN(n709) );
  INV_X1 U764 ( .A(n710), .ZN(n708) );
  NAND2_X1 U765 ( .A1(n709), .A2(n708), .ZN(n713) );
  NAND2_X1 U766 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U767 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U768 ( .A(n714), .B(KEYINPUT51), .ZN(n715) );
  XNOR2_X1 U769 ( .A(KEYINPUT119), .B(n715), .ZN(n716) );
  NOR2_X1 U770 ( .A1(n736), .A2(n716), .ZN(n732) );
  INV_X1 U771 ( .A(n717), .ZN(n721) );
  NOR2_X1 U772 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U775 ( .A(KEYINPUT120), .B(n724), .Z(n725) );
  NOR2_X1 U776 ( .A1(n726), .A2(n725), .ZN(n729) );
  BUF_X1 U777 ( .A(n727), .Z(n728) );
  NOR2_X1 U778 ( .A1(n729), .A2(n728), .ZN(n730) );
  XOR2_X1 U779 ( .A(KEYINPUT121), .B(n730), .Z(n731) );
  NOR2_X1 U780 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U781 ( .A(n733), .B(KEYINPUT52), .ZN(n735) );
  NOR2_X1 U782 ( .A1(n735), .A2(n734), .ZN(n741) );
  NOR2_X1 U783 ( .A1(n736), .A2(n728), .ZN(n737) );
  XOR2_X1 U784 ( .A(KEYINPUT122), .B(n737), .Z(n739) );
  INV_X1 U785 ( .A(G953), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U787 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U788 ( .A1(n743), .A2(n742), .ZN(n745) );
  XNOR2_X1 U789 ( .A(KEYINPUT123), .B(KEYINPUT53), .ZN(n744) );
  XNOR2_X1 U790 ( .A(n745), .B(n744), .ZN(G75) );
  NOR2_X1 U791 ( .A1(n759), .A2(n747), .ZN(n746) );
  XOR2_X1 U792 ( .A(G104), .B(n746), .Z(G6) );
  NOR2_X1 U793 ( .A1(n747), .A2(n761), .ZN(n751) );
  XOR2_X1 U794 ( .A(KEYINPUT27), .B(KEYINPUT113), .Z(n749) );
  XNOR2_X1 U795 ( .A(G107), .B(KEYINPUT26), .ZN(n748) );
  XNOR2_X1 U796 ( .A(n749), .B(n748), .ZN(n750) );
  XNOR2_X1 U797 ( .A(n751), .B(n750), .ZN(G9) );
  XNOR2_X1 U798 ( .A(KEYINPUT115), .B(KEYINPUT29), .ZN(n754) );
  INV_X1 U799 ( .A(n761), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n757), .A2(n752), .ZN(n753) );
  XNOR2_X1 U801 ( .A(n754), .B(n753), .ZN(n755) );
  XNOR2_X1 U802 ( .A(G128), .B(n755), .ZN(G30) );
  INV_X1 U803 ( .A(n759), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U805 ( .A(G146), .B(n758), .ZN(G48) );
  NOR2_X1 U806 ( .A1(n762), .A2(n759), .ZN(n760) );
  XOR2_X1 U807 ( .A(G113), .B(n760), .Z(G15) );
  NOR2_X1 U808 ( .A1(n762), .A2(n761), .ZN(n764) );
  XNOR2_X1 U809 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n763) );
  XNOR2_X1 U810 ( .A(n764), .B(n763), .ZN(n765) );
  XNOR2_X1 U811 ( .A(G116), .B(n765), .ZN(G18) );
  XOR2_X1 U812 ( .A(G125), .B(KEYINPUT37), .Z(n766) );
  XNOR2_X1 U813 ( .A(n767), .B(n766), .ZN(G27) );
  XOR2_X1 U814 ( .A(G137), .B(n768), .Z(G39) );
endmodule

