//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  INV_X1    g000(.A(KEYINPUT96), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT74), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n192), .A2(G227), .ZN(new_n193));
  XOR2_X1   g007(.A(new_n191), .B(new_n193), .Z(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G146), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n198), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT68), .A3(new_n196), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n204), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n199), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  OAI21_X1  g023(.A(G128), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT79), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n195), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT79), .B1(new_n213), .B2(new_n204), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n206), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  AND2_X1   g030(.A1(KEYINPUT75), .A2(G107), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT75), .A2(G107), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT78), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n216), .B2(G107), .ZN(new_n221));
  INV_X1    g035(.A(G107), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT78), .A3(G104), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n219), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(G104), .B2(new_n222), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n217), .A2(new_n218), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n216), .A2(KEYINPUT3), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(G101), .B1(new_n216), .B2(G107), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n224), .A2(G101), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT10), .B1(new_n215), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G101), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n216), .A2(G107), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n233), .B1(new_n229), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT75), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n222), .ZN(new_n237));
  NAND2_X1  g051(.A1(KEYINPUT75), .A2(G107), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n228), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT3), .B1(new_n216), .B2(G107), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(new_n230), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT4), .ZN(new_n242));
  OAI21_X1  g056(.A(KEYINPUT76), .B1(new_n235), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n239), .A2(new_n240), .A3(new_n234), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G101), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT76), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n245), .A2(new_n246), .A3(KEYINPUT4), .A4(new_n241), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT64), .B1(new_n197), .B2(G143), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT64), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(new_n199), .A3(G146), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n198), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n204), .A2(new_n255), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT77), .B(KEYINPUT4), .Z(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n235), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n232), .B1(new_n248), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT80), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n221), .A2(new_n223), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n233), .B1(new_n265), .B2(new_n219), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n239), .A2(new_n240), .A3(new_n230), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(G104), .B1(new_n237), .B2(new_n238), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n221), .A2(new_n223), .ZN(new_n270));
  OAI21_X1  g084(.A(G101), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT80), .A3(new_n241), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT10), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n253), .A2(new_n210), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n274), .B1(new_n275), .B2(new_n206), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT81), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n271), .A2(KEYINPUT80), .A3(new_n241), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT80), .B1(new_n271), .B2(new_n241), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n276), .B(KEYINPUT81), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n263), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT11), .ZN(new_n283));
  INV_X1    g097(.A(G134), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(G137), .ZN(new_n285));
  INV_X1    g099(.A(G137), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT11), .A3(G134), .ZN(new_n287));
  INV_X1    g101(.A(G131), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n284), .A2(G137), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n285), .A2(new_n287), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT65), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n290), .A2(new_n291), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n287), .A2(new_n289), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(new_n285), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n285), .A2(new_n287), .A3(new_n294), .A4(new_n289), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G131), .ZN(new_n298));
  OAI22_X1  g112(.A1(new_n292), .A2(new_n293), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n282), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT81), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n280), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n285), .A2(new_n287), .A3(new_n289), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT66), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n297), .A2(G131), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n295), .A2(KEYINPUT65), .A3(new_n288), .A4(new_n285), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n290), .A2(new_n291), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n306), .A2(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n304), .A2(new_n310), .A3(new_n263), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n194), .B1(new_n300), .B2(new_n311), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n210), .A2(new_n253), .B1(new_n203), .B2(new_n205), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n268), .A2(new_n313), .A3(new_n272), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n215), .A2(new_n231), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n299), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT12), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT83), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n316), .A2(KEYINPUT12), .A3(new_n299), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT12), .B1(new_n316), .B2(new_n299), .ZN(new_n323));
  AOI211_X1 g137(.A(new_n318), .B(new_n310), .C1(new_n314), .C2(new_n315), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT83), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n322), .A2(new_n325), .A3(new_n311), .A4(new_n194), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT84), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n312), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n311), .A2(new_n194), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n329), .A2(KEYINPUT84), .A3(new_n322), .A4(new_n325), .ZN(new_n330));
  AOI211_X1 g144(.A(G469), .B(G902), .C1(new_n328), .C2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n194), .ZN(new_n332));
  AND3_X1   g146(.A1(new_n304), .A2(new_n310), .A3(new_n263), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n323), .A2(new_n324), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n311), .A2(KEYINPUT82), .A3(new_n194), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n300), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT82), .B1(new_n311), .B2(new_n194), .ZN(new_n338));
  OAI211_X1 g152(.A(G469), .B(new_n335), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(G469), .A2(G902), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n189), .B1(new_n331), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(G237), .A2(G953), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(G143), .A3(G214), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(G143), .B1(new_n343), .B2(G214), .ZN(new_n346));
  OAI21_X1  g160(.A(G131), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT17), .ZN(new_n348));
  INV_X1    g162(.A(G237), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n192), .A3(G214), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n199), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n288), .A3(new_n344), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n347), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT91), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT16), .ZN(new_n355));
  INV_X1    g169(.A(G140), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(G125), .ZN(new_n358));
  INV_X1    g172(.A(G125), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G140), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n357), .B1(new_n361), .B2(new_n355), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n197), .ZN(new_n363));
  OAI211_X1 g177(.A(G146), .B(new_n357), .C1(new_n361), .C2(new_n355), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT91), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n347), .A2(new_n366), .A3(new_n348), .A4(new_n352), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n347), .A2(new_n348), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n354), .A2(new_n365), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n345), .A2(new_n346), .ZN(new_n370));
  AND2_X1   g184(.A1(KEYINPUT18), .A2(G131), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n371), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n358), .A2(new_n360), .A3(new_n197), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT90), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n361), .A2(G146), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n361), .A2(KEYINPUT90), .A3(G146), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n374), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G113), .B(G122), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(new_n216), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n369), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n383), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n361), .B(KEYINPUT19), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n364), .B1(new_n386), .B2(G146), .ZN(new_n387));
  AND2_X1   g201(.A1(new_n347), .A2(new_n352), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI22_X1  g203(.A1(new_n372), .A2(new_n373), .B1(new_n378), .B2(new_n379), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n384), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G475), .ZN(new_n393));
  INV_X1    g207(.A(G902), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  XOR2_X1   g209(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT20), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n392), .A2(new_n399), .A3(new_n393), .A4(new_n394), .ZN(new_n400));
  INV_X1    g214(.A(new_n384), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n383), .B1(new_n369), .B2(new_n381), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n394), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n398), .A2(new_n400), .B1(G475), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G116), .B(G122), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G122), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(G116), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n222), .B1(new_n409), .B2(KEYINPUT14), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n407), .A2(new_n410), .B1(new_n227), .B2(new_n405), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT92), .B1(new_n195), .B2(G143), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT92), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n199), .A3(G128), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT93), .B1(new_n199), .B2(G128), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT93), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(new_n195), .A3(G143), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n415), .A2(new_n419), .A3(new_n284), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n284), .B1(new_n415), .B2(new_n419), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n411), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT94), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n411), .B(KEYINPUT94), .C1(new_n420), .C2(new_n421), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n227), .A2(new_n405), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n227), .A2(new_n405), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n420), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT13), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n419), .B1(new_n415), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT13), .B1(new_n412), .B2(new_n414), .ZN(new_n432));
  OAI21_X1  g246(.A(G134), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G217), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n188), .A2(new_n435), .A3(G953), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n426), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n426), .B2(new_n434), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n394), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT95), .ZN(new_n440));
  INV_X1    g254(.A(G478), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(KEYINPUT15), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT95), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n443), .B(new_n394), .C1(new_n437), .C2(new_n438), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n440), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n439), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(KEYINPUT15), .B2(new_n441), .ZN(new_n447));
  NAND2_X1  g261(.A1(G234), .A2(G237), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(G952), .A3(new_n192), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(G902), .A3(G953), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(G898), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AND4_X1   g269(.A1(new_n404), .A2(new_n445), .A3(new_n447), .A4(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G214), .B1(G237), .B2(G902), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G122), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT85), .ZN(new_n460));
  INV_X1    g274(.A(G119), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G116), .ZN(new_n462));
  INV_X1    g276(.A(G116), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G119), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(KEYINPUT2), .B(G113), .Z(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n462), .A2(new_n464), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT2), .B(G113), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT69), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n467), .A2(KEYINPUT69), .A3(new_n470), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n473), .A2(new_n474), .B1(new_n235), .B2(new_n261), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n248), .A2(new_n460), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n465), .A2(KEYINPUT5), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n477), .B(G113), .C1(KEYINPUT5), .C2(new_n462), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n273), .A2(new_n467), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n460), .B1(new_n248), .B2(new_n475), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n459), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n248), .A2(new_n475), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT85), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n484), .A2(new_n458), .A3(new_n479), .A4(new_n476), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(KEYINPUT6), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT68), .B1(new_n204), .B2(new_n196), .ZN(new_n487));
  AND4_X1   g301(.A1(KEYINPUT68), .A2(new_n196), .A3(new_n198), .A4(new_n200), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n208), .B1(new_n249), .B2(new_n251), .ZN(new_n489));
  OAI22_X1  g303(.A1(new_n487), .A2(new_n488), .B1(new_n489), .B2(new_n213), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT86), .B1(new_n490), .B2(G125), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n313), .A2(new_n492), .A3(new_n359), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n260), .A2(G125), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n192), .A2(G224), .ZN(new_n497));
  XOR2_X1   g311(.A(new_n496), .B(new_n497), .Z(new_n498));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n499), .B(new_n459), .C1(new_n480), .C2(new_n481), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n486), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n497), .B1(new_n502), .B2(KEYINPUT7), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n502), .B2(KEYINPUT7), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n494), .A2(KEYINPUT87), .B1(G125), .B2(new_n260), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT87), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n491), .A2(new_n493), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n504), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n458), .B(KEYINPUT8), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n478), .A2(new_n467), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n268), .B2(new_n272), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n231), .B1(new_n467), .B2(new_n478), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n509), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n494), .A2(KEYINPUT7), .A3(new_n495), .A4(new_n497), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(G902), .B1(new_n516), .B2(new_n485), .ZN(new_n517));
  OAI21_X1  g331(.A(G210), .B1(G237), .B2(G902), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n501), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n518), .B1(new_n501), .B2(new_n517), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n456), .B(new_n457), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n187), .B1(new_n342), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n521), .ZN(new_n523));
  INV_X1    g337(.A(new_n189), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n326), .A2(new_n327), .ZN(new_n525));
  INV_X1    g339(.A(new_n312), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n330), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G469), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n394), .ZN(new_n529));
  INV_X1    g343(.A(new_n341), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n524), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n523), .A2(new_n531), .A3(KEYINPUT96), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT25), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n363), .A2(new_n364), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT23), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n461), .B2(G128), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n536), .B(new_n537), .C1(G119), .C2(new_n195), .ZN(new_n538));
  XNOR2_X1  g352(.A(G119), .B(G128), .ZN(new_n539));
  XOR2_X1   g353(.A(KEYINPUT24), .B(G110), .Z(new_n540));
  AOI22_X1  g354(.A1(new_n538), .A2(G110), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n538), .A2(G110), .B1(new_n539), .B2(new_n540), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(new_n364), .A3(new_n375), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT71), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT22), .B(G137), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n542), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n542), .B2(new_n544), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n533), .B1(new_n551), .B2(G902), .ZN(new_n552));
  OAI211_X1 g366(.A(KEYINPUT25), .B(new_n394), .C1(new_n549), .C2(new_n550), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n435), .B1(G234), .B2(new_n394), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n554), .A2(KEYINPUT72), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT72), .B1(new_n554), .B2(new_n555), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n555), .A2(G902), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT73), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n556), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n343), .A2(G210), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n563), .B(KEYINPUT27), .Z(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT26), .B(G101), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n258), .A2(new_n259), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n299), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n474), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT69), .B1(new_n467), .B2(new_n470), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n286), .A2(G134), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n289), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n308), .A2(new_n309), .B1(G131), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n490), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n569), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT70), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT28), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n577), .B2(new_n579), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n574), .A2(G131), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n292), .B2(new_n293), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT67), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT67), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n575), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n587), .A3(new_n490), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n572), .B1(new_n588), .B2(new_n569), .ZN(new_n589));
  INV_X1    g403(.A(new_n577), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT28), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n567), .B1(new_n582), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT30), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n569), .B2(new_n576), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n308), .A2(new_n309), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n307), .A2(new_n306), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n260), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n313), .B1(new_n584), .B2(KEYINPUT67), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n598), .B2(new_n587), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n594), .B1(new_n599), .B2(new_n593), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n577), .B(new_n567), .C1(new_n600), .C2(new_n572), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT31), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n490), .B1(new_n575), .B2(new_n586), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n584), .A2(KEYINPUT67), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n593), .B(new_n569), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n569), .A2(new_n576), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT30), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n572), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n590), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(KEYINPUT31), .A3(new_n567), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n592), .B1(new_n603), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(G472), .A2(G902), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(KEYINPUT32), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n582), .A2(new_n591), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n566), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT31), .B1(new_n611), .B2(new_n567), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n572), .B1(new_n606), .B2(new_n608), .ZN(new_n620));
  NOR4_X1   g434(.A1(new_n620), .A2(new_n602), .A3(new_n590), .A4(new_n566), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n618), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT32), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n623), .A3(new_n614), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n572), .B1(new_n569), .B2(new_n576), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT28), .B1(new_n590), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n582), .A2(KEYINPUT29), .A3(new_n567), .A4(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n617), .A2(new_n566), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT29), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n611), .B2(new_n567), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n394), .B(new_n628), .C1(new_n629), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G472), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n562), .B1(new_n625), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n522), .A2(new_n532), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  OAI211_X1 g450(.A(new_n457), .B(new_n455), .C1(new_n519), .C2(new_n520), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n440), .A2(new_n441), .A3(new_n444), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n441), .A2(G902), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  INV_X1    g454(.A(new_n438), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n426), .A2(new_n434), .A3(new_n436), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT33), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n639), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n398), .A2(new_n400), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n403), .A2(G475), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n637), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(G472), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n622), .B2(new_n394), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n613), .A2(new_n615), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n651), .A2(new_n561), .A3(new_n531), .A4(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT34), .B(G104), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT97), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n656), .B(new_n658), .ZN(G6));
  NOR2_X1   g473(.A1(new_n342), .A2(new_n562), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n445), .A2(new_n447), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n395), .A2(new_n397), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n395), .A2(new_n397), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n648), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n637), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n660), .A2(new_n655), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT35), .B(G107), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  INV_X1    g483(.A(new_n557), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n554), .A2(KEYINPUT72), .A3(new_n555), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n548), .A2(KEYINPUT36), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n542), .A2(new_n544), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n559), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n670), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n522), .A2(new_n532), .A3(new_n655), .A4(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  AOI22_X1  g494(.A1(new_n616), .A2(new_n624), .B1(G472), .B2(new_n632), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n677), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n501), .A2(new_n517), .ZN(new_n684));
  INV_X1    g498(.A(new_n518), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n501), .A2(new_n517), .A3(new_n518), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n451), .A2(G900), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n449), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n648), .B(new_n690), .C1(new_n663), .C2(new_n664), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n662), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n688), .A2(new_n457), .A3(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n683), .A2(new_n342), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n195), .ZN(G30));
  XNOR2_X1  g509(.A(new_n690), .B(KEYINPUT39), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n531), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT40), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT98), .ZN(new_n699));
  INV_X1    g513(.A(new_n601), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n590), .A2(new_n626), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n701), .A2(new_n567), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n699), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n601), .B(KEYINPUT98), .C1(new_n567), .C2(new_n701), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n394), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G472), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n677), .B1(new_n625), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n519), .A2(new_n520), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT38), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT38), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n710), .B1(new_n519), .B2(new_n520), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n457), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n662), .A2(new_n404), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n698), .A2(new_n707), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G143), .ZN(G45));
  NAND3_X1  g532(.A1(new_n646), .A2(new_n649), .A3(new_n690), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT99), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n646), .A2(new_n649), .A3(KEYINPUT99), .A4(new_n690), .ZN(new_n722));
  AND4_X1   g536(.A1(new_n457), .A2(new_n688), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n677), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n681), .A2(new_n724), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n723), .A2(new_n725), .A3(new_n531), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n197), .ZN(G48));
  NAND2_X1  g541(.A1(new_n527), .A2(new_n394), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT100), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n528), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n527), .B(new_n394), .C1(new_n729), .C2(new_n528), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n189), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT101), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT101), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n731), .A2(new_n735), .A3(new_n732), .A4(new_n189), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n734), .A2(new_n634), .A3(new_n651), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT102), .ZN(new_n738));
  XNOR2_X1  g552(.A(KEYINPUT41), .B(G113), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G15));
  NAND4_X1  g554(.A1(new_n734), .A2(new_n634), .A3(new_n666), .A4(new_n736), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G116), .ZN(G18));
  INV_X1    g556(.A(new_n456), .ZN(new_n743));
  NOR3_X1   g557(.A1(new_n681), .A2(new_n743), .A3(new_n724), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n708), .A2(new_n713), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n734), .A2(new_n744), .A3(new_n745), .A4(new_n736), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT103), .B(G119), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G21));
  AND2_X1   g562(.A1(new_n582), .A2(new_n627), .ZN(new_n749));
  OAI22_X1  g563(.A1(new_n619), .A2(new_n621), .B1(new_n749), .B2(new_n567), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n614), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n603), .A2(new_n612), .ZN(new_n752));
  AOI21_X1  g566(.A(G902), .B1(new_n752), .B2(new_n618), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n751), .B(new_n561), .C1(new_n753), .C2(new_n652), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n754), .A2(new_n637), .A3(new_n715), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n734), .A2(new_n755), .A3(new_n736), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G122), .ZN(G24));
  NAND2_X1  g571(.A1(new_n721), .A2(new_n722), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n751), .B(new_n677), .C1(new_n753), .C2(new_n652), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n734), .A2(new_n745), .A3(new_n736), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  NAND2_X1  g576(.A1(new_n311), .A2(new_n194), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT82), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n300), .A3(new_n336), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT104), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n335), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g582(.A(KEYINPUT104), .B(new_n332), .C1(new_n333), .C2(new_n334), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n766), .A2(new_n768), .A3(G469), .A4(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n340), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n524), .B1(new_n771), .B2(new_n529), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n686), .A2(new_n457), .A3(new_n687), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT105), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n708), .A2(KEYINPUT105), .A3(new_n457), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n634), .A2(new_n772), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n758), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(KEYINPUT42), .A3(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT42), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n634), .A2(new_n772), .A3(new_n775), .A4(new_n776), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n780), .B1(new_n781), .B2(new_n758), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  INV_X1    g598(.A(new_n692), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n284), .ZN(G36));
  NAND2_X1  g601(.A1(new_n766), .A2(new_n335), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n766), .A2(new_n768), .A3(KEYINPUT45), .A4(new_n769), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(G469), .A3(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n792), .A2(new_n340), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n793), .A2(KEYINPUT46), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(KEYINPUT46), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n794), .A2(new_n529), .A3(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(new_n189), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n797), .A2(new_n696), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n776), .A2(new_n775), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n646), .A2(new_n404), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(KEYINPUT43), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(KEYINPUT43), .ZN(new_n802));
  OR4_X1    g616(.A1(new_n655), .A2(new_n801), .A3(new_n802), .A4(new_n724), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n799), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n804), .B2(new_n803), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n798), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(KEYINPUT106), .B(G137), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n807), .B(new_n808), .ZN(G39));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(KEYINPUT107), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n796), .A2(new_n189), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n796), .B2(new_n189), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n682), .A2(new_n758), .A3(new_n561), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n814), .A2(new_n799), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  NOR4_X1   g634(.A1(new_n562), .A2(new_n800), .A3(new_n524), .A4(new_n713), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT108), .Z(new_n822));
  NAND2_X1  g636(.A1(new_n731), .A2(new_n732), .ZN(new_n823));
  XOR2_X1   g637(.A(new_n823), .B(KEYINPUT49), .Z(new_n824));
  NAND2_X1  g638(.A1(new_n625), .A2(new_n706), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n822), .A2(new_n824), .A3(new_n826), .A4(new_n712), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n801), .A2(new_n802), .A3(new_n449), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n799), .A2(new_n734), .A3(new_n736), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n634), .ZN(new_n830));
  XOR2_X1   g644(.A(KEYINPUT121), .B(KEYINPUT48), .Z(new_n831));
  OR3_X1    g645(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n831), .B1(new_n829), .B2(new_n830), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n825), .A2(new_n562), .A3(new_n449), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n799), .A3(new_n734), .A4(new_n736), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n835), .A2(new_n650), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n192), .A2(G952), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n734), .A2(new_n745), .A3(new_n736), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n754), .A2(new_n801), .A3(new_n802), .A4(new_n449), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n832), .A2(new_n833), .A3(new_n836), .A4(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n823), .A2(new_n189), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT114), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n813), .B2(new_n816), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(new_n799), .A3(new_n839), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n457), .B1(new_n709), .B2(new_n711), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n734), .A2(new_n736), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT115), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n734), .A2(new_n846), .A3(new_n849), .A4(new_n736), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n839), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n851), .A2(KEYINPUT117), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(KEYINPUT50), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT50), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n853), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n835), .A2(new_n649), .A3(new_n646), .ZN(new_n860));
  OR3_X1    g674(.A1(new_n829), .A2(KEYINPUT118), .A3(new_n759), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT118), .B1(new_n829), .B2(new_n759), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n845), .A2(new_n857), .A3(new_n859), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n841), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n635), .A2(new_n656), .A3(new_n756), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n746), .A2(new_n741), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT109), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n661), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n445), .A2(new_n447), .A3(KEYINPUT109), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n649), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n637), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n660), .A2(new_n655), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT110), .B1(new_n678), .B2(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n678), .A2(KEYINPUT110), .A3(new_n876), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n869), .B(new_n738), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  INV_X1    g695(.A(new_n693), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n725), .B(new_n531), .C1(new_n723), .C2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n688), .A2(new_n714), .A3(new_n457), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(new_n707), .A3(new_n772), .A4(new_n690), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n761), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT52), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT52), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n761), .A2(new_n883), .A3(new_n889), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n881), .B1(new_n891), .B2(KEYINPUT112), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n772), .A2(new_n775), .A3(new_n776), .ZN(new_n893));
  AOI22_X1  g707(.A1(new_n777), .A2(new_n692), .B1(new_n893), .B2(new_n760), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT111), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n871), .A2(new_n872), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n691), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n531), .A2(new_n776), .A3(new_n775), .A4(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n895), .B1(new_n898), .B2(new_n683), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n529), .A2(new_n530), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n897), .A2(new_n900), .A3(new_n189), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n799), .A2(new_n901), .A3(KEYINPUT111), .A4(new_n725), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT42), .B1(new_n777), .B2(new_n778), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n781), .A2(new_n780), .A3(new_n758), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n894), .B(new_n903), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n891), .A2(new_n906), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n880), .A2(new_n892), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n892), .B1(new_n880), .B2(new_n907), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT54), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n878), .A2(new_n877), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n756), .A2(new_n656), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(new_n635), .A3(new_n741), .A4(new_n746), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT102), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n737), .B(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n907), .A2(new_n881), .A3(new_n913), .A4(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n760), .A2(new_n775), .A3(new_n776), .A4(new_n772), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n781), .B2(new_n785), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n899), .B2(new_n902), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(new_n888), .A3(new_n783), .A4(new_n890), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT53), .B1(new_n879), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n912), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n866), .A2(new_n910), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n856), .A2(KEYINPUT50), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT117), .B1(new_n851), .B2(new_n852), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n859), .B(new_n863), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(KEYINPUT119), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n857), .A2(new_n933), .A3(new_n859), .A4(new_n863), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n842), .B1(new_n814), .B2(new_n817), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n839), .A2(new_n799), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT51), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n928), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  AOI211_X1 g754(.A(KEYINPUT120), .B(new_n938), .C1(new_n932), .C2(new_n934), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n927), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(G952), .A2(G953), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n827), .B1(new_n942), .B2(new_n943), .ZN(G75));
  INV_X1    g758(.A(new_n924), .ZN(new_n945));
  NOR3_X1   g759(.A1(new_n879), .A2(new_n923), .A3(KEYINPUT53), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n947), .A2(G210), .A3(G902), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT56), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n486), .A2(new_n500), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(new_n498), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT55), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n948), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n948), .B2(new_n949), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n192), .A2(G952), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(G51));
  XOR2_X1   g770(.A(new_n340), .B(KEYINPUT57), .Z(new_n957));
  AND3_X1   g771(.A1(new_n919), .A2(new_n924), .A3(new_n912), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n957), .B1(new_n958), .B2(new_n925), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT122), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  OAI211_X1 g775(.A(new_n961), .B(new_n957), .C1(new_n958), .C2(new_n925), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n527), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n792), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n947), .A2(G902), .A3(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n955), .B1(new_n963), .B2(new_n965), .ZN(G54));
  NAND4_X1  g780(.A1(new_n947), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n967));
  INV_X1    g781(.A(new_n392), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n969), .A2(new_n970), .A3(new_n955), .ZN(G60));
  OR2_X1    g785(.A1(new_n643), .A2(new_n644), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n910), .A2(new_n926), .ZN(new_n973));
  NAND2_X1  g787(.A1(G478), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT59), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n972), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n972), .B(new_n975), .C1(new_n958), .C2(new_n925), .ZN(new_n977));
  INV_X1    g791(.A(new_n955), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n976), .A2(new_n979), .ZN(G63));
  NAND2_X1  g794(.A1(G217), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT60), .Z(new_n982));
  NAND4_X1  g796(.A1(new_n919), .A2(new_n924), .A3(new_n674), .A4(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT123), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  OAI21_X1  g800(.A(KEYINPUT124), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n919), .A2(new_n924), .A3(new_n982), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n955), .B1(new_n988), .B2(new_n551), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(new_n985), .B2(new_n986), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT61), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n987), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  OAI221_X1 g806(.A(new_n989), .B1(KEYINPUT124), .B2(KEYINPUT61), .C1(new_n985), .C2(new_n986), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(G66));
  XNOR2_X1  g808(.A(new_n879), .B(KEYINPUT125), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n192), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n995), .A2(KEYINPUT126), .A3(new_n192), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(G224), .ZN(new_n1001));
  OAI21_X1  g815(.A(G953), .B1(new_n453), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n192), .A2(G898), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n950), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1000), .A2(new_n950), .A3(new_n1004), .A4(new_n1002), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(G69));
  NAND3_X1  g822(.A1(new_n717), .A2(new_n761), .A3(new_n883), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n874), .A2(new_n650), .ZN(new_n1011));
  AND4_X1   g825(.A1(new_n634), .A2(new_n697), .A3(new_n799), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(new_n798), .B2(new_n806), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1010), .A2(new_n1013), .A3(new_n819), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n192), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n609), .B(new_n386), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT127), .Z(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1017), .B1(G900), .B2(G953), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n786), .B1(new_n798), .B2(new_n806), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n761), .A2(new_n883), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n830), .A2(new_n884), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1022), .B1(new_n798), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1021), .A2(new_n1024), .A3(new_n783), .A4(new_n819), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1020), .B1(new_n1025), .B2(G953), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1019), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n192), .B1(G227), .B2(G900), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1027), .B(new_n1028), .ZN(G72));
  NAND2_X1  g843(.A1(G472), .A2(G902), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT63), .Z(new_n1031));
  OAI21_X1  g845(.A(new_n1031), .B1(new_n1015), .B2(new_n995), .ZN(new_n1032));
  OAI211_X1 g846(.A(new_n1032), .B(new_n567), .C1(new_n590), .C2(new_n620), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n611), .A2(new_n567), .ZN(new_n1034));
  OAI221_X1 g848(.A(new_n1031), .B1(new_n700), .B2(new_n1034), .C1(new_n908), .C2(new_n909), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1031), .B1(new_n1025), .B2(new_n995), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1036), .A2(new_n566), .A3(new_n611), .ZN(new_n1037));
  AND4_X1   g851(.A1(new_n978), .A2(new_n1033), .A3(new_n1035), .A4(new_n1037), .ZN(G57));
endmodule


