//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n558, new_n559, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND3_X1   g035(.A1(KEYINPUT67), .A2(G113), .A3(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(KEYINPUT67), .B1(G113), .B2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n460), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n460), .C1(new_n464), .C2(new_n465), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n460), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  OAI21_X1  g047(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G112), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT69), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n464), .A2(new_n465), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n476), .B1(G136), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(KEYINPUT68), .B1(new_n477), .B2(new_n460), .ZN(new_n480));
  XNOR2_X1  g055(.A(KEYINPUT3), .B(G2104), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n481), .A2(new_n482), .A3(G2105), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n495), .B1(new_n464), .B2(new_n465), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n495), .B(new_n498), .C1(new_n465), .C2(new_n464), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n493), .B1(new_n497), .B2(new_n499), .ZN(G164));
  NAND2_X1  g075(.A1(KEYINPUT70), .A2(G651), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n504));
  OR2_X1    g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G88), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n509), .B1(new_n505), .B2(new_n506), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g087(.A(G651), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  AND3_X1   g088(.A1(KEYINPUT70), .A2(KEYINPUT6), .A3(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT6), .B1(KEYINPUT70), .B2(G651), .ZN(new_n515));
  OAI211_X1 g090(.A(G50), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n508), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(G166));
  NAND2_X1  g093(.A1(new_n507), .A2(G89), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n520), .B1(new_n503), .B2(new_n504), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G51), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n505), .A2(new_n506), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n526));
  AND4_X1   g101(.A1(new_n519), .A2(new_n522), .A3(new_n524), .A4(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  INV_X1    g103(.A(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT71), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n507), .A2(G90), .B1(new_n521), .B2(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(KEYINPUT71), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(G171));
  NAND2_X1  g110(.A1(new_n507), .A2(G81), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n521), .A2(G43), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n525), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n536), .B(new_n537), .C1(new_n529), .C2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G860), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n539), .A2(new_n540), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  INV_X1    g120(.A(G65), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n546), .B1(new_n505), .B2(new_n506), .ZN(new_n547));
  AND2_X1   g122(.A1(G78), .A2(G543), .ZN(new_n548));
  OAI21_X1  g123(.A(G651), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g124(.A(G53), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT9), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n503), .A2(new_n504), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n553), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n553), .A2(new_n525), .A3(G91), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n549), .A2(new_n552), .A3(new_n554), .A4(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n558));
  XNOR2_X1  g133(.A(G168), .B(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(G286));
  AND2_X1   g135(.A1(KEYINPUT5), .A2(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(KEYINPUT5), .A2(G543), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n514), .A2(new_n515), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G88), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n516), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(G62), .B1(new_n561), .B2(new_n562), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n529), .B1(new_n566), .B2(new_n511), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT73), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n508), .A2(new_n513), .A3(new_n569), .A4(new_n516), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n568), .A2(new_n570), .ZN(G303));
  OAI211_X1 g146(.A(KEYINPUT75), .B(G651), .C1(new_n525), .C2(G74), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n573));
  NAND2_X1  g148(.A1(G74), .A2(G651), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n561), .A2(new_n562), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n573), .B(new_n574), .C1(new_n575), .C2(new_n529), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n572), .A2(new_n576), .B1(new_n521), .B2(G49), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n507), .A2(new_n578), .A3(G87), .ZN(new_n579));
  INV_X1    g154(.A(G87), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT74), .B1(new_n563), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n577), .A2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n575), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(new_n507), .B2(G86), .ZN(new_n587));
  OAI211_X1 g162(.A(G48), .B(G543), .C1(new_n514), .C2(new_n515), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT76), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n553), .A2(new_n590), .A3(G48), .A4(G543), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n587), .A2(new_n592), .ZN(G305));
  NAND2_X1  g168(.A1(new_n507), .A2(G85), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n521), .A2(G47), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n594), .B(new_n595), .C1(new_n529), .C2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n507), .A2(KEYINPUT10), .A3(G92), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n563), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n575), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(G54), .B2(new_n521), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT77), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n598), .B1(G868), .B2(new_n610), .ZN(G284));
  OAI21_X1  g186(.A(new_n598), .B1(G868), .B2(new_n610), .ZN(G321));
  NOR2_X1   g187(.A1(G299), .A2(G868), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n559), .B2(G868), .ZN(G297));
  AOI21_X1  g189(.A(new_n613), .B1(new_n559), .B2(G868), .ZN(G280));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n610), .B1(new_n616), .B2(G860), .ZN(G148));
  NAND2_X1  g192(.A1(new_n610), .A2(new_n616), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  OR3_X1    g195(.A1(new_n619), .A2(KEYINPUT78), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(KEYINPUT78), .B1(new_n619), .B2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n539), .A2(new_n620), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(G323));
  XOR2_X1   g199(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n625));
  XNOR2_X1  g200(.A(G323), .B(new_n625), .ZN(G282));
  NAND2_X1  g201(.A1(new_n481), .A2(new_n469), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT13), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n484), .A2(G123), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n478), .A2(G135), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n460), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n631), .A2(G2100), .B1(G2096), .B2(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n637), .B(new_n638), .C1(G2100), .C2(new_n631), .ZN(G156));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n644), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n647), .B2(new_n646), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n643), .B(new_n649), .Z(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  AND3_X1   g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(KEYINPUT81), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT17), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT82), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n661), .B(new_n663), .C1(new_n660), .C2(new_n656), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n656), .A2(new_n658), .A3(new_n662), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT18), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n659), .A2(new_n662), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n664), .B(new_n666), .C1(new_n657), .C2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2096), .B(G2100), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1961), .B(G1966), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT20), .ZN(new_n678));
  INV_X1    g253(.A(new_n673), .ZN(new_n679));
  INV_X1    g254(.A(new_n676), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n675), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n678), .B(new_n682), .C1(new_n679), .C2(new_n681), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT84), .Z(new_n684));
  XOR2_X1   g259(.A(G1981), .B(G1986), .Z(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n684), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G35), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G162), .B2(new_n692), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G2090), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(G32), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n469), .A2(G105), .ZN(new_n698));
  NAND3_X1  g273(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT26), .ZN(new_n700));
  AOI211_X1 g275(.A(new_n698), .B(new_n700), .C1(G141), .C2(new_n478), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n484), .A2(G129), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n697), .B1(new_n703), .B2(new_n692), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT27), .B(G1996), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n706), .ZN(new_n708));
  NOR2_X1   g283(.A1(G29), .A2(G33), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT91), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT92), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT25), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n478), .A2(G139), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n713), .B(new_n714), .C1(new_n460), .C2(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n710), .B1(new_n716), .B2(new_n692), .ZN(new_n717));
  INV_X1    g292(.A(G2072), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n696), .A2(new_n707), .A3(new_n708), .A4(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G34), .ZN(new_n721));
  AOI21_X1  g296(.A(G29), .B1(new_n721), .B2(KEYINPUT24), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(KEYINPUT24), .B2(new_n721), .ZN(new_n723));
  INV_X1    g298(.A(G160), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n692), .ZN(new_n725));
  INV_X1    g300(.A(G2084), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT95), .ZN(new_n728));
  INV_X1    g303(.A(G28), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(KEYINPUT30), .ZN(new_n730));
  AOI21_X1  g305(.A(G29), .B1(new_n729), .B2(KEYINPUT30), .ZN(new_n731));
  OR2_X1    g306(.A1(KEYINPUT31), .A2(G11), .ZN(new_n732));
  NAND2_X1  g307(.A1(KEYINPUT31), .A2(G11), .ZN(new_n733));
  AOI22_X1  g308(.A1(new_n730), .A2(new_n731), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n636), .B2(new_n692), .ZN(new_n735));
  INV_X1    g310(.A(G2078), .ZN(new_n736));
  NAND2_X1  g311(.A1(G164), .A2(G29), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G27), .B2(G29), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n739), .B1(new_n736), .B2(new_n738), .C1(new_n726), .C2(new_n725), .ZN(new_n740));
  MUX2_X1   g315(.A(G19), .B(new_n539), .S(G16), .Z(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(G1341), .Z(new_n742));
  OR2_X1    g317(.A1(new_n717), .A2(new_n718), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n742), .B1(new_n744), .B2(KEYINPUT93), .ZN(new_n745));
  NOR4_X1   g320(.A1(new_n720), .A2(new_n728), .A3(new_n740), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n692), .A2(G26), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT28), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n484), .A2(G128), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G116), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G2105), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n478), .B2(G140), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(G29), .ZN(new_n755));
  INV_X1    g330(.A(G2067), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n744), .B2(KEYINPUT93), .ZN(new_n758));
  INV_X1    g333(.A(G16), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G4), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n610), .B2(new_n759), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(G1348), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n759), .A2(G5), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G171), .B2(new_n759), .ZN(new_n764));
  INV_X1    g339(.A(G1961), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n758), .A2(new_n762), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G1348), .B2(new_n761), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n695), .A2(G2090), .ZN(new_n769));
  NAND2_X1  g344(.A1(G299), .A2(G16), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n759), .A2(G20), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT23), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1956), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n759), .A2(G21), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G168), .B2(new_n759), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT94), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1966), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n746), .A2(new_n768), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n780), .A2(KEYINPUT96), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(KEYINPUT96), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n692), .A2(G25), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n484), .A2(G119), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n785));
  INV_X1    g360(.A(G107), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G2105), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n478), .B2(G131), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n783), .B1(new_n790), .B2(new_n692), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT35), .B(G1991), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  MUX2_X1   g368(.A(G24), .B(G290), .S(G16), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT85), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1986), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n759), .A2(G22), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT88), .Z(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G166), .B2(new_n759), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT89), .B(G1971), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(G6), .A2(G16), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G305), .B2(new_n759), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT32), .B(G1981), .Z(new_n804));
  OAI21_X1  g379(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g380(.A1(new_n759), .A2(G23), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G288), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT33), .B(G1976), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT87), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n807), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n803), .A2(new_n804), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n805), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n793), .B(new_n796), .C1(new_n815), .C2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT90), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n815), .A2(new_n817), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(KEYINPUT36), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n819), .A2(new_n823), .A3(new_n820), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n781), .A2(new_n782), .B1(new_n822), .B2(new_n824), .ZN(G311));
  NAND2_X1  g400(.A1(new_n781), .A2(new_n782), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(new_n824), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(G150));
  NAND2_X1  g403(.A1(new_n507), .A2(G93), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n521), .A2(G55), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n829), .B(new_n830), .C1(new_n529), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G860), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT98), .B(KEYINPUT37), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n610), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n539), .B(new_n832), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(KEYINPUT97), .Z(new_n842));
  OAI21_X1  g417(.A(new_n540), .B1(new_n840), .B2(KEYINPUT39), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n835), .B1(new_n842), .B2(new_n843), .ZN(G145));
  XNOR2_X1  g419(.A(new_n486), .B(new_n636), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(new_n724), .ZN(new_n846));
  XNOR2_X1  g421(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n846), .B(new_n847), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n703), .B(new_n754), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n497), .A2(new_n499), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n488), .A2(new_n492), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT101), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n716), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n849), .A2(new_n852), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n716), .A2(new_n854), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n478), .A2(G142), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n460), .A2(G118), .ZN(new_n860));
  OAI21_X1  g435(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(G130), .B2(new_n484), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n858), .B(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n789), .B(new_n629), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n857), .A2(new_n864), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT102), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n866), .B1(new_n865), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n848), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  INV_X1    g447(.A(new_n848), .ZN(new_n873));
  NAND4_X1  g448(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT102), .A4(new_n868), .ZN(new_n874));
  INV_X1    g449(.A(G37), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n618), .B(new_n838), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n603), .A2(new_n607), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n880), .A2(G299), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n881), .A2(KEYINPUT103), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(G299), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(KEYINPUT103), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n879), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(KEYINPUT104), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n885), .B(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n879), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n886), .A2(KEYINPUT104), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n888), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(G290), .B(KEYINPUT105), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n895), .A2(G288), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(G288), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G305), .B(new_n517), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n896), .B2(new_n897), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT42), .B1(new_n900), .B2(new_n902), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n878), .B1(new_n894), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT106), .ZN(new_n910));
  INV_X1    g485(.A(new_n893), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n890), .A2(new_n891), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n887), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n910), .B1(new_n913), .B2(new_n907), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n894), .A2(KEYINPUT106), .A3(new_n908), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(KEYINPUT107), .A3(new_n907), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n909), .A2(new_n914), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n917), .A2(new_n918), .A3(G868), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n832), .A2(new_n620), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT108), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n921), .B1(new_n917), .B2(G868), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n919), .A2(new_n922), .ZN(G295));
  NOR2_X1   g498(.A1(new_n919), .A2(new_n922), .ZN(G331));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n925));
  OR2_X1    g500(.A1(G171), .A2(G168), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n559), .A2(G171), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n926), .A2(new_n927), .A3(new_n838), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n838), .B1(new_n926), .B2(new_n927), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n885), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n930), .A2(KEYINPUT110), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n928), .A2(new_n929), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n890), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n903), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(KEYINPUT110), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n931), .A2(new_n933), .A3(new_n934), .A4(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n933), .A2(new_n930), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n936), .B(new_n875), .C1(new_n937), .C2(new_n934), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n931), .A2(new_n933), .A3(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n903), .ZN(new_n941));
  XOR2_X1   g516(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n942));
  NAND4_X1  g517(.A1(new_n941), .A2(new_n875), .A3(new_n942), .A4(new_n936), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n925), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(new_n875), .A3(new_n936), .ZN(new_n945));
  INV_X1    g520(.A(new_n942), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n938), .A2(new_n946), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n944), .B1(new_n949), .B2(new_n925), .ZN(G397));
  XNOR2_X1  g525(.A(new_n754), .B(new_n756), .ZN(new_n951));
  INV_X1    g526(.A(G1996), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n952), .B2(new_n703), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(G164), .B2(G1384), .ZN(new_n955));
  INV_X1    g530(.A(new_n467), .ZN(new_n956));
  INV_X1    g531(.A(new_n471), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n956), .A2(G40), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n953), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n952), .A3(new_n703), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n961), .A2(KEYINPUT111), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(KEYINPUT111), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT112), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n789), .B(new_n792), .ZN(new_n967));
  OR2_X1    g542(.A1(new_n967), .A2(KEYINPUT113), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(KEYINPUT113), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n968), .A2(new_n959), .A3(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT126), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT126), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n966), .A2(new_n973), .A3(new_n970), .ZN(new_n974));
  NOR2_X1   g549(.A1(G290), .A2(G1986), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n959), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT48), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n972), .A2(new_n974), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n951), .A2(new_n703), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n959), .A2(new_n952), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n979), .A2(new_n959), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n980), .B2(new_n981), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n983), .B(KEYINPUT47), .Z(new_n984));
  NAND2_X1  g559(.A1(new_n790), .A2(new_n792), .ZN(new_n985));
  OAI22_X1  g560(.A1(new_n965), .A2(new_n985), .B1(G2067), .B2(new_n754), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n986), .B2(new_n959), .ZN(new_n987));
  AND2_X1   g562(.A1(new_n978), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1981), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n587), .A2(new_n989), .A3(new_n592), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(KEYINPUT114), .ZN(new_n991));
  NOR2_X1   g566(.A1(G288), .A2(G1976), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n992), .B(KEYINPUT115), .Z(new_n993));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n587), .A2(new_n989), .A3(new_n592), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n989), .B1(new_n587), .B2(new_n592), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(G305), .A2(G1981), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n998), .A2(KEYINPUT49), .A3(new_n990), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n850), .B2(new_n851), .ZN(new_n1001));
  INV_X1    g576(.A(G40), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n467), .A2(new_n471), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1000), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n997), .A2(new_n999), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n991), .B1(new_n993), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1004), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n568), .A2(new_n570), .A3(G8), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n568), .A2(new_n570), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  INV_X1    g588(.A(new_n499), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n498), .B1(new_n481), .B2(new_n495), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1013), .B1(new_n1016), .B2(new_n493), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n958), .B1(new_n1017), .B2(new_n954), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n852), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1971), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G2090), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n852), .A2(new_n1023), .A3(new_n1013), .ZN(new_n1024));
  AND4_X1   g599(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .A4(new_n1003), .ZN(new_n1025));
  OAI211_X1 g600(.A(G8), .B(new_n1012), .C1(new_n1020), .C2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n577), .A2(new_n582), .A3(G1976), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1004), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1029));
  INV_X1    g604(.A(G1976), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(G288), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(new_n1004), .A3(new_n1027), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1005), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  OAI22_X1  g608(.A1(new_n1006), .A2(new_n1007), .B1(new_n1026), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G1971), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1003), .B1(new_n1001), .B2(KEYINPUT45), .ZN(new_n1036));
  NOR3_X1   g611(.A1(G164), .A2(new_n954), .A3(G1384), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1022), .A2(new_n1024), .A3(new_n1021), .A4(new_n1003), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1000), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1033), .B1(new_n1012), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1003), .B1(new_n1001), .B2(new_n1023), .ZN(new_n1042));
  NOR3_X1   g617(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n955), .A2(new_n1019), .A3(new_n1003), .ZN(new_n1045));
  INV_X1    g620(.A(G1966), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1044), .A2(new_n726), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n559), .A2(G8), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT117), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1022), .A2(new_n1024), .A3(new_n726), .A4(new_n1003), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1052), .A2(new_n1053), .A3(G8), .A4(new_n559), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1012), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1038), .A2(KEYINPUT116), .A3(new_n1039), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G8), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT116), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1056), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1041), .A2(new_n1055), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT118), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT63), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1041), .A2(new_n1055), .A3(new_n1060), .A4(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1040), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1063), .B1(new_n1067), .B2(new_n1056), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1041), .A2(new_n1055), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1034), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n1004), .B2(new_n1027), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1028), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1073), .B2(new_n1031), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1026), .A2(new_n1005), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(G8), .A3(new_n1057), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1075), .B1(new_n1056), .B2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1045), .B2(G2078), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1018), .A2(KEYINPUT53), .A3(new_n736), .A4(new_n1019), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1022), .A2(new_n1024), .A3(new_n1003), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n765), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1082), .A2(KEYINPUT123), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(KEYINPUT123), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1086));
  OAI211_X1 g661(.A(G301), .B(new_n1081), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1081), .A2(new_n1084), .A3(new_n1082), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(G171), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1050), .A2(G168), .A3(new_n1051), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G8), .ZN(new_n1093));
  AOI21_X1  g668(.A(G168), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT51), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1092), .A2(new_n1096), .A3(G8), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1079), .A2(new_n1091), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1081), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G171), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1089), .A2(G171), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT54), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT119), .B(G1956), .Z(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1107));
  AND3_X1   g682(.A1(G299), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n1108));
  NOR2_X1   g683(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1109));
  NAND2_X1  g684(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NOR3_X1   g686(.A1(G299), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n955), .A2(new_n1019), .A3(new_n1003), .A4(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1107), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n610), .ZN(new_n1117));
  INV_X1    g692(.A(G1348), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1083), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1001), .A2(new_n1003), .A3(new_n756), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1117), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1113), .B1(new_n1107), .B2(new_n1115), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1116), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1107), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1125), .B2(new_n1122), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1107), .A2(new_n1115), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1113), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(KEYINPUT61), .A3(new_n1116), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n955), .A2(new_n1019), .A3(new_n952), .A4(new_n1003), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  AOI22_X1  g709(.A1(new_n1131), .A2(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1018), .A2(KEYINPUT121), .A3(new_n952), .A4(new_n1019), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n539), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1126), .B(new_n1130), .C1(KEYINPUT59), .C2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1119), .A2(KEYINPUT60), .A3(new_n1120), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(new_n1117), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1119), .A2(new_n610), .A3(KEYINPUT60), .A4(new_n1120), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1137), .A2(KEYINPUT59), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1123), .B1(new_n1138), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT122), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1150), .B(new_n1123), .C1(new_n1138), .C2(new_n1147), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1104), .A2(new_n1149), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1070), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1153), .B1(new_n1070), .B2(new_n1152), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1098), .A2(KEYINPUT62), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1079), .A2(G171), .A3(new_n1100), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1098), .A2(KEYINPUT62), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1154), .A2(new_n1155), .A3(new_n1159), .ZN(new_n1160));
  AND2_X1   g735(.A1(G290), .A2(G1986), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n959), .B1(new_n975), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n966), .A2(new_n1162), .A3(new_n970), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n988), .B1(new_n1160), .B2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g739(.A(G319), .ZN(new_n1166));
  NOR4_X1   g740(.A1(G229), .A2(new_n1166), .A3(G401), .A4(G227), .ZN(new_n1167));
  OAI211_X1 g741(.A(new_n876), .B(new_n1167), .C1(new_n947), .C2(new_n948), .ZN(G225));
  INV_X1    g742(.A(G225), .ZN(G308));
endmodule


