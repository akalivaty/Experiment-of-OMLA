//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G227), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G953), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G137), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(G137), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT11), .A3(G134), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G131), .ZN(new_n198));
  INV_X1    g012(.A(G131), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n193), .A2(new_n196), .A3(new_n199), .A4(new_n194), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(new_n202), .B2(G107), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT86), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT86), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n205), .B(KEYINPUT3), .C1(new_n202), .C2(G107), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n208));
  INV_X1    g022(.A(G107), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT87), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT87), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n212), .A2(new_n208), .A3(new_n209), .A4(G104), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(G104), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n207), .A2(new_n214), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n202), .A2(G107), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n219), .B2(new_n216), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT64), .B(G146), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT1), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G128), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n223), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G143), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(new_n223), .B2(G146), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(new_n222), .B2(new_n223), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n227), .A2(KEYINPUT64), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n227), .A2(KEYINPUT64), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n231), .B(G143), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT1), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G128), .ZN(new_n239));
  AND3_X1   g053(.A1(new_n221), .A2(new_n230), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G128), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n233), .A2(new_n236), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n221), .B1(new_n239), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n201), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT12), .B1(new_n201), .B2(KEYINPUT88), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n201), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n233), .B2(new_n236), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n250), .A2(new_n238), .B1(new_n225), .B2(new_n229), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n221), .ZN(new_n252));
  AOI211_X1 g066(.A(KEYINPUT1), .B(new_n249), .C1(new_n233), .C2(new_n236), .ZN(new_n253));
  INV_X1    g067(.A(new_n243), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n218), .B(new_n220), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n248), .B1(new_n252), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n246), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n247), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT10), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n239), .B2(new_n230), .ZN(new_n261));
  INV_X1    g075(.A(new_n221), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n255), .A2(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n214), .A2(new_n217), .ZN(new_n264));
  INV_X1    g078(.A(new_n207), .ZN(new_n265));
  OAI21_X1  g079(.A(G101), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n266), .A2(KEYINPUT4), .A3(new_n218), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n237), .A2(new_n269), .ZN(new_n270));
  OR2_X1    g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n229), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n274), .B(G101), .C1(new_n264), .C2(new_n265), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n267), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n263), .A2(new_n248), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n190), .B1(new_n259), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n190), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n248), .B1(new_n263), .B2(new_n276), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT89), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n256), .A2(new_n257), .ZN(new_n284));
  AOI211_X1 g098(.A(new_n248), .B(new_n246), .C1(new_n252), .C2(new_n255), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n277), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n190), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n255), .A2(new_n260), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n261), .A2(new_n262), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n276), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n201), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n292), .A2(new_n277), .A3(new_n190), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT89), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n288), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n282), .A2(new_n283), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT90), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n296), .A2(new_n297), .A3(G469), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n296), .B2(G469), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n279), .A2(KEYINPUT91), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT91), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n277), .A2(new_n301), .A3(new_n190), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n300), .A2(new_n259), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n190), .B1(new_n292), .B2(new_n277), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT92), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT92), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n306), .B(new_n190), .C1(new_n292), .C2(new_n277), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n303), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G469), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n308), .A2(new_n309), .A3(new_n283), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n298), .A2(new_n299), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G221), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT9), .B(G234), .Z(new_n313));
  AOI21_X1  g127(.A(new_n312), .B1(new_n313), .B2(new_n283), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT93), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n296), .A2(G469), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT90), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n296), .A2(new_n297), .A3(G469), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n291), .A2(new_n201), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n287), .B1(new_n319), .B2(new_n280), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n306), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n304), .A2(KEYINPUT92), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(G902), .B1(new_n323), .B2(new_n303), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n309), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n317), .A2(new_n318), .A3(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT93), .ZN(new_n327));
  INV_X1    g141(.A(new_n314), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n315), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G214), .B1(G237), .B2(G902), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n331), .B(KEYINPUT94), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT67), .B(G116), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G119), .ZN(new_n334));
  INV_X1    g148(.A(G116), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(G119), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT2), .B(G113), .Z(new_n337));
  XNOR2_X1  g151(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n275), .A3(new_n267), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n334), .B(new_n337), .C1(new_n335), .C2(G119), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT5), .ZN(new_n342));
  INV_X1    g156(.A(G119), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(G116), .ZN(new_n344));
  OAI211_X1 g158(.A(G113), .B(new_n344), .C1(new_n336), .C2(new_n342), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n262), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G110), .B(G122), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(KEYINPUT95), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n349), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n340), .A2(new_n351), .A3(new_n346), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(KEYINPUT6), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n347), .A2(new_n354), .A3(new_n349), .ZN(new_n355));
  INV_X1    g169(.A(G125), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n251), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n270), .A2(new_n272), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G125), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G224), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(G953), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n360), .B(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n353), .A2(new_n355), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT7), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n357), .A2(new_n359), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT97), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n262), .A2(KEYINPUT96), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n345), .A2(new_n341), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n369), .B(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(new_n349), .B(KEYINPUT8), .Z(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n360), .B1(new_n365), .B2(new_n362), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n368), .A2(new_n373), .A3(new_n374), .A4(new_n352), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n364), .A2(new_n283), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G210), .B1(G237), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n364), .A2(new_n375), .A3(new_n283), .A4(new_n377), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n332), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G953), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n382), .A2(G952), .ZN(new_n383));
  NAND2_X1  g197(.A1(G234), .A2(G237), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  XOR2_X1   g200(.A(KEYINPUT21), .B(G898), .Z(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(G902), .A3(G953), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n386), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n381), .A2(new_n392), .ZN(new_n393));
  OR2_X1    g207(.A1(KEYINPUT70), .A2(G237), .ZN(new_n394));
  NAND2_X1  g208(.A1(KEYINPUT70), .A2(G237), .ZN(new_n395));
  AOI21_X1  g209(.A(G953), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(G143), .B1(new_n396), .B2(G214), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n396), .A2(G143), .A3(G214), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n199), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT18), .ZN(new_n401));
  XNOR2_X1  g215(.A(G125), .B(G140), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n234), .B2(new_n235), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n403), .B(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(new_n227), .B2(new_n402), .ZN(new_n406));
  NAND2_X1  g220(.A1(KEYINPUT18), .A2(G131), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n398), .A2(new_n399), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n401), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n399), .ZN(new_n410));
  OAI21_X1  g224(.A(G131), .B1(new_n410), .B2(new_n397), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n398), .A2(new_n199), .A3(new_n399), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n402), .A2(KEYINPUT16), .ZN(new_n414));
  OR3_X1    g228(.A1(new_n356), .A2(KEYINPUT16), .A3(G140), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(G146), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT80), .ZN(new_n417));
  XOR2_X1   g231(.A(new_n402), .B(KEYINPUT19), .Z(new_n418));
  OR2_X1    g232(.A1(new_n418), .A2(new_n222), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n413), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n409), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G113), .B(G122), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(new_n202), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT98), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT17), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n426), .B1(new_n411), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n400), .A2(KEYINPUT98), .A3(KEYINPUT17), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n411), .A2(new_n412), .A3(new_n427), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n414), .A2(new_n415), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n227), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n416), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n428), .A2(new_n429), .A3(new_n430), .A4(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n423), .A3(new_n409), .ZN(new_n436));
  AOI21_X1  g250(.A(G475), .B1(new_n425), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n283), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n437), .B2(new_n283), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(KEYINPUT99), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT99), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n437), .A2(new_n442), .A3(new_n438), .A4(new_n283), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n435), .A2(new_n409), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(new_n423), .ZN(new_n445));
  INV_X1    g259(.A(new_n436), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n283), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n441), .A2(new_n443), .B1(G475), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n333), .A2(G122), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n335), .A2(G122), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n209), .A3(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(G128), .B(G143), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(new_n192), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n450), .B1(new_n449), .B2(KEYINPUT14), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n455), .A2(KEYINPUT100), .ZN(new_n456));
  OR2_X1    g270(.A1(new_n449), .A2(KEYINPUT14), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(KEYINPUT100), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n452), .B(new_n454), .C1(new_n459), .C2(new_n209), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n453), .A2(KEYINPUT13), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n223), .A2(G128), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n461), .B(G134), .C1(KEYINPUT13), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n453), .A2(new_n192), .ZN(new_n464));
  INV_X1    g278(.A(new_n452), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n209), .B1(new_n449), .B2(new_n451), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n463), .B(new_n464), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n313), .A2(G217), .A3(new_n382), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n469), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(KEYINPUT101), .A3(new_n283), .ZN(new_n474));
  INV_X1    g288(.A(G478), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(KEYINPUT15), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n476), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n473), .A2(KEYINPUT101), .A3(new_n283), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n448), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n393), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT25), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n249), .A2(G119), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n343), .A2(G128), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT77), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT77), .B1(new_n485), .B2(new_n486), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT24), .B(G110), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(KEYINPUT79), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n490), .B1(new_n487), .B2(new_n488), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT79), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT23), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n485), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n249), .A2(KEYINPUT23), .A3(G119), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n486), .A3(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n491), .B(new_n494), .C1(G110), .C2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n405), .A3(new_n417), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n498), .B(KEYINPUT78), .ZN(new_n501));
  INV_X1    g315(.A(G110), .ZN(new_n502));
  OAI221_X1 g316(.A(new_n433), .B1(new_n489), .B2(new_n490), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT83), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n382), .A2(G221), .A3(G234), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(G137), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT82), .B(KEYINPUT22), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT83), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n510), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n505), .A2(KEYINPUT83), .A3(new_n510), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n484), .B1(new_n515), .B2(new_n283), .ZN(new_n516));
  AOI211_X1 g330(.A(KEYINPUT25), .B(G902), .C1(new_n513), .C2(new_n514), .ZN(new_n517));
  INV_X1    g331(.A(G234), .ZN(new_n518));
  OAI21_X1  g332(.A(G217), .B1(new_n518), .B2(G902), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT76), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n516), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n283), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT84), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n515), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT85), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT85), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n515), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT26), .B(G101), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n396), .A2(G210), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n533), .B(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n270), .A2(new_n272), .A3(new_n201), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n195), .A2(G134), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n192), .A2(G137), .ZN(new_n540));
  OAI21_X1  g354(.A(G131), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n200), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT68), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(KEYINPUT68), .B1(new_n200), .B2(new_n541), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT69), .B1(new_n251), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n239), .A2(new_n230), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n542), .B(new_n543), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT69), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n538), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n338), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n548), .A2(new_n200), .A3(new_n541), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n270), .A2(new_n272), .A3(KEYINPUT66), .A4(new_n201), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT66), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n537), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n339), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI211_X1 g376(.A(new_n538), .B(new_n339), .C1(new_n548), .C2(new_n549), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(KEYINPUT28), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n536), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n538), .B(new_n339), .C1(new_n547), .C2(new_n551), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT30), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n554), .A2(new_n557), .A3(new_n568), .A4(new_n555), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n552), .B2(new_n568), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n570), .B2(new_n339), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n536), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT31), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(KEYINPUT31), .A3(new_n536), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n566), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT32), .ZN(new_n577));
  NOR2_X1   g391(.A1(G472), .A2(G902), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n251), .A2(new_n546), .A3(KEYINPUT69), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n550), .B1(new_n548), .B2(new_n549), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n537), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n339), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT74), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(new_n553), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n552), .A2(KEYINPUT74), .A3(new_n338), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(KEYINPUT28), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT29), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n535), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n588), .A2(new_n565), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n283), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT75), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n564), .B1(new_n560), .B2(new_n561), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n536), .ZN(new_n596));
  INV_X1    g410(.A(new_n571), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n535), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n598), .A3(new_n589), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n591), .A2(KEYINPUT75), .A3(new_n283), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n594), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n580), .B1(new_n601), .B2(G472), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n576), .A2(KEYINPUT73), .A3(new_n579), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT73), .ZN(new_n604));
  AND3_X1   g418(.A1(new_n571), .A2(KEYINPUT31), .A3(new_n536), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT31), .B1(new_n571), .B2(new_n536), .ZN(new_n606));
  OAI22_X1  g420(.A1(new_n605), .A2(new_n606), .B1(new_n536), .B2(new_n595), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n604), .B1(new_n607), .B2(new_n578), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n577), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n530), .B1(new_n602), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n330), .A2(new_n483), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  INV_X1    g426(.A(new_n332), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n603), .A2(new_n608), .ZN(new_n614));
  OAI21_X1  g428(.A(G472), .B1(new_n576), .B2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n315), .B2(new_n329), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n379), .A2(new_n380), .ZN(new_n618));
  AND4_X1   g432(.A1(new_n613), .A2(new_n617), .A3(new_n618), .A4(new_n529), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n473), .A2(new_n475), .A3(new_n283), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n475), .A2(new_n283), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n469), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n473), .B(new_n625), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n620), .B(new_n622), .C1(new_n626), .C2(new_n475), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(new_n448), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n391), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n619), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  NAND2_X1  g447(.A1(new_n447), .A2(G475), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n391), .B(KEYINPUT103), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n440), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n439), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n480), .A2(new_n634), .A3(new_n636), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT104), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n619), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G107), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT105), .B(KEYINPUT35), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  AND2_X1   g458(.A1(new_n614), .A2(new_n615), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n515), .A2(new_n283), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT25), .ZN(new_n647));
  INV_X1    g461(.A(new_n520), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n515), .A2(new_n484), .A3(new_n283), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n510), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n504), .B(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n523), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n656), .A2(new_n393), .A3(new_n482), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n316), .A2(KEYINPUT90), .B1(new_n309), .B2(new_n324), .ZN(new_n658));
  AOI211_X1 g472(.A(KEYINPUT93), .B(new_n314), .C1(new_n658), .C2(new_n318), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n327), .B1(new_n326), .B2(new_n328), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n645), .B(new_n657), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  NAND2_X1  g477(.A1(new_n602), .A2(new_n609), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n638), .A2(new_n634), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n385), .B(KEYINPUT107), .Z(new_n666));
  OAI21_X1  g480(.A(KEYINPUT106), .B1(new_n389), .B2(G900), .ZN(new_n667));
  OR3_X1    g481(.A1(new_n389), .A2(KEYINPUT106), .A3(G900), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n481), .A2(new_n665), .A3(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n381), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n656), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n330), .A2(new_n664), .A3(new_n671), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  INV_X1    g489(.A(new_n580), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n586), .A2(new_n535), .A3(new_n587), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n572), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n678), .B2(G902), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n609), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n448), .A2(new_n481), .A3(new_n332), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n618), .B(KEYINPUT38), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n680), .A2(new_n656), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT108), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT109), .B(KEYINPUT39), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n669), .B(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(KEYINPUT40), .B1(new_n330), .B2(new_n687), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n330), .A2(KEYINPUT40), .A3(new_n687), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  NOR2_X1   g505(.A1(new_n629), .A2(new_n670), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n330), .A2(new_n664), .A3(new_n673), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G146), .ZN(G48));
  NAND2_X1  g508(.A1(new_n308), .A2(new_n283), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G469), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n381), .A2(new_n696), .A3(new_n325), .A4(new_n328), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n664), .A2(new_n529), .A3(new_n630), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NAND4_X1  g515(.A1(new_n664), .A2(new_n529), .A3(new_n640), .A4(new_n698), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  NAND3_X1  g517(.A1(new_n696), .A2(new_n328), .A3(new_n325), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n664), .A2(new_n657), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G119), .ZN(G21));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n708), .B1(new_n521), .B2(new_n528), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n605), .A2(new_n606), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n536), .B1(new_n588), .B2(new_n565), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n578), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n515), .A2(new_n526), .A3(new_n523), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n526), .B1(new_n515), .B2(new_n523), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n650), .A2(new_n715), .A3(KEYINPUT110), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n709), .A2(new_n615), .A3(new_n712), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n448), .A2(new_n332), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n480), .A3(new_n618), .A4(new_n636), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n721), .A3(new_n705), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  AND2_X1   g537(.A1(new_n615), .A2(new_n712), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n724), .A2(new_n655), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n692), .A3(new_n698), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  NAND2_X1  g541(.A1(G469), .A2(G902), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n278), .A2(new_n281), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(G469), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n325), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n328), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n379), .A2(new_n613), .A3(new_n380), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n610), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n692), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(KEYINPUT42), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n577), .B1(new_n576), .B2(new_n579), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n602), .A2(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n709), .A2(new_n716), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n734), .A3(new_n692), .A4(new_n740), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n735), .A2(new_n737), .B1(new_n741), .B2(KEYINPUT42), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT111), .B(G131), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G33));
  NAND2_X1  g558(.A1(new_n735), .A2(new_n671), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n747));
  INV_X1    g561(.A(new_n448), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n747), .B1(new_n748), .B2(KEYINPUT112), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n627), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT113), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n645), .A2(new_n656), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n751), .A2(new_n756), .A3(new_n752), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n729), .A2(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n282), .A2(new_n295), .ZN(new_n762));
  OAI211_X1 g576(.A(G469), .B(new_n761), .C1(new_n762), .C2(KEYINPUT45), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT46), .B1(new_n763), .B2(new_n728), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n310), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(KEYINPUT46), .A3(new_n728), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n328), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n686), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n760), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n733), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n758), .B2(new_n759), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g587(.A(KEYINPUT114), .B(G137), .Z(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G39));
  AND3_X1   g589(.A1(new_n767), .A2(KEYINPUT47), .A3(new_n328), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT47), .B1(new_n767), .B2(new_n328), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n664), .A2(new_n529), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n736), .A2(new_n733), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(KEYINPUT115), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(KEYINPUT115), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  AOI21_X1  g599(.A(new_n666), .B1(new_n751), .B2(new_n752), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n786), .A2(new_n718), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n705), .A2(KEYINPUT119), .A3(new_n332), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT119), .B1(new_n705), .B2(new_n332), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n682), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n696), .A2(new_n325), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n328), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n771), .B(new_n787), .C1(new_n778), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n704), .A2(new_n733), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n786), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n725), .ZN(new_n799));
  INV_X1    g613(.A(new_n680), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n386), .A3(new_n529), .A4(new_n797), .ZN(new_n801));
  INV_X1    g615(.A(new_n627), .ZN(new_n802));
  OR3_X1    g616(.A1(new_n801), .A2(new_n748), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n793), .A2(new_n796), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n804), .A2(new_n805), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n787), .A2(new_n698), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n801), .A2(new_n629), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n383), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n739), .A2(new_n740), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n798), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n812), .B(new_n813), .C1(KEYINPUT48), .C2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n806), .A2(new_n807), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n719), .A2(new_n480), .A3(new_n618), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n732), .A2(new_n819), .A3(new_n670), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n656), .A3(new_n680), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n674), .A2(new_n693), .A3(new_n726), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT117), .ZN(new_n823));
  AOI22_X1  g637(.A1(new_n315), .A2(new_n329), .B1(new_n609), .B2(new_n602), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n824), .B(new_n673), .C1(new_n671), .C2(new_n692), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(new_n826), .A3(new_n726), .A4(new_n821), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n611), .A2(new_n661), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n699), .A2(new_n702), .A3(new_n706), .A4(new_n722), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n482), .B1(new_n802), .B2(new_n448), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n635), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n617), .A2(new_n381), .A3(new_n529), .A4(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n831), .A2(new_n832), .A3(new_n742), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n655), .A2(new_n669), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n665), .A2(new_n480), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n664), .B(new_n838), .C1(new_n659), .C2(new_n660), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n724), .A2(new_n328), .A3(new_n628), .A4(new_n731), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n733), .B(new_n837), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n745), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT116), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n839), .A2(new_n840), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n655), .A3(new_n669), .A4(new_n771), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n846), .A3(new_n745), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n836), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n823), .A2(KEYINPUT52), .A3(new_n827), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n830), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(KEYINPUT53), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n822), .A2(KEYINPUT52), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n830), .A2(new_n848), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n851), .A2(KEYINPUT54), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n816), .A2(KEYINPUT48), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n850), .A2(new_n852), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n717), .A2(new_n720), .A3(new_n704), .ZN(new_n859));
  AOI211_X1 g673(.A(new_n530), .B(new_n697), .C1(new_n602), .C2(new_n609), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n630), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(KEYINPUT118), .A3(new_n702), .A4(new_n706), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n699), .A2(new_n702), .A3(new_n706), .A4(new_n722), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT118), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n865), .A3(KEYINPUT53), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n843), .B2(new_n847), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n831), .A2(new_n742), .A3(new_n835), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n830), .A3(new_n853), .A4(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n857), .A2(new_n858), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n818), .A2(new_n855), .A3(new_n856), .A4(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(G952), .B2(G953), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n740), .A2(new_n613), .A3(new_n328), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n794), .B(KEYINPUT49), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n873), .A2(new_n874), .A3(new_n682), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n875), .A2(new_n800), .A3(new_n750), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n872), .A2(new_n876), .ZN(G75));
  AND3_X1   g691(.A1(new_n823), .A2(KEYINPUT52), .A3(new_n827), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT52), .B1(new_n823), .B2(new_n827), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT53), .B1(new_n880), .B2(new_n848), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n830), .A2(new_n867), .A3(new_n853), .A4(new_n868), .ZN(new_n882));
  OAI211_X1 g696(.A(G210), .B(G902), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n353), .A2(new_n355), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n363), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT121), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT55), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n883), .A2(new_n884), .A3(new_n885), .A4(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n382), .A2(G952), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n283), .B1(new_n857), .B2(new_n869), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT56), .B1(new_n894), .B2(G210), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n884), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n889), .B1(new_n895), .B2(new_n884), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(G51));
  XOR2_X1   g712(.A(new_n728), .B(KEYINPUT57), .Z(new_n899));
  INV_X1    g713(.A(new_n870), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n858), .B1(new_n857), .B2(new_n869), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n308), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n857), .A2(new_n869), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OR3_X1    g719(.A1(new_n905), .A2(new_n283), .A3(new_n763), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n891), .B1(new_n903), .B2(new_n906), .ZN(G54));
  NAND3_X1  g721(.A1(new_n894), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n436), .A3(new_n425), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n425), .A2(new_n436), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n894), .A2(KEYINPUT58), .A3(G475), .A4(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n909), .A2(new_n892), .A3(new_n911), .ZN(G60));
  INV_X1    g726(.A(new_n626), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n621), .B(KEYINPUT59), .ZN(new_n914));
  INV_X1    g728(.A(new_n901), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n913), .B(new_n914), .C1(new_n915), .C2(new_n870), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n855), .B2(new_n870), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n892), .B1(new_n917), .B2(new_n626), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n916), .A2(new_n918), .ZN(G63));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n920));
  NAND2_X1  g734(.A1(G217), .A2(G902), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT60), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n857), .B2(new_n869), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n653), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n892), .B1(new_n923), .B2(new_n515), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n923), .A2(new_n515), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n928), .A2(KEYINPUT61), .A3(new_n892), .A4(new_n924), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(G66));
  AND3_X1   g744(.A1(new_n831), .A2(new_n835), .A3(new_n832), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n382), .B1(new_n387), .B2(G224), .ZN(new_n934));
  AOI22_X1  g748(.A1(new_n932), .A2(new_n382), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n933), .B2(new_n934), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n886), .B1(G898), .B2(new_n382), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(G69));
  XNOR2_X1  g752(.A(new_n570), .B(new_n418), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n188), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n382), .B1(new_n940), .B2(G900), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n773), .B1(new_n782), .B2(new_n783), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n769), .A2(new_n618), .A3(new_n681), .A4(new_n815), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n943), .A2(new_n742), .A3(new_n745), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n674), .A2(new_n693), .A3(new_n726), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n825), .A2(KEYINPUT124), .A3(new_n726), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n942), .A2(new_n944), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n939), .B1(new_n950), .B2(new_n382), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n188), .A2(G953), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n941), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n690), .A2(new_n947), .A3(new_n948), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n690), .A2(new_n947), .A3(KEYINPUT62), .A4(new_n948), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n610), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n959), .A2(new_n833), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(new_n330), .A3(new_n687), .A4(new_n771), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n942), .A3(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n962), .A2(new_n382), .A3(new_n939), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n953), .A2(new_n963), .ZN(G72));
  XOR2_X1   g778(.A(new_n571), .B(KEYINPUT126), .Z(new_n965));
  NAND4_X1  g779(.A1(new_n942), .A2(new_n931), .A3(new_n944), .A4(new_n949), .ZN(new_n966));
  XOR2_X1   g780(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n967));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  AOI211_X1 g783(.A(new_n536), .B(new_n965), .C1(new_n966), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n598), .A2(new_n572), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n851), .A2(new_n854), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n892), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n958), .A2(new_n942), .A3(new_n931), .A4(new_n961), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n969), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(new_n536), .A3(new_n965), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n975), .A2(KEYINPUT127), .A3(new_n536), .A4(new_n965), .ZN(new_n979));
  AOI211_X1 g793(.A(new_n970), .B(new_n973), .C1(new_n978), .C2(new_n979), .ZN(G57));
endmodule


