//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(KEYINPUT16), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  OAI211_X1 g007(.A(new_n188), .B(G146), .C1(KEYINPUT16), .C2(new_n190), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G128), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n196), .A2(G128), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n197), .B(new_n199), .C1(new_n200), .C2(KEYINPUT23), .ZN(new_n201));
  XOR2_X1   g015(.A(KEYINPUT24), .B(G110), .Z(new_n202));
  XNOR2_X1  g016(.A(G119), .B(G128), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n201), .A2(G110), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n195), .A2(new_n204), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT74), .B(G110), .Z(new_n206));
  OAI22_X1  g020(.A1(new_n201), .A2(new_n206), .B1(new_n202), .B2(new_n203), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n187), .A2(new_n192), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n194), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G137), .ZN(new_n211));
  INV_X1    g025(.A(G953), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(G221), .A3(G234), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n211), .B(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n214), .B(KEYINPUT75), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n205), .A2(new_n209), .A3(new_n214), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G217), .ZN(new_n219));
  INV_X1    g033(.A(G902), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(G234), .B2(new_n220), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n218), .A2(G902), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n216), .A2(new_n220), .A3(new_n217), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n216), .A2(KEYINPUT25), .A3(new_n220), .A4(new_n217), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n222), .B1(new_n227), .B2(new_n221), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT32), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n231));
  INV_X1    g045(.A(G113), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT2), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT2), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G116), .B(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n231), .B1(new_n238), .B2(KEYINPUT67), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n240));
  AOI211_X1 g054(.A(new_n240), .B(KEYINPUT68), .C1(new_n236), .C2(new_n237), .ZN(new_n241));
  OAI22_X1  g055(.A1(new_n239), .A2(new_n241), .B1(new_n237), .B2(new_n236), .ZN(new_n242));
  XOR2_X1   g056(.A(G116), .B(G119), .Z(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT2), .B(G113), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT67), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT68), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n236), .A2(new_n237), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n238), .A2(KEYINPUT67), .A3(new_n231), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n242), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT30), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n253), .A2(new_n254), .A3(new_n255), .A4(G134), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  OAI22_X1  g071(.A1(new_n257), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n257), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT66), .B1(new_n255), .B2(G134), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n257), .A3(G137), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n255), .A2(G134), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G131), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT69), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n262), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n192), .A2(G143), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n198), .B1(new_n273), .B2(KEYINPUT1), .ZN(new_n274));
  INV_X1    g088(.A(G143), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G146), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n273), .B(new_n276), .C1(KEYINPUT1), .C2(new_n198), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n270), .A2(new_n272), .A3(new_n280), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n273), .A2(new_n276), .A3(KEYINPUT0), .A4(G128), .ZN(new_n282));
  XNOR2_X1  g096(.A(G143), .B(G146), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT0), .B(G128), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n260), .A2(KEYINPUT65), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n259), .A2(new_n288), .A3(new_n261), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n288), .B1(new_n259), .B2(new_n261), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n252), .B1(new_n281), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n280), .A2(new_n268), .A3(new_n262), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(new_n292), .A3(new_n252), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n251), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n250), .A2(new_n281), .A3(new_n292), .ZN(new_n298));
  NOR2_X1   g112(.A1(G237), .A2(G953), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G210), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n300), .B(KEYINPUT27), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G101), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n297), .A2(new_n298), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT31), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n250), .A2(new_n281), .A3(new_n292), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n259), .A2(new_n261), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n287), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n285), .B1(new_n309), .B2(new_n289), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n278), .A2(new_n279), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n311), .B1(new_n269), .B2(KEYINPUT69), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n310), .B1(new_n312), .B2(new_n272), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n295), .B1(new_n313), .B2(new_n252), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n307), .B1(new_n314), .B2(new_n251), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT31), .A3(new_n303), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n294), .A2(new_n292), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n249), .A3(new_n242), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n298), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT28), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT71), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n307), .B2(KEYINPUT28), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n298), .A2(KEYINPUT71), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n303), .B(KEYINPUT70), .Z(new_n326));
  AOI22_X1  g140(.A1(new_n306), .A2(new_n316), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(G472), .A2(G902), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n230), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT31), .B1(new_n315), .B2(new_n303), .ZN(new_n331));
  AND4_X1   g145(.A1(KEYINPUT31), .A2(new_n297), .A3(new_n298), .A4(new_n303), .ZN(new_n332));
  INV_X1    g146(.A(new_n324), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n323), .B1(new_n298), .B2(new_n318), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT71), .B1(new_n298), .B2(new_n323), .ZN(new_n335));
  NOR3_X1   g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n326), .ZN(new_n337));
  OAI22_X1  g151(.A1(new_n331), .A2(new_n332), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT32), .A3(new_n328), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n330), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n341));
  NOR4_X1   g155(.A1(new_n333), .A2(new_n334), .A3(new_n335), .A4(new_n326), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n315), .B2(new_n303), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n341), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n313), .A2(new_n250), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT28), .B1(new_n307), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n303), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(new_n343), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n347), .A2(new_n322), .A3(new_n324), .A4(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT73), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(G902), .B1(new_n350), .B2(new_n351), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n297), .A2(new_n298), .ZN(new_n354));
  AOI21_X1  g168(.A(KEYINPUT29), .B1(new_n354), .B2(new_n348), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n320), .A2(new_n322), .A3(new_n337), .A4(new_n324), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(KEYINPUT72), .A3(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n345), .A2(new_n352), .A3(new_n353), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G472), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n229), .B1(new_n340), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G221), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT9), .B(G234), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n362), .B(KEYINPUT76), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n361), .B1(new_n363), .B2(new_n220), .ZN(new_n364));
  XNOR2_X1  g178(.A(G110), .B(G140), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n212), .A2(G227), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n290), .A2(new_n291), .ZN(new_n368));
  INV_X1    g182(.A(G107), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(G104), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(G104), .ZN(new_n371));
  OR2_X1    g185(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G101), .ZN(new_n374));
  INV_X1    g188(.A(G104), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(G107), .ZN(new_n376));
  NAND2_X1  g190(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n373), .A2(new_n374), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(G101), .B1(new_n376), .B2(new_n370), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n381), .A2(new_n279), .A3(new_n278), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT10), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT10), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n280), .A2(new_n385), .A3(new_n381), .A4(new_n382), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n374), .B1(new_n373), .B2(new_n380), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT4), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n285), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT78), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n371), .B1(new_n372), .B2(new_n377), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n375), .A2(G107), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n376), .B2(new_n379), .ZN(new_n394));
  OAI21_X1  g208(.A(G101), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(KEYINPUT4), .A3(new_n381), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n390), .A2(new_n391), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n391), .B1(new_n390), .B2(new_n396), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n368), .B(new_n387), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT12), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n381), .A2(new_n382), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n311), .ZN(new_n403));
  AOI211_X1 g217(.A(new_n401), .B(new_n368), .C1(new_n383), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n383), .ZN(new_n405));
  INV_X1    g219(.A(new_n368), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT12), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n367), .B1(new_n400), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT79), .ZN(new_n410));
  INV_X1    g224(.A(new_n367), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n399), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n387), .B1(new_n397), .B2(new_n398), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n406), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n410), .B1(new_n399), .B2(new_n411), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n409), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT80), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT80), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n409), .B(new_n419), .C1(new_n415), .C2(new_n416), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(G469), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G469), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(new_n220), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n399), .A2(new_n411), .ZN(new_n424));
  OR2_X1    g238(.A1(new_n424), .A2(new_n408), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n395), .A2(KEYINPUT4), .A3(new_n381), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n389), .B(G101), .C1(new_n392), .C2(new_n394), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n286), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT78), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n390), .A2(new_n391), .A3(new_n396), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n368), .B1(new_n431), .B2(new_n387), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n367), .B1(new_n400), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(G902), .B1(new_n425), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n423), .B1(new_n434), .B2(new_n422), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n364), .B1(new_n421), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n363), .A2(G217), .A3(new_n212), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G116), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n439), .A2(KEYINPUT14), .A3(G122), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT14), .ZN(new_n441));
  XNOR2_X1  g255(.A(G116), .B(G122), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n369), .B(new_n440), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n369), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n275), .A2(G128), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n198), .A2(G143), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(new_n257), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n257), .B1(new_n445), .B2(new_n446), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n443), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n198), .A2(G143), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(KEYINPUT88), .A3(KEYINPUT13), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n275), .A2(KEYINPUT13), .A3(G128), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT86), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT13), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n459), .B(new_n460), .C1(new_n198), .C2(G143), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n446), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n445), .B2(new_n460), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n458), .B1(new_n464), .B2(KEYINPUT87), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n462), .B2(new_n463), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n257), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n444), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n442), .A2(new_n369), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n447), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(KEYINPUT89), .B(new_n452), .C1(new_n468), .C2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT89), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n460), .B1(new_n198), .B2(G143), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT86), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n475), .A2(KEYINPUT87), .A3(new_n446), .A4(new_n461), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n455), .B(KEYINPUT88), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n467), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n471), .B1(new_n478), .B2(G134), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n473), .B1(new_n479), .B2(new_n451), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n438), .B1(new_n472), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n476), .A2(new_n477), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n275), .A2(G128), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT13), .B1(new_n275), .B2(G128), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n484), .B2(new_n459), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT87), .B1(new_n485), .B2(new_n475), .ZN(new_n486));
  OAI21_X1  g300(.A(G134), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n471), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n452), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n437), .B1(new_n490), .B2(new_n473), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n220), .B1(new_n481), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(G478), .ZN(new_n493));
  OR2_X1    g307(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n494));
  NAND2_X1  g308(.A1(KEYINPUT90), .A2(KEYINPUT15), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR2_X1    g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n496), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G237), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n212), .A3(G214), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n275), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n299), .A2(G143), .A3(G214), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(KEYINPUT82), .A2(KEYINPUT18), .A3(G131), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n503), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n507), .A2(KEYINPUT82), .A3(KEYINPUT18), .A4(G131), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n187), .B(new_n192), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(G131), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n507), .A2(G131), .ZN(new_n513));
  NOR3_X1   g327(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT17), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n507), .A2(KEYINPUT17), .A3(G131), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n193), .A2(new_n194), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n510), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(G113), .B(G122), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(new_n375), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n510), .ZN(new_n522));
  INV_X1    g336(.A(new_n516), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n504), .A2(new_n260), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n511), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n522), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n519), .B(KEYINPUT84), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n521), .A2(KEYINPUT85), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n526), .A2(new_n193), .A3(new_n194), .A4(new_n515), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n519), .B1(new_n530), .B2(new_n510), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT85), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(G902), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G475), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT20), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n530), .A2(new_n510), .A3(new_n528), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT83), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n538), .A2(KEYINPUT19), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(KEYINPUT19), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n187), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n541), .B(new_n192), .C1(new_n187), .C2(new_n540), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n542), .B(new_n194), .C1(new_n512), .C2(new_n513), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n510), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n520), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(G475), .A2(G902), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n536), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n546), .A2(new_n536), .A3(new_n547), .ZN(new_n549));
  OAI22_X1  g363(.A1(new_n534), .A2(new_n535), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n499), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n436), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n242), .A2(new_n249), .A3(new_n396), .A4(new_n427), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT5), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n196), .A3(G116), .ZN(new_n555));
  OAI211_X1 g369(.A(G113), .B(new_n555), .C1(new_n243), .C2(new_n554), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n238), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n557), .A2(new_n402), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(G110), .B(G122), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT81), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n553), .A2(new_n561), .A3(new_n558), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT6), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n285), .A2(G125), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n280), .B2(G125), .ZN(new_n567));
  INV_X1    g381(.A(G224), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(G953), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n569), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n566), .B(new_n571), .C1(new_n280), .C2(G125), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT6), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n559), .A2(new_n574), .A3(new_n562), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n565), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n570), .A2(new_n572), .B1(new_n577), .B2(new_n571), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT8), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n561), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n557), .A2(new_n402), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n558), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n567), .A2(new_n577), .A3(new_n571), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n578), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(G902), .B1(new_n584), .B2(new_n564), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n576), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(G210), .B1(G237), .B2(G902), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n576), .A2(new_n585), .A3(new_n587), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G214), .B1(G237), .B2(G902), .ZN(new_n592));
  NAND2_X1  g406(.A1(G234), .A2(G237), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n593), .A2(G952), .A3(new_n212), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT21), .B(G898), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT91), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n593), .A2(G902), .A3(G953), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n595), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n591), .A2(new_n592), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n360), .A2(new_n552), .A3(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  OAI21_X1  g418(.A(G472), .B1(new_n327), .B2(G902), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n338), .A2(new_n328), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n607), .A2(new_n228), .A3(new_n436), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT92), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n490), .B1(new_n610), .B2(new_n438), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n489), .A2(KEYINPUT92), .A3(new_n437), .A4(new_n452), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n609), .B1(new_n481), .B2(new_n491), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n493), .A2(G902), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n492), .A2(new_n618), .A3(new_n493), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n492), .B2(new_n493), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n550), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n601), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n608), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT34), .B(G104), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G6));
  OAI21_X1  g440(.A(new_n537), .B1(new_n531), .B2(new_n532), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n521), .A2(KEYINPUT85), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n220), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n546), .A2(new_n547), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT20), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n546), .A2(new_n536), .A3(new_n547), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n629), .A2(G475), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n499), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n601), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n608), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT35), .B(G107), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT94), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n636), .B(new_n638), .ZN(G9));
  NAND2_X1  g453(.A1(new_n227), .A2(new_n221), .ZN(new_n640));
  OR3_X1    g454(.A1(new_n215), .A2(KEYINPUT95), .A3(KEYINPUT36), .ZN(new_n641));
  INV_X1    g455(.A(new_n210), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT95), .B1(new_n215), .B2(KEYINPUT36), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n642), .B1(new_n641), .B2(new_n643), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n221), .A2(G902), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n591), .A2(new_n592), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n551), .A2(new_n600), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n651), .A2(new_n436), .A3(new_n607), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  NAND2_X1  g469(.A1(new_n340), .A2(new_n359), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n595), .B1(new_n599), .B2(G900), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT96), .Z(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n499), .A2(new_n633), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n656), .A2(new_n661), .A3(new_n436), .A4(new_n651), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  OAI21_X1  g477(.A(new_n326), .B1(new_n307), .B2(new_n346), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n304), .A2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n665), .B2(G902), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n330), .A2(new_n339), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT97), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT97), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n330), .A2(new_n339), .A3(new_n669), .A4(new_n666), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n499), .A2(new_n550), .A3(new_n592), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n649), .ZN(new_n673));
  INV_X1    g487(.A(new_n590), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n587), .B1(new_n576), .B2(new_n585), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT38), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT38), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n591), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n673), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n671), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT40), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT98), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n421), .A2(new_n435), .ZN(new_n684));
  INV_X1    g498(.A(new_n364), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n658), .B(KEYINPUT39), .Z(new_n686));
  AND4_X1   g500(.A1(new_n683), .A2(new_n684), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n683), .B1(new_n436), .B2(new_n686), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n682), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT98), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n436), .A2(new_n683), .A3(new_n686), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n691), .A2(KEYINPUT40), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n681), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n275), .ZN(G45));
  AOI21_X1  g509(.A(new_n650), .B1(new_n340), .B2(new_n359), .ZN(new_n696));
  AOI21_X1  g510(.A(KEYINPUT89), .B1(new_n489), .B2(new_n452), .ZN(new_n697));
  NOR3_X1   g511(.A1(new_n479), .A2(new_n473), .A3(new_n451), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n437), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n480), .A2(new_n438), .ZN(new_n700));
  AOI21_X1  g514(.A(G902), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(KEYINPUT93), .B1(new_n701), .B2(G478), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n492), .A2(new_n618), .A3(new_n493), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n633), .B1(new_n704), .B2(new_n617), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT99), .B1(new_n705), .B2(new_n659), .ZN(new_n706));
  AND4_X1   g520(.A1(KEYINPUT99), .A2(new_n621), .A3(new_n550), .A4(new_n659), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n696), .A2(new_n708), .A3(new_n436), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  NAND2_X1  g524(.A1(new_n434), .A2(new_n422), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n411), .B1(new_n414), .B2(new_n399), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n424), .A2(new_n408), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n220), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(G469), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n711), .A2(new_n685), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n360), .A2(new_n623), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND3_X1  g534(.A1(new_n360), .A2(new_n635), .A3(new_n717), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  NAND3_X1  g536(.A1(new_n696), .A2(new_n652), .A3(new_n717), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NOR2_X1   g538(.A1(new_n676), .A2(new_n672), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n725), .A2(new_n600), .A3(new_n717), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n347), .A2(new_n322), .A3(new_n324), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n306), .A2(new_n316), .B1(new_n727), .B2(new_n326), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n728), .A2(new_n329), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n228), .A3(new_n605), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n730), .A2(KEYINPUT100), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(KEYINPUT100), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n726), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  INV_X1    g548(.A(new_n707), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n729), .A2(new_n605), .A3(new_n649), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n591), .A2(new_n592), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n716), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT99), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n622), .B2(new_n658), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n735), .A2(new_n736), .A3(new_n738), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n339), .B(new_n743), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n358), .A2(G472), .B1(new_n230), .B2(new_n606), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n229), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n589), .A2(new_n592), .A3(new_n590), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT101), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n417), .A2(new_n422), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n364), .B1(new_n435), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n589), .A2(KEYINPUT101), .A3(new_n592), .A4(new_n590), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n749), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n746), .A2(KEYINPUT42), .A3(new_n708), .A4(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n360), .A2(new_n753), .A3(new_n708), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT103), .ZN(new_n756));
  XNOR2_X1  g570(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n756), .B1(new_n755), .B2(new_n758), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n754), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  AND2_X1   g576(.A1(new_n360), .A2(new_n753), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n661), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n550), .B1(new_n704), .B2(new_n617), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n767), .B1(new_n768), .B2(KEYINPUT43), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n621), .A2(new_n633), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(KEYINPUT105), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n621), .A2(KEYINPUT43), .A3(new_n633), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT106), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT106), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n621), .A2(new_n776), .A3(KEYINPUT43), .A4(new_n633), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT107), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n773), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n649), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n607), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n779), .B1(new_n773), .B2(new_n778), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n766), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n773), .A2(new_n778), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT107), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(KEYINPUT44), .A3(new_n780), .A4(new_n782), .ZN(new_n788));
  INV_X1    g602(.A(new_n423), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT45), .B1(new_n418), .B2(new_n420), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT45), .ZN(new_n791));
  OAI21_X1  g605(.A(G469), .B1(new_n417), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n789), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT46), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  OAI211_X1 g609(.A(KEYINPUT46), .B(new_n789), .C1(new_n790), .C2(new_n792), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n711), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n749), .A2(new_n752), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AND4_X1   g613(.A1(new_n685), .A2(new_n797), .A3(new_n686), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n785), .A2(new_n788), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G137), .ZN(G39));
  INV_X1    g616(.A(new_n656), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(new_n708), .A3(new_n229), .A4(new_n799), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n797), .A2(KEYINPUT47), .A3(new_n685), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT47), .B1(new_n797), .B2(new_n685), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G140), .ZN(G42));
  AOI21_X1  g623(.A(new_n595), .B1(new_n773), .B2(new_n778), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n798), .A2(new_n716), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n746), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT48), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n229), .A2(new_n595), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n811), .A2(new_n668), .A3(new_n670), .A4(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n622), .ZN(new_n816));
  INV_X1    g630(.A(G952), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n816), .A2(new_n817), .A3(G953), .ZN(new_n818));
  INV_X1    g632(.A(new_n738), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n731), .A2(new_n732), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n810), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n813), .B(new_n818), .C1(new_n819), .C2(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n810), .A2(new_n736), .A3(new_n811), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n815), .A2(new_n550), .A3(new_n621), .ZN(new_n824));
  OR2_X1    g638(.A1(new_n716), .A2(new_n592), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n825), .A2(new_n826), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n677), .A2(new_n679), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n820), .A3(new_n810), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n823), .B(new_n824), .C1(KEYINPUT50), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n806), .A2(new_n807), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n711), .A2(new_n715), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n833), .B1(new_n685), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT50), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n835), .A2(new_n799), .B1(new_n836), .B2(new_n830), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n832), .B1(new_n837), .B2(new_n821), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT51), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT51), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n840), .B(new_n832), .C1(new_n837), .C2(new_n821), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n822), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n622), .A2(KEYINPUT108), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT108), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n705), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT109), .B1(new_n847), .B2(new_n601), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT109), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n602), .A2(new_n849), .A3(new_n844), .A4(new_n846), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n608), .A3(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(new_n603), .A3(new_n636), .A4(new_n653), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n733), .A2(new_n723), .A3(new_n718), .A4(new_n721), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI211_X1 g668(.A(new_n781), .B(new_n658), .C1(new_n340), .C2(new_n359), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n552), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n736), .A2(new_n751), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n708), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n859), .A2(new_n799), .B1(new_n661), .B2(new_n763), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n854), .A2(new_n761), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n649), .A2(new_n658), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT110), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n667), .A3(new_n725), .A4(new_n751), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n709), .A2(new_n865), .A3(new_n662), .A4(new_n741), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT52), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n843), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n855), .A2(new_n552), .B1(new_n857), .B2(new_n708), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n764), .B1(new_n869), .B2(new_n798), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n755), .A2(new_n758), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT103), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n870), .B1(new_n874), .B2(new_n754), .ZN(new_n875));
  XNOR2_X1  g689(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n866), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(KEYINPUT52), .B2(new_n866), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT115), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n853), .B(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n852), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n875), .A2(new_n880), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n868), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(KEYINPUT54), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n883), .B1(new_n861), .B2(new_n879), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT112), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT112), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n891), .B(new_n883), .C1(new_n861), .C2(new_n879), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n866), .A2(KEYINPUT52), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n866), .A2(KEYINPUT52), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n843), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n875), .A2(new_n854), .A3(new_n895), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT114), .ZN(new_n898));
  INV_X1    g712(.A(new_n861), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT114), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(new_n900), .A3(new_n895), .A4(new_n896), .ZN(new_n901));
  AOI22_X1  g715(.A1(new_n890), .A2(new_n892), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n842), .B(new_n888), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n817), .A2(new_n212), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n228), .A2(new_n685), .A3(new_n592), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n834), .B2(KEYINPUT49), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(KEYINPUT49), .B2(new_n834), .ZN(new_n909));
  OR4_X1    g723(.A1(new_n671), .A2(new_n909), .A3(new_n829), .A4(new_n770), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n906), .A2(new_n910), .ZN(G75));
  AOI21_X1  g725(.A(new_n220), .B1(new_n868), .B2(new_n885), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n913), .A3(G210), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT56), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n565), .A2(new_n575), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n573), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT55), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n914), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n913), .B1(new_n912), .B2(G210), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n212), .A2(G952), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT56), .B1(new_n912), .B2(G210), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n918), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n921), .A2(new_n925), .ZN(G51));
  AOI21_X1  g740(.A(new_n903), .B1(new_n868), .B2(new_n885), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n887), .A2(new_n927), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n423), .B(KEYINPUT57), .Z(new_n929));
  OAI22_X1  g743(.A1(new_n928), .A2(new_n929), .B1(new_n712), .B2(new_n713), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n886), .A2(G902), .ZN(new_n931));
  OR3_X1    g745(.A1(new_n931), .A2(new_n790), .A3(new_n792), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n922), .B1(new_n930), .B2(new_n932), .ZN(G54));
  AND3_X1   g747(.A1(new_n912), .A2(KEYINPUT58), .A3(G475), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n923), .B1(new_n934), .B2(new_n546), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n546), .B2(new_n934), .ZN(G60));
  NAND2_X1  g750(.A1(new_n699), .A2(new_n700), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n613), .B1(new_n937), .B2(new_n609), .ZN(new_n938));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n923), .B1(new_n928), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n890), .A2(new_n892), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n898), .A2(new_n901), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n903), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n941), .B1(new_n946), .B2(new_n887), .ZN(new_n947));
  INV_X1    g761(.A(new_n938), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(G63));
  INV_X1    g763(.A(new_n886), .ZN(new_n950));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT60), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n218), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n868), .B2(new_n885), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n922), .B1(new_n954), .B2(new_n646), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT118), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n954), .B2(new_n646), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n958), .A2(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n953), .B(new_n955), .C1(new_n958), .C2(KEYINPUT61), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(G66));
  INV_X1    g776(.A(new_n597), .ZN(new_n963));
  OAI21_X1  g777(.A(G953), .B1(new_n963), .B2(new_n568), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n854), .B2(G953), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n916), .B1(G898), .B2(new_n212), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G69));
  AOI21_X1  g781(.A(new_n212), .B1(G227), .B2(G900), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT121), .Z(new_n969));
  OAI21_X1  g783(.A(new_n541), .B1(new_n187), .B2(new_n540), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n314), .B(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n212), .A2(G900), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT122), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n709), .A2(new_n662), .A3(new_n741), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n801), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n797), .A2(new_n685), .A3(new_n686), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n746), .A2(new_n725), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT123), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n725), .ZN(new_n981));
  AOI211_X1 g795(.A(new_n229), .B(new_n981), .C1(new_n744), .C2(new_n745), .ZN(new_n982));
  AOI22_X1  g796(.A1(new_n793), .A2(new_n794), .B1(new_n422), .B2(new_n434), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n364), .B1(new_n983), .B2(new_n796), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT123), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n982), .A2(new_n984), .A3(new_n985), .A4(new_n686), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n980), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n761), .A2(new_n987), .A3(new_n808), .A4(new_n764), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n975), .B1(new_n801), .B2(new_n976), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n977), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n974), .B1(new_n990), .B2(G953), .ZN(new_n991));
  INV_X1    g805(.A(new_n681), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n687), .A2(new_n688), .A3(new_n682), .ZN(new_n993));
  AOI21_X1  g807(.A(KEYINPUT40), .B1(new_n691), .B2(new_n692), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT62), .B1(new_n995), .B2(new_n976), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n709), .A2(new_n662), .A3(new_n741), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT62), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n694), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n808), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n687), .A2(new_n688), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n847), .A2(new_n634), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1001), .A2(new_n360), .A3(new_n799), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n801), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT119), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n801), .A2(new_n1003), .A3(KEYINPUT119), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1000), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n971), .B1(new_n1008), .B2(G953), .ZN(new_n1009));
  INV_X1    g823(.A(KEYINPUT120), .ZN(new_n1010));
  AOI22_X1  g824(.A1(new_n972), .A2(new_n991), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(KEYINPUT120), .B(new_n971), .C1(new_n1008), .C2(G953), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n969), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n977), .A2(new_n988), .ZN(new_n1014));
  INV_X1    g828(.A(new_n989), .ZN(new_n1015));
  AOI21_X1  g829(.A(G953), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n972), .B1(new_n1016), .B2(new_n973), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1018));
  AND4_X1   g832(.A1(new_n969), .A2(new_n1017), .A3(new_n1018), .A4(new_n1012), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1013), .A2(new_n1019), .ZN(G72));
  NAND2_X1  g834(.A1(new_n354), .A2(new_n303), .ZN(new_n1021));
  INV_X1    g835(.A(new_n808), .ZN(new_n1022));
  INV_X1    g836(.A(new_n999), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n998), .B1(new_n694), .B2(new_n997), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1007), .ZN(new_n1026));
  AOI21_X1  g840(.A(KEYINPUT119), .B1(new_n801), .B2(new_n1003), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n1025), .B(new_n854), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(G472), .A2(G902), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT63), .Z(new_n1030));
  AOI21_X1  g844(.A(new_n1021), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT124), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1031), .B(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(new_n988), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n801), .A2(new_n975), .A3(new_n976), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1034), .A2(new_n1015), .A3(new_n854), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(KEYINPUT125), .ZN(new_n1037));
  AND3_X1   g851(.A1(new_n1036), .A2(new_n1037), .A3(new_n1030), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1037), .B1(new_n1036), .B2(new_n1030), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n354), .A2(new_n303), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1040), .ZN(new_n1041));
  NOR3_X1   g855(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n1041), .A2(new_n1021), .A3(new_n1030), .ZN(new_n1043));
  XOR2_X1   g857(.A(new_n1043), .B(KEYINPUT126), .Z(new_n1044));
  OAI21_X1  g858(.A(new_n923), .B1(new_n902), .B2(new_n1044), .ZN(new_n1045));
  NOR3_X1   g859(.A1(new_n1033), .A2(new_n1042), .A3(new_n1045), .ZN(G57));
endmodule


