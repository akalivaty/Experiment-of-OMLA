//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1339,
    new_n1340, new_n1341, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1424, new_n1425,
    new_n1426, new_n1427;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT66), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n209), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n214), .A2(new_n225), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(new_n217), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n202), .A2(G68), .ZN(new_n244));
  INV_X1    g0044(.A(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n243), .B(new_n249), .ZN(G351));
  NAND2_X1  g0050(.A1(new_n208), .A2(G274), .ZN(new_n251));
  XOR2_X1   g0051(.A(KEYINPUT67), .B(G45), .Z(new_n252));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT68), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n256), .A2(new_n260), .A3(new_n257), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n254), .B1(new_n262), .B2(G244), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT69), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  OAI211_X1 g0067(.A(G232), .B(new_n265), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(G238), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(G107), .A3(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n268), .A2(new_n269), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n256), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n263), .A2(new_n264), .A3(new_n277), .ZN(new_n278));
  AND3_X1   g0078(.A1(new_n256), .A2(new_n260), .A3(new_n257), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n260), .B1(new_n256), .B2(new_n257), .ZN(new_n280));
  OAI21_X1  g0080(.A(G244), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT67), .B(G45), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n208), .B(G274), .C1(new_n282), .C2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n277), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT69), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n278), .A2(new_n285), .A3(G200), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n228), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(KEYINPUT8), .B(G58), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n291), .A2(new_n292), .B1(G20), .B2(G77), .ZN(new_n293));
  XOR2_X1   g0093(.A(KEYINPUT15), .B(G87), .Z(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(new_n209), .A3(G33), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n289), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(new_n288), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n208), .A2(G20), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G77), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(G77), .B2(new_n297), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n286), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT70), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n278), .A2(new_n285), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(G190), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  AOI211_X1 g0108(.A(KEYINPUT70), .B(new_n308), .C1(new_n278), .C2(new_n285), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n304), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n202), .B1(new_n208), .B2(G20), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n299), .A2(new_n311), .B1(new_n202), .B2(new_n298), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n209), .A2(G33), .ZN(new_n313));
  INV_X1    g0113(.A(G150), .ZN(new_n314));
  INV_X1    g0114(.A(new_n292), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n290), .A2(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(G20), .B2(new_n203), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n312), .B1(new_n317), .B2(new_n289), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(KEYINPUT9), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(KEYINPUT9), .ZN(new_n321));
  NAND2_X1  g0121(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT71), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT10), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n254), .B1(new_n262), .B2(G226), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n272), .A2(new_n273), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(G222), .A3(new_n265), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(G223), .A3(G1698), .ZN(new_n330));
  INV_X1    g0130(.A(G77), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n329), .B(new_n330), .C1(new_n331), .C2(new_n328), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n276), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G200), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n327), .A2(new_n333), .A3(G190), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n323), .A2(new_n326), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n335), .A2(new_n336), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n324), .B(new_n325), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n306), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n303), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n278), .A2(new_n285), .A3(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n319), .B1(new_n334), .B2(new_n345), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G179), .B2(new_n334), .ZN(new_n349));
  AND4_X1   g0149(.A1(new_n310), .A2(new_n341), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT78), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT74), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n272), .A2(new_n209), .A3(new_n273), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n272), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n273), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n245), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n216), .A2(new_n245), .ZN(new_n358));
  OAI21_X1  g0158(.A(G20), .B1(new_n358), .B2(new_n201), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n292), .A2(G159), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(KEYINPUT16), .A3(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n352), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n266), .A2(new_n267), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n363), .B2(new_n209), .ZN(new_n364));
  INV_X1    g0164(.A(new_n356), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n359), .A2(KEYINPUT16), .A3(new_n360), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(KEYINPUT74), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n289), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n359), .A2(new_n360), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT76), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n372), .B1(new_n357), .B2(new_n373), .ZN(new_n374));
  AOI211_X1 g0174(.A(KEYINPUT76), .B(new_n245), .C1(new_n355), .C2(new_n356), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n370), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n369), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n299), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n291), .A2(new_n300), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n378), .A2(new_n379), .B1(new_n297), .B2(new_n291), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G200), .ZN(new_n382));
  OR2_X1    g0182(.A1(G223), .A2(G1698), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(G226), .B2(new_n265), .ZN(new_n384));
  INV_X1    g0184(.A(G87), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n384), .A2(new_n363), .B1(new_n271), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n276), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n283), .B1(new_n217), .B2(new_n258), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n382), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n258), .A2(new_n217), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT77), .B1(new_n254), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT77), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n283), .B(new_n393), .C1(new_n217), .C2(new_n258), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n392), .A2(new_n394), .A3(new_n308), .A4(new_n387), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  AND4_X1   g0196(.A1(KEYINPUT17), .A2(new_n377), .A3(new_n381), .A4(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n380), .B1(new_n369), .B2(new_n376), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT17), .B1(new_n398), .B2(new_n396), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n351), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT18), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT74), .B1(new_n366), .B2(new_n367), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n357), .A2(new_n352), .A3(new_n361), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n288), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n370), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n371), .B1(new_n366), .B2(KEYINPUT76), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n357), .A2(new_n373), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n381), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n345), .B1(new_n388), .B2(new_n389), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n392), .A2(new_n394), .A3(new_n342), .A4(new_n387), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n401), .B1(new_n409), .B2(new_n413), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n398), .A2(KEYINPUT18), .A3(new_n412), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n377), .A2(new_n381), .A3(new_n396), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n398), .A2(KEYINPUT17), .A3(new_n396), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(KEYINPUT78), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n400), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n298), .A2(new_n245), .ZN(new_n424));
  XNOR2_X1  g0224(.A(new_n424), .B(KEYINPUT12), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n292), .A2(G50), .B1(G20), .B2(new_n245), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n331), .B2(new_n313), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n427), .A2(KEYINPUT11), .A3(new_n288), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n299), .A2(G68), .A3(new_n300), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n425), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT11), .B1(new_n427), .B2(new_n288), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT73), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT14), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G97), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT72), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(KEYINPUT72), .A2(G33), .A3(G97), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n217), .A2(G1698), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(G226), .B2(G1698), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n437), .B(new_n438), .C1(new_n440), .C2(new_n363), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n254), .B1(new_n441), .B2(new_n276), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT13), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n262), .A2(G238), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n443), .B1(new_n442), .B2(new_n444), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n434), .B(G169), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n441), .A2(new_n276), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n283), .ZN(new_n449));
  INV_X1    g0249(.A(G238), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(new_n259), .B2(new_n261), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT13), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n442), .A2(new_n444), .A3(new_n443), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(G179), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n447), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n453), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n434), .B1(new_n456), .B2(G169), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n433), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(G169), .B1(new_n445), .B2(new_n446), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT14), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n460), .A2(KEYINPUT73), .A3(new_n454), .A4(new_n447), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n432), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n456), .A2(G200), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n452), .A2(G190), .A3(new_n453), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n432), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n350), .A2(new_n423), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G244), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n272), .B2(new_n273), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT4), .B1(new_n470), .B2(new_n265), .ZN(new_n471));
  AOI21_X1  g0271(.A(KEYINPUT82), .B1(G33), .B2(G283), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(KEYINPUT82), .A2(G33), .A3(G283), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G250), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT83), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT4), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n480), .A2(G1698), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n481), .B(G244), .C1(new_n267), .C2(new_n266), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT81), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n328), .A2(KEYINPUT81), .A3(G244), .A4(new_n481), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n478), .A2(new_n479), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(G244), .B(new_n265), .C1(new_n266), .C2(new_n267), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n480), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n475), .A3(new_n476), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n484), .A2(new_n485), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT83), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n486), .A2(new_n491), .A3(new_n276), .ZN(new_n492));
  OR2_X1    g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G45), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(G1), .ZN(new_n497));
  INV_X1    g0297(.A(new_n228), .ZN(new_n498));
  AOI22_X1  g0298(.A1(new_n495), .A2(new_n497), .B1(new_n498), .B2(new_n255), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n208), .A2(G45), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n493), .B2(new_n494), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n499), .A2(G257), .B1(G274), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n492), .A2(G190), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT84), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n492), .A2(new_n502), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G200), .ZN(new_n506));
  INV_X1    g0306(.A(new_n502), .ZN(new_n507));
  AND2_X1   g0307(.A1(new_n475), .A2(new_n476), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n508), .A2(new_n488), .A3(new_n484), .A4(new_n485), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n256), .B1(new_n509), .B2(KEYINPUT83), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n510), .B2(new_n486), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT84), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n512), .A3(G190), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n297), .A2(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n208), .A2(G33), .ZN(new_n515));
  AND4_X1   g0315(.A1(new_n228), .A2(new_n297), .A3(new_n287), .A4(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(G97), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  OR3_X1    g0318(.A1(new_n315), .A2(KEYINPUT79), .A3(new_n331), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT79), .B1(new_n315), .B2(new_n331), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT6), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n521), .A2(new_n218), .A3(G107), .ZN(new_n522));
  XNOR2_X1  g0322(.A(G97), .B(G107), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n519), .B(new_n520), .C1(new_n524), .C2(new_n209), .ZN(new_n525));
  INV_X1    g0325(.A(G107), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n355), .B2(new_n356), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n288), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(KEYINPUT80), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT80), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n530), .B(new_n288), .C1(new_n525), .C2(new_n527), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n518), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n504), .A2(new_n506), .A3(new_n513), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n511), .A2(new_n342), .ZN(new_n534));
  OAI21_X1  g0334(.A(G107), .B1(new_n364), .B2(new_n365), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n523), .A2(new_n521), .ZN(new_n536));
  INV_X1    g0336(.A(new_n522), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G20), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n535), .A2(new_n539), .A3(new_n519), .A4(new_n520), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n530), .B1(new_n540), .B2(new_n288), .ZN(new_n541));
  INV_X1    g0341(.A(new_n531), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n517), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n534), .B(new_n543), .C1(G169), .C2(new_n511), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n497), .A2(G274), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT85), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n497), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n500), .A2(KEYINPUT85), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n256), .A2(G250), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n545), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n450), .A2(G1698), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n266), .B2(new_n267), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT86), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G116), .ZN(new_n556));
  OAI211_X1 g0356(.A(G244), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n552), .B(KEYINPUT86), .C1(new_n267), .C2(new_n266), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n555), .A2(new_n556), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n551), .B1(new_n559), .B2(new_n276), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n560), .A2(G169), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n342), .ZN(new_n562));
  NOR3_X1   g0362(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n563), .A2(KEYINPUT87), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n563), .A2(KEYINPUT87), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n437), .B2(new_n438), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n564), .A2(new_n565), .B1(new_n567), .B2(G20), .ZN(new_n568));
  AOI21_X1  g0368(.A(G20), .B1(new_n272), .B2(new_n273), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n209), .A2(G33), .A3(G97), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n569), .A2(G68), .B1(new_n570), .B2(new_n566), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n289), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n294), .A2(new_n297), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n516), .ZN(new_n575));
  INV_X1    g0375(.A(new_n294), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n561), .B(new_n562), .C1(new_n574), .C2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n575), .A2(new_n385), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n572), .A2(new_n573), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n560), .A2(G190), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(new_n382), .C2(new_n560), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n533), .A2(new_n544), .A3(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(G264), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n585));
  OAI211_X1 g0385(.A(G257), .B(new_n265), .C1(new_n266), .C2(new_n267), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n272), .A2(G303), .A3(new_n273), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT88), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT88), .A4(new_n587), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n276), .ZN(new_n593));
  INV_X1    g0393(.A(new_n494), .ZN(new_n594));
  NOR2_X1   g0394(.A1(KEYINPUT5), .A2(G41), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n497), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(G270), .A3(new_n256), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n501), .A2(G274), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(G190), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n297), .A2(G116), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n516), .B2(G116), .ZN(new_n603));
  AOI21_X1  g0403(.A(G20), .B1(new_n271), .B2(G97), .ZN(new_n604));
  AND3_X1   g0404(.A1(KEYINPUT82), .A2(G33), .A3(G283), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n604), .B1(new_n605), .B2(new_n472), .ZN(new_n606));
  INV_X1    g0406(.A(G116), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n287), .A2(new_n228), .B1(G20), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(KEYINPUT20), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT20), .B1(new_n606), .B2(new_n608), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n603), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n256), .B1(new_n590), .B2(new_n591), .ZN(new_n614));
  OAI21_X1  g0414(.A(G200), .B1(new_n614), .B2(new_n599), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n601), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT23), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n209), .B2(G107), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n526), .A2(KEYINPUT23), .A3(G20), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n209), .B(G87), .C1(new_n266), .C2(new_n267), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT22), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT22), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n328), .A2(new_n625), .A3(new_n209), .A4(G87), .ZN(new_n626));
  AOI211_X1 g0426(.A(KEYINPUT24), .B(new_n622), .C1(new_n624), .C2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT24), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n624), .A2(new_n626), .ZN(new_n629));
  INV_X1    g0429(.A(new_n622), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n288), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n575), .A2(new_n526), .ZN(new_n633));
  XOR2_X1   g0433(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n634));
  NOR2_X1   g0434(.A1(new_n297), .A2(G107), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT90), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(G294), .ZN(new_n640));
  INV_X1    g0440(.A(G294), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(KEYINPUT90), .ZN(new_n642));
  OAI21_X1  g0442(.A(G33), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(G257), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n644));
  OAI211_X1 g0444(.A(G250), .B(new_n265), .C1(new_n266), .C2(new_n267), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n276), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n499), .A2(G264), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n308), .A2(new_n647), .A3(new_n598), .A4(new_n648), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n646), .A2(new_n276), .B1(new_n499), .B2(G264), .ZN(new_n650));
  AOI21_X1  g0450(.A(G200), .B1(new_n650), .B2(new_n598), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT91), .B1(new_n638), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n650), .A2(new_n308), .A3(new_n598), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n647), .A2(new_n598), .A3(new_n648), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n654), .B1(new_n655), .B2(G200), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT91), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(new_n632), .A4(new_n637), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n616), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n599), .B1(new_n592), .B2(new_n276), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n612), .A2(G169), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT21), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n606), .A2(new_n608), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT20), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n609), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n345), .B1(new_n666), .B2(new_n603), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT21), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n667), .B(new_n668), .C1(new_n599), .C2(new_n614), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n599), .A2(new_n342), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n593), .A2(new_n612), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n650), .A2(new_n598), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n345), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n655), .A2(new_n342), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n625), .B1(new_n569), .B2(G87), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n623), .A2(KEYINPUT22), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n630), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT24), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n629), .A2(new_n628), .A3(new_n630), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n289), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n637), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n674), .B(new_n675), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n670), .A2(new_n672), .A3(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n659), .A2(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n468), .A2(new_n584), .A3(new_n685), .ZN(G372));
  NAND3_X1  g0486(.A1(new_n533), .A2(new_n544), .A3(new_n583), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n653), .A2(new_n658), .ZN(new_n688));
  INV_X1    g0488(.A(new_n683), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n670), .A2(new_n672), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n687), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT26), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n578), .A2(new_n582), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n544), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n544), .A2(new_n693), .A3(new_n694), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n578), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n468), .B1(new_n692), .B2(new_n698), .ZN(new_n699));
  AND3_X1   g0499(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n462), .B1(new_n465), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n400), .A2(new_n421), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n416), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n341), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n704), .A2(new_n349), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n699), .A2(new_n705), .ZN(G369));
  NAND3_X1  g0506(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT27), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT27), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G213), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(G343), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n613), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n690), .B(new_n714), .Z(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n616), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n653), .A2(new_n658), .B1(new_n638), .B2(new_n712), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(new_n689), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n689), .A2(new_n713), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n718), .A2(new_n690), .A3(new_n683), .A4(new_n713), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n724), .A2(new_n720), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT92), .ZN(G399));
  INV_X1    g0527(.A(new_n212), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G41), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n564), .A2(new_n565), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G116), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(new_n732), .A3(G1), .ZN(new_n733));
  INV_X1    g0533(.A(new_n227), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n733), .B1(new_n734), .B2(new_n730), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT95), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n697), .B1(new_n737), .B2(new_n695), .ZN(new_n738));
  NOR4_X1   g0538(.A1(new_n544), .A2(new_n694), .A3(KEYINPUT95), .A4(new_n693), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n578), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT96), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n692), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(KEYINPUT96), .B1(new_n687), .B2(new_n691), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(KEYINPUT29), .B(new_n713), .C1(new_n740), .C2(new_n744), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n687), .A2(new_n691), .ZN(new_n746));
  INV_X1    g0546(.A(new_n578), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n532), .B1(new_n345), .B2(new_n505), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n583), .A2(new_n748), .A3(KEYINPUT26), .A4(new_n534), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n747), .B1(new_n749), .B2(new_n695), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n712), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT29), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n745), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT94), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT30), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n593), .A2(new_n560), .A3(new_n671), .A4(new_n650), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n755), .B1(new_n505), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n560), .A2(new_n671), .A3(new_n650), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n614), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(new_n511), .A3(KEYINPUT30), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n559), .A2(new_n276), .ZN(new_n762));
  INV_X1    g0562(.A(new_n551), .ZN(new_n763));
  AOI21_X1  g0563(.A(G179), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n764), .B(new_n673), .C1(new_n599), .C2(new_n614), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n511), .ZN(new_n766));
  OAI211_X1 g0566(.A(KEYINPUT31), .B(new_n712), .C1(new_n761), .C2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT93), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(new_n765), .B2(new_n511), .ZN(new_n769));
  INV_X1    g0569(.A(new_n660), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n655), .A2(new_n560), .A3(G179), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n505), .A2(KEYINPUT93), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n505), .A2(new_n755), .A3(new_n756), .ZN(new_n774));
  AOI21_X1  g0574(.A(KEYINPUT30), .B1(new_n759), .B2(new_n511), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n713), .B1(new_n773), .B2(new_n776), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n754), .B(new_n767), .C1(new_n777), .C2(KEYINPUT31), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n769), .A2(new_n757), .A3(new_n772), .A4(new_n760), .ZN(new_n779));
  AOI21_X1  g0579(.A(KEYINPUT31), .B1(new_n779), .B2(new_n712), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n712), .A2(KEYINPUT31), .ZN(new_n781));
  INV_X1    g0581(.A(new_n766), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(KEYINPUT94), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n584), .A2(new_n685), .A3(new_n713), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n778), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G330), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n753), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n736), .B1(new_n789), .B2(G1), .ZN(G364));
  AND2_X1   g0590(.A1(new_n209), .A2(G13), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n208), .B1(new_n791), .B2(G45), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n729), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n728), .A2(new_n363), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n796), .A2(G355), .B1(new_n607), .B2(new_n728), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n728), .A2(new_n328), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n734), .B2(new_n282), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n249), .A2(new_n496), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G13), .A2(G33), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n228), .B1(G20), .B2(new_n345), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT97), .Z(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n795), .B1(new_n801), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n805), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n308), .A2(G179), .A3(G200), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n209), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n209), .A2(new_n342), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G200), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n308), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G97), .A2(new_n813), .B1(new_n816), .B2(G50), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n209), .A2(G179), .ZN(new_n818));
  NOR2_X1   g0618(.A1(G190), .A2(G200), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G159), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT32), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n818), .A2(G190), .A3(G200), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n822), .A2(new_n823), .B1(new_n825), .B2(G87), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n817), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n822), .A2(new_n823), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n815), .A2(G190), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n818), .A2(new_n308), .A3(G200), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n830), .A2(new_n245), .B1(new_n831), .B2(new_n526), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n814), .A2(new_n819), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n814), .A2(G190), .A3(new_n382), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n328), .B1(new_n833), .B2(new_n331), .C1(new_n216), .C2(new_n834), .ZN(new_n835));
  NOR4_X1   g0635(.A1(new_n827), .A2(new_n828), .A3(new_n832), .A4(new_n835), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(KEYINPUT98), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(KEYINPUT98), .ZN(new_n838));
  INV_X1    g0638(.A(new_n816), .ZN(new_n839));
  INV_X1    g0639(.A(G326), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n640), .A2(new_n642), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n839), .A2(new_n840), .B1(new_n841), .B2(new_n812), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT99), .ZN(new_n843));
  INV_X1    g0643(.A(G311), .ZN(new_n844));
  INV_X1    g0644(.A(G329), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n833), .A2(new_n844), .B1(new_n820), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n834), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n328), .B(new_n846), .C1(G322), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G317), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT33), .ZN(new_n850));
  OR2_X1    g0650(.A1(new_n849), .A2(KEYINPUT33), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n829), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n831), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n825), .A2(G303), .B1(new_n853), .B2(G283), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n843), .A2(new_n848), .A3(new_n852), .A4(new_n854), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n837), .A2(new_n838), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n804), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n809), .B1(new_n810), .B2(new_n856), .C1(new_n716), .C2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n717), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n859), .A2(new_n794), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n716), .A2(G330), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(G396));
  NOR2_X1   g0663(.A1(new_n303), .A2(new_n713), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n700), .B1(new_n310), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n347), .A2(new_n712), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n866), .A2(KEYINPUT101), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT101), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n286), .A2(new_n303), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n264), .B1(new_n263), .B2(new_n277), .ZN(new_n871));
  AND4_X1   g0671(.A1(new_n264), .A2(new_n277), .A3(new_n283), .A4(new_n281), .ZN(new_n872));
  OAI21_X1  g0672(.A(G190), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT70), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n306), .A2(new_n305), .A3(G190), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n347), .B1(new_n876), .B2(new_n864), .ZN(new_n877));
  INV_X1    g0677(.A(new_n867), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n869), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n868), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n751), .B(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(new_n787), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT102), .Z(new_n883));
  AOI21_X1  g0683(.A(new_n794), .B1(new_n881), .B2(new_n787), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n833), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n816), .A2(G303), .B1(new_n886), .B2(G116), .ZN(new_n887));
  INV_X1    g0687(.A(G283), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n887), .B1(new_n888), .B2(new_n830), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT100), .Z(new_n890));
  OAI221_X1 g0690(.A(new_n363), .B1(new_n820), .B2(new_n844), .C1(new_n834), .C2(new_n641), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n813), .A2(G97), .B1(new_n853), .B2(G87), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n526), .B2(new_n824), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n847), .A2(G143), .B1(new_n886), .B2(G159), .ZN(new_n895));
  INV_X1    g0695(.A(G137), .ZN(new_n896));
  OAI221_X1 g0696(.A(new_n895), .B1(new_n830), .B2(new_n314), .C1(new_n896), .C2(new_n839), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT34), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  INV_X1    g0700(.A(G132), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n328), .B1(new_n820), .B2(new_n901), .C1(new_n202), .C2(new_n824), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n831), .A2(new_n245), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n216), .B2(new_n812), .ZN(new_n905));
  NOR4_X1   g0705(.A1(new_n899), .A2(new_n900), .A3(new_n902), .A4(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n805), .B1(new_n894), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n805), .A2(new_n802), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n795), .B1(new_n331), .B2(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n907), .B(new_n909), .C1(new_n880), .C2(new_n803), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n885), .A2(new_n910), .ZN(G384));
  OR2_X1    g0711(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n912), .A2(G116), .A3(new_n229), .A4(new_n913), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT36), .Z(new_n915));
  OAI211_X1 g0715(.A(new_n227), .B(G77), .C1(new_n216), .C2(new_n245), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n208), .B(G13), .C1(new_n916), .C2(new_n244), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT107), .ZN(new_n919));
  INV_X1    g0719(.A(new_n710), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n409), .B1(new_n413), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n921), .B(new_n417), .C1(KEYINPUT106), .C2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n922), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n377), .A2(new_n381), .B1(new_n412), .B2(new_n710), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT106), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n377), .A2(new_n381), .A3(new_n396), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(new_n926), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n919), .B1(new_n924), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n921), .A2(new_n417), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n933), .B(new_n925), .C1(new_n927), .C2(new_n926), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(KEYINPUT107), .A3(new_n923), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n398), .A2(new_n710), .ZN(new_n936));
  INV_X1    g0736(.A(new_n416), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n419), .A2(new_n420), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n932), .A2(new_n935), .A3(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT38), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n370), .B1(new_n357), .B2(new_n371), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n288), .B(new_n943), .C1(new_n402), .C2(new_n403), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n381), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n920), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n413), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n947), .A3(new_n417), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT37), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT103), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n921), .A2(new_n417), .A3(new_n922), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT103), .ZN(new_n952));
  INV_X1    g0752(.A(new_n396), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n380), .B1(new_n369), .B2(new_n943), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n409), .A2(new_n953), .B1(new_n954), .B2(new_n710), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n412), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n952), .B(KEYINPUT37), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n950), .A2(new_n951), .A3(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n946), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n422), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n958), .A2(new_n960), .A3(KEYINPUT38), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n942), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT39), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n958), .A2(KEYINPUT38), .A3(new_n960), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT38), .B1(new_n958), .B2(new_n960), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n965), .A2(new_n966), .A3(new_n963), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n458), .A2(new_n461), .ZN(new_n969));
  INV_X1    g0769(.A(new_n432), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(new_n712), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n964), .A2(new_n968), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n867), .B1(new_n751), .B2(new_n880), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n432), .A2(new_n713), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n971), .A2(new_n465), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n975), .B1(new_n462), .B2(new_n466), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n974), .A2(new_n980), .ZN(new_n981));
  NOR3_X1   g0781(.A1(new_n965), .A2(new_n966), .A3(KEYINPUT105), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT105), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n422), .A2(new_n959), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n957), .A2(new_n951), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n952), .B1(new_n948), .B2(KEYINPUT37), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n941), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n983), .B1(new_n988), .B2(new_n961), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n981), .B1(new_n982), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n937), .A2(new_n710), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n973), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n745), .A2(new_n468), .A3(new_n752), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n705), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n992), .B(new_n994), .Z(new_n995));
  INV_X1    g0795(.A(new_n780), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n779), .A2(KEYINPUT31), .A3(new_n712), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n785), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AND4_X1   g0798(.A1(KEYINPUT40), .A2(new_n998), .A3(new_n979), .A4(new_n880), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT108), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n962), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(new_n962), .B2(new_n999), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n998), .A2(new_n979), .A3(new_n880), .ZN(new_n1003));
  OAI21_X1  g0803(.A(KEYINPUT105), .B1(new_n965), .B2(new_n966), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n988), .A2(new_n983), .A3(new_n961), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n1001), .A2(new_n1002), .B1(new_n1006), .B2(KEYINPUT40), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n468), .A2(new_n998), .ZN(new_n1008));
  OAI21_X1  g0808(.A(G330), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n1008), .B2(new_n1007), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n995), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n995), .A2(new_n1010), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT109), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1011), .B1(new_n208), .B2(new_n791), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1012), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(KEYINPUT109), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n918), .B1(new_n1014), .B2(new_n1016), .ZN(G367));
  INV_X1    g0817(.A(new_n544), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n533), .A2(new_n544), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n543), .A2(new_n712), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT110), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1019), .A2(new_n1023), .A3(new_n1020), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1018), .B1(new_n1025), .B2(new_n689), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(new_n712), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT42), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1018), .A2(new_n712), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1022), .A2(new_n1029), .A3(new_n1024), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n724), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT43), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n712), .B1(new_n574), .B2(new_n579), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n583), .A2(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n578), .A2(new_n1035), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1030), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1033), .A2(new_n1034), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1032), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1042), .B(new_n1040), .C1(new_n712), .C2(new_n1026), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1039), .A2(new_n1034), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1038), .A2(KEYINPUT43), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1030), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n723), .A2(new_n1047), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1041), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1048), .B1(new_n1041), .B2(new_n1046), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n729), .B(KEYINPUT41), .Z(new_n1052));
  INV_X1    g0852(.A(KEYINPUT44), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n725), .B1(KEYINPUT111), .B2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1047), .B(new_n1054), .C1(KEYINPUT111), .C2(new_n1053), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT111), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1056), .B(KEYINPUT44), .C1(new_n1030), .C2(new_n725), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1030), .A2(new_n725), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT45), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(KEYINPUT45), .B1(new_n1030), .B2(new_n725), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1055), .B(new_n1057), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n722), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1058), .B(new_n1059), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1064), .A2(new_n723), .A3(new_n1057), .A4(new_n1055), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n712), .B1(new_n670), .B2(new_n672), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n721), .B(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(new_n859), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n788), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1063), .A2(new_n1065), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1052), .B1(new_n1070), .B2(new_n789), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1051), .B1(new_n1071), .B2(new_n793), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n808), .B1(new_n212), .B2(new_n576), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n798), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(new_n239), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n794), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n833), .A2(new_n202), .B1(new_n820), .B2(new_n896), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n363), .B(new_n1077), .C1(G150), .C2(new_n847), .ZN(new_n1078));
  INV_X1    g0878(.A(G143), .ZN(new_n1079));
  OAI221_X1 g0879(.A(new_n1078), .B1(new_n1079), .B2(new_n839), .C1(new_n821), .C2(new_n830), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n853), .A2(G77), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1081), .B1(new_n216), .B2(new_n824), .C1(new_n245), .C2(new_n812), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n841), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n829), .A2(new_n1083), .B1(new_n853), .B2(G97), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1084), .B1(new_n526), .B2(new_n812), .C1(new_n844), .C2(new_n839), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n820), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n847), .A2(G303), .B1(new_n1086), .B2(G317), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT46), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n824), .B2(new_n607), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n825), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n328), .B1(new_n886), .B2(G283), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1080), .A2(new_n1082), .B1(new_n1085), .B2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT47), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1076), .B1(new_n1094), .B2(new_n805), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n857), .B2(new_n1038), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1072), .A2(new_n1096), .ZN(G387));
  NAND2_X1  g0897(.A1(new_n788), .A2(new_n1068), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1069), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1098), .A2(new_n1099), .A3(new_n729), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n798), .B1(new_n236), .B2(new_n252), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n796), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1101), .B1(new_n732), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n290), .A2(G50), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT50), .ZN(new_n1105));
  AOI21_X1  g0905(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n732), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1103), .A2(new_n1107), .B1(new_n526), .B2(new_n728), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n794), .B1(new_n1108), .B2(new_n807), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n847), .A2(G317), .B1(new_n886), .B2(G303), .ZN(new_n1110));
  INV_X1    g0910(.A(G322), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1110), .B1(new_n830), .B2(new_n844), .C1(new_n1111), .C2(new_n839), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT48), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n813), .A2(G283), .B1(new_n1083), .B2(new_n825), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1118), .A2(KEYINPUT49), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n363), .B1(new_n820), .B2(new_n840), .C1(new_n607), .C2(new_n831), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1121), .B1(KEYINPUT49), .B2(new_n1118), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n813), .A2(new_n294), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n202), .B2(new_n834), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT112), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n328), .B1(new_n820), .B2(new_n314), .C1(new_n245), .C2(new_n833), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n830), .A2(new_n290), .B1(new_n218), .B2(new_n831), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n839), .A2(new_n821), .B1(new_n824), .B2(new_n331), .ZN(new_n1128));
  OR4_X1    g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n810), .B1(new_n1122), .B2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1109), .B(new_n1130), .C1(new_n721), .C2(new_n804), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1068), .B2(new_n792), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1100), .A2(new_n1134), .ZN(G393));
  NAND2_X1  g0935(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n1099), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1137), .A2(new_n729), .A3(new_n1070), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1063), .A2(new_n1065), .A3(new_n793), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n808), .B1(new_n218), .B2(new_n212), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n1074), .A2(new_n243), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n794), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n839), .A2(new_n849), .B1(new_n844), .B2(new_n834), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT52), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n824), .A2(new_n888), .B1(new_n820), .B2(new_n1111), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT113), .Z(new_n1146));
  OAI21_X1  g0946(.A(new_n363), .B1(new_n833), .B2(new_n641), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G107), .B2(new_n853), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G116), .A2(new_n813), .B1(new_n829), .B2(G303), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT114), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G150), .A2(new_n816), .B1(new_n847), .B2(G159), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT51), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n328), .B1(new_n820), .B2(new_n1079), .C1(new_n290), .C2(new_n833), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n830), .A2(new_n202), .B1(new_n831), .B2(new_n385), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n812), .A2(new_n331), .B1(new_n824), .B2(new_n245), .ZN(new_n1157));
  OR4_X1    g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1152), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1142), .B1(new_n1160), .B2(new_n805), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n1030), .B2(new_n857), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1138), .A2(new_n1139), .A3(new_n1162), .ZN(G390));
  NAND2_X1  g0963(.A1(new_n979), .A2(new_n880), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n996), .A2(new_n997), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n659), .A2(new_n684), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n687), .A2(new_n1166), .A3(new_n712), .ZN(new_n1167));
  OAI21_X1  g0967(.A(G330), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1164), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n713), .B1(new_n698), .B2(new_n692), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n879), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n877), .A2(new_n869), .A3(new_n878), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n878), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n979), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n972), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n964), .A2(new_n968), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n713), .B(new_n880), .C1(new_n740), .C2(new_n744), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n980), .B1(new_n1178), .B2(new_n878), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n962), .A2(new_n1176), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1169), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT39), .B1(new_n942), .B2(new_n961), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n972), .A2(new_n981), .B1(new_n1183), .B2(new_n967), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n786), .A2(G330), .A3(new_n880), .A4(new_n979), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT115), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1185), .B(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1184), .B(new_n1187), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1182), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n802), .B1(new_n1183), .B2(new_n967), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n824), .A2(new_n385), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n839), .A2(new_n888), .B1(new_n331), .B2(new_n812), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n363), .B1(new_n820), .B2(new_n641), .C1(new_n834), .C2(new_n607), .ZN(new_n1194));
  OR4_X1    g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n903), .A4(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n829), .A2(G107), .B1(new_n886), .B2(G97), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT119), .Z(new_n1197));
  NAND2_X1  g0997(.A1(new_n825), .A2(G150), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT53), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G159), .A2(new_n813), .B1(new_n829), .B2(G137), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n816), .A2(G128), .B1(new_n853), .B2(G50), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT54), .B(G143), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n363), .B1(new_n886), .B2(new_n1203), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n847), .A2(G132), .B1(new_n1086), .B2(G125), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1200), .A2(new_n1201), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n1195), .A2(new_n1197), .B1(new_n1199), .B2(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1207), .A2(new_n805), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n795), .B(new_n1208), .C1(new_n290), .C2(new_n908), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1190), .A2(new_n793), .B1(new_n1191), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n786), .A2(G330), .A3(new_n880), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n980), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT116), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1169), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT116), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1211), .A2(new_n1215), .A3(new_n980), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n980), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(new_n1178), .A3(new_n878), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1217), .A2(new_n1174), .B1(new_n1187), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n468), .A2(G330), .A3(new_n998), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n993), .A2(new_n1222), .A3(new_n705), .ZN(new_n1223));
  OAI21_X1  g1023(.A(KEYINPUT118), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT118), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1223), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1169), .B1(new_n1212), .B2(KEYINPUT116), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n974), .B1(new_n1227), .B2(new_n1216), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1219), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1225), .B(new_n1226), .C1(new_n1228), .C2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1224), .A2(new_n1189), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT117), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1226), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1234), .B(new_n729), .C1(new_n1189), .C2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1217), .A2(new_n1174), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1187), .A2(new_n1220), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1240), .A2(new_n1188), .A3(new_n1182), .A4(new_n1226), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1234), .B1(new_n1241), .B2(new_n729), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1210), .B1(new_n1237), .B2(new_n1242), .ZN(G378));
  NAND2_X1  g1043(.A1(new_n271), .A2(new_n253), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT120), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n202), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n253), .B2(new_n363), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n839), .A2(new_n607), .B1(new_n831), .B2(new_n216), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G97), .B2(new_n829), .ZN(new_n1249));
  AOI211_X1 g1049(.A(G41), .B(new_n328), .C1(new_n1086), .C2(G283), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n847), .A2(G107), .B1(new_n886), .B2(new_n294), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n813), .A2(G68), .B1(new_n825), .B2(G77), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT58), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1247), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1245), .B1(G124), .B2(new_n1086), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n816), .A2(G125), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n830), .B2(new_n901), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n847), .A2(G128), .B1(new_n886), .B2(G137), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n824), .B2(new_n1202), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1258), .B(new_n1260), .C1(G150), .C2(new_n813), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT59), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1256), .B1(new_n821), .B2(new_n831), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1261), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(KEYINPUT59), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1255), .B1(new_n1254), .B2(new_n1253), .C1(new_n1263), .C2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n805), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n795), .B1(new_n202), .B2(new_n908), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n341), .A2(new_n349), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n319), .A2(new_n710), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1269), .B(new_n1270), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1271), .B(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1267), .B(new_n1268), .C1(new_n1274), .C2(new_n803), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT40), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1003), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n982), .B2(new_n989), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n965), .B1(new_n941), .B2(new_n940), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n998), .A2(new_n979), .A3(new_n880), .A4(KEYINPUT40), .ZN(new_n1281));
  OAI21_X1  g1081(.A(KEYINPUT108), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n962), .A2(new_n999), .A3(new_n1000), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n1277), .A2(new_n1279), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1274), .B1(new_n1284), .B2(G330), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1279), .A2(new_n1277), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1287));
  AND4_X1   g1087(.A1(G330), .A2(new_n1286), .A3(new_n1287), .A4(new_n1274), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n992), .B1(new_n1285), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(G330), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1273), .B1(new_n1007), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n992), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1286), .A2(new_n1287), .A3(new_n1274), .A4(G330), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1289), .A2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1276), .B1(new_n1295), .B2(new_n793), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1226), .B1(new_n1189), .B2(new_n1221), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1292), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1299));
  OAI211_X1 g1099(.A(KEYINPUT57), .B(new_n1297), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n729), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT57), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1296), .B1(new_n1301), .B2(new_n1302), .ZN(G375));
  AOI21_X1  g1103(.A(new_n792), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n980), .A2(new_n802), .ZN(new_n1305));
  OAI22_X1  g1105(.A1(new_n607), .A2(new_n830), .B1(new_n839), .B2(new_n641), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1306), .B1(G97), .B2(new_n825), .ZN(new_n1307));
  OAI22_X1  g1107(.A1(new_n834), .A2(new_n888), .B1(new_n833), .B2(new_n526), .ZN(new_n1308));
  AOI211_X1 g1108(.A(new_n328), .B(new_n1308), .C1(G303), .C2(new_n1086), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1307), .A2(new_n1081), .A3(new_n1123), .A4(new_n1309), .ZN(new_n1310));
  OAI22_X1  g1110(.A1(new_n812), .A2(new_n202), .B1(new_n824), .B2(new_n821), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(G132), .B2(new_n816), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n363), .B1(new_n1086), .B2(G128), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n847), .A2(G137), .B1(new_n886), .B2(G150), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n829), .A2(new_n1203), .B1(new_n853), .B2(G58), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .A4(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n810), .B1(new_n1310), .B2(new_n1316), .ZN(new_n1317));
  AOI211_X1 g1117(.A(new_n795), .B(new_n1317), .C1(new_n245), .C2(new_n908), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1305), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT121), .B1(new_n1304), .B2(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n793), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT121), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1322), .A2(new_n1323), .A3(new_n1319), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1224), .A2(new_n1232), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1052), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1325), .B1(new_n1326), .B2(new_n1329), .ZN(G381));
  INV_X1    g1130(.A(G375), .ZN(new_n1331));
  INV_X1    g1131(.A(G378), .ZN(new_n1332));
  INV_X1    g1132(.A(G390), .ZN(new_n1333));
  INV_X1    g1133(.A(G384), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(G393), .A2(G396), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  NOR3_X1   g1136(.A1(new_n1336), .A2(G387), .A3(G381), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1331), .A2(new_n1332), .A3(new_n1337), .ZN(G407));
  NAND2_X1  g1138(.A1(new_n711), .A2(G213), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(new_n1339), .B(KEYINPUT122), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1331), .A2(new_n1332), .A3(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(G407), .A2(new_n1341), .A3(G213), .ZN(G409));
  INV_X1    g1142(.A(KEYINPUT127), .ZN(new_n1343));
  OAI211_X1 g1143(.A(G378), .B(new_n1296), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1328), .B(new_n1297), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n793), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1345), .A2(new_n1346), .A3(new_n1275), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1241), .A2(new_n729), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(KEYINPUT117), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1349), .A2(new_n1233), .A3(new_n1236), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1347), .A2(new_n1350), .A3(new_n1210), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1344), .A2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1340), .ZN(new_n1353));
  NOR3_X1   g1153(.A1(new_n1228), .A2(new_n1226), .A3(new_n1231), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1354), .B1(KEYINPUT60), .B2(new_n1235), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1238), .A2(KEYINPUT60), .A3(new_n1223), .A4(new_n1239), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n729), .ZN(new_n1357));
  AND3_X1   g1157(.A1(new_n1322), .A2(new_n1323), .A3(new_n1319), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1323), .B1(new_n1322), .B2(new_n1319), .ZN(new_n1359));
  OAI22_X1  g1159(.A1(new_n1355), .A2(new_n1357), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(new_n1334), .ZN(new_n1361));
  AND2_X1   g1161(.A1(new_n1356), .A2(new_n729), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1223), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT60), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1327), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1362), .A2(new_n1365), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1366), .A2(new_n1325), .A3(G384), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1361), .A2(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1368), .ZN(new_n1369));
  NAND4_X1  g1169(.A1(new_n1352), .A2(KEYINPUT62), .A3(new_n1353), .A4(new_n1369), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1339), .ZN(new_n1371));
  AOI211_X1 g1171(.A(new_n1371), .B(new_n1368), .C1(new_n1344), .C2(new_n1351), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1370), .B1(new_n1372), .B2(KEYINPUT62), .ZN(new_n1373));
  INV_X1    g1173(.A(KEYINPUT125), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1340), .A2(G2897), .ZN(new_n1375));
  INV_X1    g1175(.A(new_n1375), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1366), .A2(new_n1325), .A3(G384), .ZN(new_n1377));
  AOI21_X1  g1177(.A(G384), .B1(new_n1366), .B2(new_n1325), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1376), .B1(new_n1377), .B2(new_n1378), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1371), .A2(G2897), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1361), .A2(new_n1367), .A3(new_n1380), .ZN(new_n1381));
  NAND3_X1  g1181(.A1(new_n1379), .A2(new_n1381), .A3(KEYINPUT123), .ZN(new_n1382));
  INV_X1    g1182(.A(KEYINPUT123), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(new_n1368), .A2(new_n1383), .A3(new_n1376), .ZN(new_n1384));
  NAND2_X1  g1184(.A1(new_n1382), .A2(new_n1384), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1352), .A2(new_n1353), .ZN(new_n1386));
  AOI21_X1  g1186(.A(KEYINPUT61), .B1(new_n1385), .B2(new_n1386), .ZN(new_n1387));
  AND3_X1   g1187(.A1(new_n1373), .A2(new_n1374), .A3(new_n1387), .ZN(new_n1388));
  AOI21_X1  g1188(.A(new_n1374), .B1(new_n1373), .B2(new_n1387), .ZN(new_n1389));
  AND2_X1   g1189(.A1(G393), .A2(G396), .ZN(new_n1390));
  NOR2_X1   g1190(.A1(new_n1390), .A2(new_n1335), .ZN(new_n1391));
  INV_X1    g1191(.A(new_n1391), .ZN(new_n1392));
  AND3_X1   g1192(.A1(G390), .A2(new_n1072), .A3(new_n1096), .ZN(new_n1393));
  AOI21_X1  g1193(.A(G390), .B1(new_n1072), .B2(new_n1096), .ZN(new_n1394));
  OAI21_X1  g1194(.A(new_n1392), .B1(new_n1393), .B2(new_n1394), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(G387), .A2(new_n1333), .ZN(new_n1396));
  NAND3_X1  g1196(.A1(G390), .A2(new_n1072), .A3(new_n1096), .ZN(new_n1397));
  NAND3_X1  g1197(.A1(new_n1396), .A2(new_n1391), .A3(new_n1397), .ZN(new_n1398));
  AND2_X1   g1198(.A1(new_n1395), .A2(new_n1398), .ZN(new_n1399));
  XNOR2_X1  g1199(.A(new_n1399), .B(KEYINPUT126), .ZN(new_n1400));
  INV_X1    g1200(.A(new_n1400), .ZN(new_n1401));
  NOR3_X1   g1201(.A1(new_n1388), .A2(new_n1389), .A3(new_n1401), .ZN(new_n1402));
  NAND3_X1  g1202(.A1(new_n1352), .A2(new_n1339), .A3(new_n1369), .ZN(new_n1403));
  INV_X1    g1203(.A(KEYINPUT63), .ZN(new_n1404));
  NAND2_X1  g1204(.A1(new_n1403), .A2(new_n1404), .ZN(new_n1405));
  NAND2_X1  g1205(.A1(new_n1352), .A2(new_n1339), .ZN(new_n1406));
  NAND2_X1  g1206(.A1(new_n1385), .A2(new_n1406), .ZN(new_n1407));
  INV_X1    g1207(.A(KEYINPUT61), .ZN(new_n1408));
  NAND3_X1  g1208(.A1(new_n1395), .A2(new_n1398), .A3(new_n1408), .ZN(new_n1409));
  AOI21_X1  g1209(.A(new_n1340), .B1(new_n1344), .B2(new_n1351), .ZN(new_n1410));
  NOR2_X1   g1210(.A1(new_n1368), .A2(new_n1404), .ZN(new_n1411));
  AOI21_X1  g1211(.A(new_n1409), .B1(new_n1410), .B2(new_n1411), .ZN(new_n1412));
  NAND3_X1  g1212(.A1(new_n1405), .A2(new_n1407), .A3(new_n1412), .ZN(new_n1413));
  XNOR2_X1  g1213(.A(new_n1413), .B(KEYINPUT124), .ZN(new_n1414));
  OAI21_X1  g1214(.A(new_n1343), .B1(new_n1402), .B2(new_n1414), .ZN(new_n1415));
  INV_X1    g1215(.A(KEYINPUT124), .ZN(new_n1416));
  XNOR2_X1  g1216(.A(new_n1413), .B(new_n1416), .ZN(new_n1417));
  NAND2_X1  g1217(.A1(new_n1373), .A2(new_n1387), .ZN(new_n1418));
  NAND2_X1  g1218(.A1(new_n1418), .A2(KEYINPUT125), .ZN(new_n1419));
  NAND3_X1  g1219(.A1(new_n1373), .A2(new_n1387), .A3(new_n1374), .ZN(new_n1420));
  NAND3_X1  g1220(.A1(new_n1419), .A2(new_n1420), .A3(new_n1400), .ZN(new_n1421));
  NAND3_X1  g1221(.A1(new_n1417), .A2(new_n1421), .A3(KEYINPUT127), .ZN(new_n1422));
  NAND2_X1  g1222(.A1(new_n1415), .A2(new_n1422), .ZN(G405));
  NOR2_X1   g1223(.A1(new_n1331), .A2(G378), .ZN(new_n1424));
  INV_X1    g1224(.A(new_n1424), .ZN(new_n1425));
  NAND2_X1  g1225(.A1(new_n1425), .A2(new_n1344), .ZN(new_n1426));
  XNOR2_X1  g1226(.A(new_n1426), .B(new_n1368), .ZN(new_n1427));
  XNOR2_X1  g1227(.A(new_n1427), .B(new_n1399), .ZN(G402));
endmodule


