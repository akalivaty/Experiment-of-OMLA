

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606;

  XNOR2_X1 U325 ( .A(n309), .B(n308), .ZN(n311) );
  XNOR2_X1 U326 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U327 ( .A(n484), .B(n483), .ZN(n567) );
  XNOR2_X1 U328 ( .A(n482), .B(KEYINPUT48), .ZN(n483) );
  XNOR2_X1 U329 ( .A(n357), .B(G71GAT), .ZN(n358) );
  XNOR2_X1 U330 ( .A(n465), .B(KEYINPUT107), .ZN(n548) );
  XOR2_X2 U331 ( .A(n346), .B(n345), .Z(n580) );
  XOR2_X1 U332 ( .A(KEYINPUT97), .B(n455), .Z(n293) );
  XNOR2_X1 U333 ( .A(n307), .B(n306), .ZN(n308) );
  INV_X1 U334 ( .A(KEYINPUT111), .ZN(n482) );
  XNOR2_X1 U335 ( .A(n383), .B(KEYINPUT26), .ZN(n384) );
  NOR2_X1 U336 ( .A1(n432), .A2(n431), .ZN(n513) );
  XNOR2_X1 U337 ( .A(n385), .B(n384), .ZN(n502) );
  XNOR2_X1 U338 ( .A(n298), .B(n297), .ZN(n344) );
  XNOR2_X1 U339 ( .A(n316), .B(n315), .ZN(n596) );
  INV_X1 U340 ( .A(G106GAT), .ZN(n466) );
  XNOR2_X1 U341 ( .A(n457), .B(n456), .ZN(n530) );
  XNOR2_X1 U342 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U343 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U344 ( .A(n462), .B(G50GAT), .ZN(n463) );
  XNOR2_X1 U345 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U346 ( .A(n500), .B(n499), .ZN(G1351GAT) );
  XNOR2_X1 U347 ( .A(n464), .B(n463), .ZN(G1331GAT) );
  XOR2_X1 U348 ( .A(KEYINPUT98), .B(KEYINPUT38), .Z(n457) );
  XNOR2_X1 U349 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n294) );
  XNOR2_X1 U350 ( .A(n294), .B(G29GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(G50GAT), .ZN(n296) );
  INV_X1 U352 ( .A(KEYINPUT7), .ZN(n295) );
  XNOR2_X1 U353 ( .A(G22GAT), .B(G197GAT), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n299), .B(G141GAT), .ZN(n378) );
  XNOR2_X1 U355 ( .A(n344), .B(n378), .ZN(n303) );
  INV_X1 U356 ( .A(n303), .ZN(n301) );
  XOR2_X1 U357 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n302) );
  INV_X1 U358 ( .A(n302), .ZN(n300) );
  NAND2_X1 U359 ( .A1(n301), .A2(n300), .ZN(n305) );
  NAND2_X1 U360 ( .A1(n303), .A2(n302), .ZN(n304) );
  NAND2_X1 U361 ( .A1(n305), .A2(n304), .ZN(n309) );
  XOR2_X1 U362 ( .A(G169GAT), .B(G8GAT), .Z(n388) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(n388), .ZN(n307) );
  INV_X1 U364 ( .A(KEYINPUT29), .ZN(n306) );
  INV_X1 U365 ( .A(n311), .ZN(n310) );
  XOR2_X1 U366 ( .A(G15GAT), .B(G1GAT), .Z(n436) );
  NAND2_X1 U367 ( .A1(n310), .A2(n436), .ZN(n314) );
  INV_X1 U368 ( .A(n436), .ZN(n312) );
  NAND2_X1 U369 ( .A1(n312), .A2(n311), .ZN(n313) );
  NAND2_X1 U370 ( .A1(n314), .A2(n313), .ZN(n316) );
  NAND2_X1 U371 ( .A1(G229GAT), .A2(G233GAT), .ZN(n315) );
  XOR2_X1 U372 ( .A(KEYINPUT67), .B(n596), .Z(n550) );
  XOR2_X1 U373 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n318) );
  NAND2_X1 U374 ( .A1(G230GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U376 ( .A(n319), .B(KEYINPUT33), .Z(n323) );
  XNOR2_X1 U377 ( .A(G71GAT), .B(G57GAT), .ZN(n320) );
  XNOR2_X1 U378 ( .A(n320), .B(KEYINPUT13), .ZN(n435) );
  XNOR2_X1 U379 ( .A(G176GAT), .B(G92GAT), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n321), .B(G64GAT), .ZN(n392) );
  XNOR2_X1 U381 ( .A(n435), .B(n392), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U383 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n325) );
  XNOR2_X1 U384 ( .A(G120GAT), .B(KEYINPUT72), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U386 ( .A(n327), .B(n326), .Z(n333) );
  XOR2_X1 U387 ( .A(G78GAT), .B(G148GAT), .Z(n329) );
  XNOR2_X1 U388 ( .A(KEYINPUT69), .B(G204GAT), .ZN(n328) );
  XNOR2_X1 U389 ( .A(n329), .B(n328), .ZN(n373) );
  XOR2_X1 U390 ( .A(G85GAT), .B(KEYINPUT70), .Z(n331) );
  XNOR2_X1 U391 ( .A(G99GAT), .B(G106GAT), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n373), .B(n336), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n600) );
  NOR2_X1 U395 ( .A1(n550), .A2(n600), .ZN(n515) );
  XOR2_X1 U396 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n335) );
  XNOR2_X1 U397 ( .A(G92GAT), .B(KEYINPUT73), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n343) );
  XOR2_X1 U399 ( .A(G218GAT), .B(G162GAT), .Z(n377) );
  XOR2_X1 U400 ( .A(n336), .B(n377), .Z(n338) );
  NAND2_X1 U401 ( .A1(G232GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U403 ( .A(n339), .B(KEYINPUT64), .Z(n341) );
  XOR2_X1 U404 ( .A(G190GAT), .B(G134GAT), .Z(n356) );
  XNOR2_X1 U405 ( .A(n356), .B(KEYINPUT11), .ZN(n340) );
  XNOR2_X1 U406 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U407 ( .A(n343), .B(n342), .ZN(n346) );
  INV_X1 U408 ( .A(n344), .ZN(n345) );
  INV_X1 U409 ( .A(n580), .ZN(n509) );
  XNOR2_X1 U410 ( .A(KEYINPUT36), .B(n509), .ZN(n505) );
  INV_X1 U411 ( .A(KEYINPUT90), .ZN(n406) );
  XOR2_X1 U412 ( .A(KEYINPUT77), .B(G120GAT), .Z(n348) );
  XNOR2_X1 U413 ( .A(G113GAT), .B(G127GAT), .ZN(n347) );
  XNOR2_X1 U414 ( .A(n348), .B(n347), .ZN(n350) );
  XOR2_X1 U415 ( .A(KEYINPUT0), .B(KEYINPUT78), .Z(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n423) );
  XOR2_X1 U417 ( .A(KEYINPUT80), .B(G176GAT), .Z(n352) );
  XNOR2_X1 U418 ( .A(G169GAT), .B(G15GAT), .ZN(n351) );
  XNOR2_X1 U419 ( .A(n352), .B(n351), .ZN(n365) );
  XOR2_X1 U420 ( .A(KEYINPUT79), .B(KEYINPUT65), .Z(n354) );
  XNOR2_X1 U421 ( .A(G43GAT), .B(G99GAT), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U423 ( .A(n356), .B(n355), .ZN(n359) );
  AND2_X1 U424 ( .A1(G227GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U426 ( .A(G183GAT), .B(KEYINPUT18), .Z(n361) );
  XNOR2_X1 U427 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n360) );
  XNOR2_X1 U428 ( .A(n361), .B(n360), .ZN(n393) );
  XOR2_X1 U429 ( .A(n393), .B(KEYINPUT20), .Z(n362) );
  XNOR2_X1 U430 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U431 ( .A(n365), .B(n364), .Z(n366) );
  XOR2_X2 U432 ( .A(n423), .B(n366), .Z(n551) );
  XOR2_X1 U433 ( .A(KEYINPUT81), .B(KEYINPUT23), .Z(n368) );
  XNOR2_X1 U434 ( .A(G50GAT), .B(G106GAT), .ZN(n367) );
  XNOR2_X1 U435 ( .A(n368), .B(n367), .ZN(n382) );
  XOR2_X1 U436 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n370) );
  NAND2_X1 U437 ( .A1(G228GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U439 ( .A(n371), .B(KEYINPUT82), .Z(n375) );
  XNOR2_X1 U440 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n372) );
  XNOR2_X1 U441 ( .A(n372), .B(KEYINPUT2), .ZN(n418) );
  XNOR2_X1 U442 ( .A(n418), .B(n373), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U444 ( .A(KEYINPUT21), .B(G211GAT), .Z(n397) );
  XOR2_X1 U445 ( .A(n376), .B(n397), .Z(n380) );
  XNOR2_X1 U446 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U447 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n382), .B(n381), .ZN(n491) );
  NOR2_X1 U449 ( .A1(n551), .A2(n491), .ZN(n385) );
  INV_X1 U450 ( .A(KEYINPUT87), .ZN(n383) );
  XOR2_X1 U451 ( .A(KEYINPUT86), .B(G204GAT), .Z(n387) );
  XNOR2_X1 U452 ( .A(G197GAT), .B(G190GAT), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n391) );
  XNOR2_X1 U454 ( .A(G36GAT), .B(n388), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n389), .B(G218GAT), .ZN(n390) );
  XOR2_X1 U456 ( .A(n391), .B(n390), .Z(n395) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U459 ( .A(n397), .B(n396), .Z(n399) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n546) );
  XNOR2_X1 U462 ( .A(n546), .B(KEYINPUT27), .ZN(n428) );
  NAND2_X1 U463 ( .A1(n502), .A2(n428), .ZN(n569) );
  XNOR2_X1 U464 ( .A(KEYINPUT89), .B(KEYINPUT25), .ZN(n403) );
  NAND2_X1 U465 ( .A1(n551), .A2(n546), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n400), .B(KEYINPUT88), .ZN(n401) );
  NAND2_X1 U467 ( .A1(n401), .A2(n491), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n403), .B(n402), .ZN(n404) );
  NAND2_X1 U469 ( .A1(n569), .A2(n404), .ZN(n405) );
  XNOR2_X1 U470 ( .A(n406), .B(n405), .ZN(n427) );
  XOR2_X1 U471 ( .A(G57GAT), .B(G148GAT), .Z(n408) );
  XNOR2_X1 U472 ( .A(G1GAT), .B(G141GAT), .ZN(n407) );
  XNOR2_X1 U473 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U474 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n410) );
  XNOR2_X1 U475 ( .A(KEYINPUT84), .B(KEYINPUT6), .ZN(n409) );
  XNOR2_X1 U476 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U477 ( .A(n412), .B(n411), .Z(n417) );
  XOR2_X1 U478 ( .A(KEYINPUT4), .B(KEYINPUT85), .Z(n414) );
  NAND2_X1 U479 ( .A1(G225GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U480 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U481 ( .A(KEYINPUT83), .B(n415), .ZN(n416) );
  XNOR2_X1 U482 ( .A(n417), .B(n416), .ZN(n422) );
  XOR2_X1 U483 ( .A(G85GAT), .B(G162GAT), .Z(n420) );
  XNOR2_X1 U484 ( .A(G29GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U485 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U486 ( .A(n422), .B(n421), .Z(n426) );
  INV_X1 U487 ( .A(n423), .ZN(n424) );
  XNOR2_X1 U488 ( .A(n424), .B(G134GAT), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n566) );
  NOR2_X1 U490 ( .A1(n427), .A2(n566), .ZN(n432) );
  INV_X1 U491 ( .A(n428), .ZN(n429) );
  XOR2_X1 U492 ( .A(KEYINPUT28), .B(n491), .Z(n541) );
  NOR2_X1 U493 ( .A1(n429), .A2(n541), .ZN(n430) );
  NAND2_X1 U494 ( .A1(n566), .A2(n430), .ZN(n553) );
  NOR2_X1 U495 ( .A1(n551), .A2(n553), .ZN(n431) );
  XOR2_X1 U496 ( .A(G211GAT), .B(G78GAT), .Z(n434) );
  XNOR2_X1 U497 ( .A(G22GAT), .B(G155GAT), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n449) );
  XOR2_X1 U499 ( .A(n435), .B(G183GAT), .Z(n438) );
  XNOR2_X1 U500 ( .A(n436), .B(G127GAT), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U502 ( .A(KEYINPUT75), .B(KEYINPUT12), .Z(n440) );
  NAND2_X1 U503 ( .A1(G231GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U504 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U505 ( .A(n442), .B(n441), .Z(n447) );
  XOR2_X1 U506 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n444) );
  XNOR2_X1 U507 ( .A(G8GAT), .B(G64GAT), .ZN(n443) );
  XNOR2_X1 U508 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U509 ( .A(n445), .B(KEYINPUT74), .ZN(n446) );
  XNOR2_X1 U510 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U511 ( .A(n449), .B(n448), .Z(n470) );
  INV_X1 U512 ( .A(n470), .ZN(n603) );
  NOR2_X1 U513 ( .A1(n513), .A2(n603), .ZN(n451) );
  INV_X1 U514 ( .A(KEYINPUT96), .ZN(n450) );
  XNOR2_X1 U515 ( .A(n451), .B(n450), .ZN(n452) );
  NOR2_X1 U516 ( .A1(n505), .A2(n452), .ZN(n454) );
  INV_X1 U517 ( .A(KEYINPUT37), .ZN(n453) );
  XNOR2_X1 U518 ( .A(n454), .B(n453), .ZN(n455) );
  NAND2_X1 U519 ( .A1(n515), .A2(n293), .ZN(n456) );
  NAND2_X1 U520 ( .A1(n530), .A2(n551), .ZN(n461) );
  XOR2_X1 U521 ( .A(KEYINPUT101), .B(KEYINPUT40), .Z(n459) );
  XNOR2_X1 U522 ( .A(G43GAT), .B(KEYINPUT100), .ZN(n458) );
  XNOR2_X1 U523 ( .A(n461), .B(n460), .ZN(G1330GAT) );
  NAND2_X1 U524 ( .A1(n530), .A2(n541), .ZN(n464) );
  XOR2_X1 U525 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n462) );
  INV_X1 U526 ( .A(n596), .ZN(n571) );
  XNOR2_X1 U527 ( .A(n600), .B(KEYINPUT41), .ZN(n555) );
  NOR2_X1 U528 ( .A1(n571), .A2(n555), .ZN(n533) );
  NAND2_X1 U529 ( .A1(n533), .A2(n293), .ZN(n465) );
  NAND2_X1 U530 ( .A1(n548), .A2(n541), .ZN(n469) );
  XOR2_X1 U531 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n467) );
  XNOR2_X1 U532 ( .A(n469), .B(n468), .ZN(G1339GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT54), .B(KEYINPUT119), .Z(n486) );
  NOR2_X1 U534 ( .A1(n505), .A2(n470), .ZN(n471) );
  XOR2_X1 U535 ( .A(KEYINPUT45), .B(n471), .Z(n472) );
  NOR2_X1 U536 ( .A1(n600), .A2(n472), .ZN(n473) );
  NAND2_X1 U537 ( .A1(n473), .A2(n550), .ZN(n481) );
  NOR2_X1 U538 ( .A1(n596), .A2(n555), .ZN(n474) );
  XNOR2_X1 U539 ( .A(n474), .B(KEYINPUT46), .ZN(n475) );
  NOR2_X1 U540 ( .A1(n603), .A2(n475), .ZN(n476) );
  XNOR2_X1 U541 ( .A(n476), .B(KEYINPUT109), .ZN(n477) );
  NOR2_X1 U542 ( .A1(n477), .A2(n580), .ZN(n478) );
  XNOR2_X1 U543 ( .A(n478), .B(KEYINPUT110), .ZN(n479) );
  XNOR2_X1 U544 ( .A(n479), .B(KEYINPUT47), .ZN(n480) );
  NAND2_X1 U545 ( .A1(n481), .A2(n480), .ZN(n484) );
  NAND2_X1 U546 ( .A1(n546), .A2(n567), .ZN(n485) );
  NAND2_X1 U547 ( .A1(n486), .A2(n485), .ZN(n490) );
  INV_X1 U548 ( .A(n485), .ZN(n488) );
  INV_X1 U549 ( .A(n486), .ZN(n487) );
  NAND2_X1 U550 ( .A1(n488), .A2(n487), .ZN(n489) );
  NAND2_X1 U551 ( .A1(n490), .A2(n489), .ZN(n501) );
  INV_X1 U552 ( .A(n491), .ZN(n492) );
  OR2_X1 U553 ( .A1(n566), .A2(n492), .ZN(n493) );
  NOR2_X1 U554 ( .A1(n501), .A2(n493), .ZN(n494) );
  XNOR2_X1 U555 ( .A(KEYINPUT55), .B(n494), .ZN(n496) );
  INV_X1 U556 ( .A(n551), .ZN(n495) );
  NOR2_X1 U557 ( .A1(n496), .A2(n495), .ZN(n590) );
  NAND2_X1 U558 ( .A1(n590), .A2(n580), .ZN(n500) );
  XOR2_X1 U559 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n498) );
  XNOR2_X1 U560 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n497) );
  NOR2_X1 U561 ( .A1(n501), .A2(n566), .ZN(n503) );
  NAND2_X1 U562 ( .A1(n503), .A2(n502), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n504), .B(KEYINPUT124), .ZN(n599) );
  NOR2_X1 U564 ( .A1(n599), .A2(n505), .ZN(n506) );
  XNOR2_X1 U565 ( .A(KEYINPUT62), .B(n506), .ZN(n508) );
  INV_X1 U566 ( .A(G218GAT), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n508), .B(n507), .ZN(G1355GAT) );
  XNOR2_X1 U568 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n517) );
  NAND2_X1 U569 ( .A1(n603), .A2(n509), .ZN(n510) );
  XNOR2_X1 U570 ( .A(n510), .B(KEYINPUT76), .ZN(n511) );
  XNOR2_X1 U571 ( .A(n511), .B(KEYINPUT16), .ZN(n512) );
  NOR2_X1 U572 ( .A1(n513), .A2(n512), .ZN(n514) );
  XOR2_X1 U573 ( .A(KEYINPUT91), .B(n514), .Z(n532) );
  AND2_X1 U574 ( .A1(n515), .A2(n532), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n566), .A2(n524), .ZN(n516) );
  XNOR2_X1 U576 ( .A(n517), .B(n516), .ZN(G1324GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n519) );
  NAND2_X1 U578 ( .A1(n524), .A2(n546), .ZN(n518) );
  XNOR2_X1 U579 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U580 ( .A(G8GAT), .B(n520), .ZN(G1325GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT94), .B(KEYINPUT35), .Z(n522) );
  NAND2_X1 U582 ( .A1(n524), .A2(n551), .ZN(n521) );
  XNOR2_X1 U583 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U584 ( .A(G15GAT), .B(n523), .ZN(G1326GAT) );
  XOR2_X1 U585 ( .A(G22GAT), .B(KEYINPUT95), .Z(n526) );
  NAND2_X1 U586 ( .A1(n524), .A2(n541), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n526), .B(n525), .ZN(G1327GAT) );
  NAND2_X1 U588 ( .A1(n530), .A2(n566), .ZN(n529) );
  XNOR2_X1 U589 ( .A(G29GAT), .B(KEYINPUT99), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(KEYINPUT39), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n529), .B(n528), .ZN(G1328GAT) );
  NAND2_X1 U592 ( .A1(n530), .A2(n546), .ZN(n531) );
  XNOR2_X1 U593 ( .A(n531), .B(G36GAT), .ZN(G1329GAT) );
  AND2_X1 U594 ( .A1(n533), .A2(n532), .ZN(n542) );
  NAND2_X1 U595 ( .A1(n542), .A2(n566), .ZN(n537) );
  XOR2_X1 U596 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n535) );
  XNOR2_X1 U597 ( .A(G57GAT), .B(KEYINPUT105), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n537), .B(n536), .ZN(G1332GAT) );
  NAND2_X1 U600 ( .A1(n542), .A2(n546), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n538), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U602 ( .A1(n551), .A2(n542), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n539), .B(KEYINPUT106), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G71GAT), .B(n540), .ZN(G1334GAT) );
  XOR2_X1 U605 ( .A(G78GAT), .B(KEYINPUT43), .Z(n544) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(G1335GAT) );
  NAND2_X1 U608 ( .A1(n566), .A2(n548), .ZN(n545) );
  XNOR2_X1 U609 ( .A(G85GAT), .B(n545), .ZN(G1336GAT) );
  NAND2_X1 U610 ( .A1(n548), .A2(n546), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n547), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U612 ( .A1(n551), .A2(n548), .ZN(n549) );
  XNOR2_X1 U613 ( .A(n549), .B(G99GAT), .ZN(G1338GAT) );
  INV_X1 U614 ( .A(n550), .ZN(n583) );
  NAND2_X1 U615 ( .A1(n567), .A2(n551), .ZN(n552) );
  NOR2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n562) );
  NAND2_X1 U617 ( .A1(n583), .A2(n562), .ZN(n554) );
  XNOR2_X1 U618 ( .A(n554), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n557) );
  INV_X1 U620 ( .A(n555), .ZN(n585) );
  NAND2_X1 U621 ( .A1(n562), .A2(n585), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G120GAT), .B(n558), .ZN(G1341GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT50), .B(KEYINPUT113), .Z(n560) );
  NAND2_X1 U625 ( .A1(n562), .A2(n603), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G127GAT), .B(n561), .ZN(G1342GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n564) );
  NAND2_X1 U629 ( .A1(n562), .A2(n580), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G134GAT), .B(n565), .ZN(G1343GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U634 ( .A(KEYINPUT115), .B(n570), .Z(n581) );
  NAND2_X1 U635 ( .A1(n571), .A2(n581), .ZN(n572) );
  XNOR2_X1 U636 ( .A(n572), .B(KEYINPUT116), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G141GAT), .B(n573), .ZN(G1344GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n575) );
  NAND2_X1 U639 ( .A1(n581), .A2(n585), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n577) );
  XOR2_X1 U641 ( .A(G148GAT), .B(KEYINPUT53), .Z(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1345GAT) );
  NAND2_X1 U643 ( .A1(n603), .A2(n581), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n578), .B(KEYINPUT118), .ZN(n579) );
  XNOR2_X1 U645 ( .A(G155GAT), .B(n579), .ZN(G1346GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U648 ( .A1(n590), .A2(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G169GAT), .B(n584), .ZN(G1348GAT) );
  NAND2_X1 U650 ( .A1(n590), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(G176GAT), .B(KEYINPUT120), .Z(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n589) );
  XNOR2_X1 U653 ( .A(KEYINPUT57), .B(KEYINPUT56), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1349GAT) );
  XOR2_X1 U655 ( .A(G183GAT), .B(KEYINPUT121), .Z(n592) );
  NAND2_X1 U656 ( .A1(n590), .A2(n603), .ZN(n591) );
  XNOR2_X1 U657 ( .A(n592), .B(n591), .ZN(G1350GAT) );
  XOR2_X1 U658 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n594) );
  XNOR2_X1 U659 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n594), .B(n593), .ZN(n595) );
  XNOR2_X1 U661 ( .A(KEYINPUT125), .B(n595), .ZN(n598) );
  NOR2_X1 U662 ( .A1(n596), .A2(n599), .ZN(n597) );
  XNOR2_X1 U663 ( .A(n598), .B(n597), .ZN(G1352GAT) );
  XOR2_X1 U664 ( .A(G204GAT), .B(KEYINPUT61), .Z(n602) );
  INV_X1 U665 ( .A(n599), .ZN(n604) );
  NAND2_X1 U666 ( .A1(n600), .A2(n604), .ZN(n601) );
  XNOR2_X1 U667 ( .A(n602), .B(n601), .ZN(G1353GAT) );
  XOR2_X1 U668 ( .A(G211GAT), .B(KEYINPUT127), .Z(n606) );
  NAND2_X1 U669 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U670 ( .A(n606), .B(n605), .ZN(G1354GAT) );
endmodule

