//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n208), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT64), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n211), .B1(new_n221), .B2(KEYINPUT1), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n202), .A2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n239), .B(new_n245), .ZN(G351));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G274), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n248), .A2(new_n251), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(new_n254), .A2(G226), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G223), .A3(G1698), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1698), .B1(new_n258), .B2(new_n259), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G222), .ZN(new_n263));
  INV_X1    g0063(.A(G77), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n261), .B(new_n263), .C1(new_n264), .C2(new_n260), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n266));
  AOI211_X1 g0066(.A(new_n252), .B(new_n255), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G200), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT71), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n222), .B1(new_n208), .B2(new_n257), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT65), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G13), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n274), .A2(new_n223), .A3(G1), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n250), .A2(G20), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G50), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n223), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT8), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(new_n213), .B2(KEYINPUT66), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT66), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(KEYINPUT8), .A3(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n280), .B1(new_n281), .B2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n287), .A2(new_n273), .B1(new_n202), .B2(new_n275), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n278), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT9), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT70), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n289), .A2(new_n290), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(G190), .B2(new_n267), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n270), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  INV_X1    g0096(.A(G179), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n267), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n298), .B(new_n289), .C1(G169), .C2(new_n267), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n286), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n277), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n276), .A2(new_n303), .B1(new_n275), .B2(new_n286), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n271), .B(KEYINPUT65), .ZN(new_n305));
  AND2_X1   g0105(.A1(KEYINPUT3), .A2(G33), .ZN(new_n306));
  NOR2_X1   g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT7), .B1(new_n308), .B2(new_n223), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n223), .A4(new_n259), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(G68), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n213), .A2(new_n241), .ZN(new_n313));
  OAI21_X1  g0113(.A(G20), .B1(new_n313), .B2(new_n201), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n279), .A2(G159), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT16), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n305), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT78), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n310), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n308), .A2(KEYINPUT78), .A3(KEYINPUT7), .A4(new_n223), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n258), .A2(new_n223), .A3(new_n259), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n322), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G68), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n314), .A2(KEYINPUT16), .A3(new_n315), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT79), .B1(new_n320), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n241), .B1(new_n326), .B2(new_n310), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n319), .B1(new_n333), .B2(new_n316), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n273), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT79), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n329), .B1(new_n327), .B2(G68), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n304), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT17), .ZN(new_n340));
  INV_X1    g0140(.A(G223), .ZN(new_n341));
  INV_X1    g0141(.A(G1698), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n260), .B(new_n343), .C1(G226), .C2(new_n342), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G87), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n248), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n214), .A2(new_n253), .B1(new_n249), .B2(new_n251), .ZN(new_n347));
  OAI21_X1  g0147(.A(G200), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n345), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n266), .ZN(new_n350));
  INV_X1    g0150(.A(new_n347), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G190), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n348), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n339), .A2(new_n340), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n304), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n336), .B1(new_n335), .B2(new_n337), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n331), .A2(KEYINPUT79), .A3(new_n273), .A4(new_n334), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n354), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT17), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT18), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n346), .A2(new_n297), .A3(new_n347), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(G169), .B2(new_n352), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n363), .B1(new_n359), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n365), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n339), .A2(KEYINPUT18), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT80), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n366), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n359), .A2(new_n365), .ZN(new_n371));
  AOI21_X1  g0171(.A(KEYINPUT80), .B1(new_n371), .B2(KEYINPUT18), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n362), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n260), .A2(G232), .A3(new_n342), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n260), .A2(G238), .A3(G1698), .ZN(new_n375));
  INV_X1    g0175(.A(G107), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n374), .B(new_n375), .C1(new_n376), .C2(new_n260), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n248), .B1(new_n377), .B2(KEYINPUT67), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(KEYINPUT67), .B2(new_n377), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n252), .B1(G244), .B2(new_n254), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(KEYINPUT68), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT68), .B1(new_n379), .B2(new_n380), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n297), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n383), .ZN(new_n385));
  INV_X1    g0185(.A(G169), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n386), .A3(new_n381), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n276), .A2(G77), .A3(new_n277), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G20), .A2(G77), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT15), .B(G87), .ZN(new_n390));
  INV_X1    g0190(.A(new_n279), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT8), .B(G58), .ZN(new_n392));
  OAI221_X1 g0192(.A(new_n389), .B1(new_n390), .B2(new_n281), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(new_n273), .B1(new_n264), .B2(new_n275), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n384), .A2(new_n387), .A3(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(G190), .B1(new_n382), .B2(new_n383), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n385), .A2(G200), .A3(new_n381), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n395), .B(KEYINPUT69), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n300), .A2(new_n373), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n275), .A2(new_n241), .ZN(new_n403));
  XOR2_X1   g0203(.A(new_n403), .B(KEYINPUT12), .Z(new_n404));
  AOI21_X1  g0204(.A(new_n241), .B1(new_n250), .B2(G20), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n404), .B1(new_n276), .B2(new_n405), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n281), .A2(new_n264), .B1(new_n223), .B2(G68), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT74), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n407), .A2(new_n408), .B1(new_n202), .B2(new_n391), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n407), .A2(new_n408), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n273), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT11), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OR2_X1    g0213(.A1(new_n411), .A2(new_n412), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n406), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT75), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n406), .A2(new_n414), .A3(KEYINPUT75), .A4(new_n413), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI211_X1 g0219(.A(G226), .B(new_n342), .C1(new_n306), .C2(new_n307), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT72), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT72), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n260), .A2(new_n422), .A3(G226), .A4(new_n342), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g0224(.A(G232), .B(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G97), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n248), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G238), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n429), .A2(new_n253), .B1(new_n249), .B2(new_n251), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT13), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n430), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT13), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n425), .A2(new_n426), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n434), .B1(new_n423), .B2(new_n421), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n432), .B(new_n433), .C1(new_n435), .C2(new_n248), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n386), .B1(new_n431), .B2(new_n436), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT14), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n438), .A2(G179), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT77), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT76), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n422), .B1(new_n262), .B2(G226), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n420), .A2(KEYINPUT72), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n427), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n266), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n433), .B1(new_n447), .B2(new_n432), .ZN(new_n448));
  INV_X1    g0248(.A(new_n436), .ZN(new_n449));
  OAI21_X1  g0249(.A(G169), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n443), .B1(new_n450), .B2(KEYINPUT14), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n439), .A2(KEYINPUT76), .A3(new_n440), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n441), .B(new_n442), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n450), .A2(new_n443), .A3(KEYINPUT14), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT76), .B1(new_n439), .B2(new_n440), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n442), .B1(new_n457), .B2(new_n441), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n419), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n437), .A2(new_n353), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n460), .B(KEYINPUT73), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n417), .A2(new_n418), .B1(G200), .B2(new_n437), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n402), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n223), .B(G87), .C1(new_n306), .C2(new_n307), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT85), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT22), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n260), .A2(new_n223), .A3(G87), .A4(new_n469), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT23), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n223), .B2(G107), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n376), .A2(KEYINPUT23), .A3(G20), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n257), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n223), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n473), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(KEYINPUT86), .B1(new_n483), .B2(KEYINPUT24), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(KEYINPUT87), .A3(KEYINPUT24), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT87), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n481), .B1(new_n471), .B2(new_n472), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT24), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT86), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n487), .A2(new_n490), .A3(new_n488), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n484), .A2(new_n485), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n273), .ZN(new_n493));
  INV_X1    g0293(.A(new_n275), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n250), .A2(G33), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n305), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G107), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n275), .A2(new_n376), .ZN(new_n499));
  XOR2_X1   g0299(.A(new_n499), .B(KEYINPUT25), .Z(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(G257), .B(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n503));
  OAI211_X1 g0303(.A(G250), .B(new_n342), .C1(new_n306), .C2(new_n307), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G294), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g0306(.A(KEYINPUT5), .B(G41), .ZN(new_n507));
  INV_X1    g0307(.A(G45), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(G1), .ZN(new_n509));
  INV_X1    g0309(.A(new_n222), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n507), .A2(new_n509), .B1(new_n510), .B2(new_n247), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n506), .A2(new_n266), .B1(new_n511), .B2(G264), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n507), .A2(G274), .A3(new_n248), .A4(new_n509), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n268), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G190), .B2(new_n514), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n493), .A2(new_n502), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT6), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n215), .A2(new_n376), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(new_n205), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n376), .A2(KEYINPUT6), .A3(G97), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(G20), .B1(G77), .B2(new_n279), .ZN(new_n523));
  OAI21_X1  g0323(.A(G107), .B1(new_n309), .B2(new_n311), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n525), .A2(new_n273), .B1(new_n215), .B2(new_n275), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n497), .A2(G97), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(KEYINPUT5), .A2(G41), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(KEYINPUT5), .A2(G41), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n509), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n248), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n513), .B1(new_n533), .B2(new_n216), .ZN(new_n534));
  OAI211_X1 g0334(.A(G244), .B(new_n342), .C1(new_n306), .C2(new_n307), .ZN(new_n535));
  NOR2_X1   g0335(.A1(KEYINPUT81), .A2(KEYINPUT4), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(new_n536), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n260), .A2(G244), .A3(new_n342), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G283), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n260), .A2(G250), .A3(G1698), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n537), .A2(new_n539), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n534), .B1(new_n542), .B2(new_n266), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n386), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n297), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT82), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT82), .B1(new_n543), .B2(new_n297), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n528), .B(new_n545), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n544), .A2(G200), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n543), .A2(G190), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n551), .A2(new_n527), .A3(new_n526), .A4(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n517), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n250), .A2(G45), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n248), .A2(G250), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n248), .A2(G274), .A3(new_n509), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(G238), .B(new_n342), .C1(new_n306), .C2(new_n307), .ZN(new_n559));
  OAI211_X1 g0359(.A(G244), .B(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n560));
  INV_X1    g0360(.A(new_n479), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n558), .B1(new_n562), .B2(new_n266), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G179), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n563), .A2(new_n386), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT83), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n260), .A2(new_n223), .A3(G68), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT19), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n223), .B1(new_n426), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(G87), .B2(new_n206), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n281), .B2(new_n215), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n273), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n390), .A2(new_n275), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n574), .B(new_n575), .C1(new_n496), .C2(new_n390), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT83), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n564), .B(new_n577), .C1(new_n386), .C2(new_n563), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n567), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n575), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(G87), .B2(new_n497), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n562), .A2(new_n266), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(new_n556), .A3(new_n557), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G200), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n581), .B(new_n584), .C1(new_n353), .C2(new_n583), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n501), .B1(new_n492), .B2(new_n273), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n514), .A2(new_n386), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G179), .B2(new_n514), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n579), .B(new_n585), .C1(new_n586), .C2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n275), .A2(G116), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n496), .B2(G116), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n540), .B(new_n223), .C1(G33), .C2(new_n215), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT20), .ZN(new_n593));
  AOI22_X1  g0393(.A1(KEYINPUT84), .A2(new_n593), .B1(new_n478), .B2(G20), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n594), .A3(new_n271), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n593), .A2(KEYINPUT84), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n248), .A2(G274), .ZN(new_n599));
  INV_X1    g0399(.A(new_n531), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n555), .B1(new_n600), .B2(new_n529), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n511), .A2(G270), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(G264), .B(G1698), .C1(new_n306), .C2(new_n307), .ZN(new_n603));
  OAI211_X1 g0403(.A(G257), .B(new_n342), .C1(new_n306), .C2(new_n307), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n258), .A2(G303), .A3(new_n259), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n266), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n602), .A2(new_n607), .A3(G179), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n598), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT21), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n602), .A2(new_n607), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(G169), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n610), .B1(new_n598), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n612), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n614), .B(KEYINPUT21), .C1(new_n591), .C2(new_n597), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(G200), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n602), .A2(new_n607), .A3(G190), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n598), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n609), .A2(new_n613), .A3(new_n615), .A4(new_n618), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n554), .A2(new_n589), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n466), .A2(new_n620), .ZN(G372));
  OAI21_X1  g0421(.A(new_n564), .B1(new_n386), .B2(new_n563), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n576), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n585), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(new_n517), .A3(new_n550), .A4(new_n553), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n586), .A2(new_n588), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n609), .A2(new_n613), .A3(new_n615), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT88), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT88), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n627), .B2(new_n628), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n626), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n546), .B(new_n547), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n526), .A2(new_n527), .B1(new_n544), .B2(new_n386), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(new_n623), .A4(new_n585), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n623), .B1(new_n636), .B2(KEYINPUT26), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n579), .A2(new_n585), .ZN(new_n639));
  INV_X1    g0439(.A(new_n550), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n633), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n466), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n359), .A2(new_n360), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n340), .ZN(new_n646));
  AOI211_X1 g0446(.A(new_n356), .B(new_n354), .C1(new_n357), .C2(new_n358), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT17), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n396), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n463), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n649), .B1(new_n459), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n368), .A2(new_n366), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n296), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n655), .A2(new_n299), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n644), .A2(new_n656), .ZN(G369));
  INV_X1    g0457(.A(new_n628), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n250), .A2(new_n223), .A3(G13), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n598), .A2(new_n665), .ZN(new_n666));
  MUX2_X1   g0466(.A(new_n619), .B(new_n658), .S(new_n666), .Z(new_n667));
  INV_X1    g0467(.A(G330), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n627), .A2(new_n665), .ZN(new_n670));
  INV_X1    g0470(.A(new_n517), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n586), .A2(new_n665), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n671), .A2(new_n672), .B1(new_n586), .B2(new_n588), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n658), .A2(new_n664), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n675), .A2(new_n673), .A3(new_n670), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n670), .A3(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n209), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n250), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n681));
  INV_X1    g0481(.A(new_n226), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n680), .A2(new_n681), .B1(new_n682), .B2(new_n679), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT28), .Z(new_n684));
  NAND2_X1  g0484(.A1(new_n620), .A2(new_n665), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n583), .A2(new_n611), .A3(new_n297), .ZN(new_n686));
  INV_X1    g0486(.A(new_n514), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n686), .A2(new_n687), .A3(new_n543), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT90), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n608), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n563), .A2(new_n512), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n602), .A2(new_n607), .A3(KEYINPUT90), .A4(G179), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n690), .A2(new_n691), .A3(new_n543), .A4(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n688), .B1(new_n694), .B2(KEYINPUT30), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT30), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g0498(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n698), .A2(new_n664), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n693), .A2(KEYINPUT91), .A3(new_n696), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT91), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n695), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n664), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n685), .B(new_n701), .C1(KEYINPUT31), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT92), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(KEYINPUT92), .A3(G330), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n623), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n636), .B2(KEYINPUT26), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n639), .A2(new_n638), .A3(new_n640), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n715), .B(new_n716), .C1(new_n625), .C2(new_n629), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .A3(new_n665), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n664), .B1(new_n633), .B2(new_n642), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(KEYINPUT29), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n684), .B1(new_n722), .B2(G1), .ZN(G364));
  NOR2_X1   g0523(.A1(new_n274), .A2(G20), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT93), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G45), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n680), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n667), .A2(new_n730), .ZN(new_n731));
  NOR4_X1   g0531(.A1(new_n223), .A2(new_n353), .A3(new_n268), .A4(G179), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT96), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT96), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G303), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n223), .A2(new_n297), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n738), .A2(new_n268), .A3(G190), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT33), .B(G317), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(new_n353), .A3(new_n268), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n739), .A2(new_n740), .B1(new_n742), .B2(G311), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G179), .A2(G200), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(G20), .A3(new_n353), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI211_X1 g0547(.A(new_n260), .B(new_n744), .C1(G329), .C2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n737), .A2(G190), .A3(G200), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR4_X1   g0550(.A1(new_n223), .A2(new_n268), .A3(G179), .A4(G190), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n750), .A2(G326), .B1(G283), .B2(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n738), .A2(new_n353), .A3(G200), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n223), .B1(new_n745), .B2(G190), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n753), .A2(G322), .B1(G294), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n736), .A2(new_n748), .A3(new_n752), .A4(new_n756), .ZN(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(KEYINPUT97), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(KEYINPUT97), .ZN(new_n759));
  INV_X1    g0559(.A(new_n751), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n376), .ZN(new_n761));
  INV_X1    g0561(.A(new_n739), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n260), .B1(new_n754), .B2(new_n215), .C1(new_n762), .C2(new_n241), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT32), .ZN(new_n764));
  INV_X1    g0564(.A(G159), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n746), .A2(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n761), .B(new_n763), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n742), .A2(KEYINPUT95), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n742), .A2(KEYINPUT95), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G77), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n735), .A2(G87), .ZN(new_n773));
  INV_X1    g0573(.A(new_n753), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n774), .A2(new_n213), .B1(new_n764), .B2(new_n766), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G50), .B2(new_n750), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n767), .A2(new_n772), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n758), .A2(new_n759), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n222), .B1(G20), .B2(new_n386), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n730), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n678), .A2(new_n308), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n781), .A2(G355), .B1(new_n478), .B2(new_n678), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n308), .A2(new_n209), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(G45), .B2(new_n226), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n245), .A2(new_n508), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n782), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n727), .B1(new_n731), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n667), .B(new_n668), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(new_n790), .B2(new_n727), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT98), .ZN(G396));
  INV_X1    g0592(.A(new_n727), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n395), .A2(new_n664), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n400), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n396), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n650), .A2(new_n665), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g0598(.A(new_n719), .B(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n793), .B1(new_n713), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n713), .B2(new_n799), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n779), .A2(new_n728), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n727), .B1(new_n264), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n779), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n739), .A2(G150), .B1(new_n750), .B2(G137), .ZN(new_n805));
  INV_X1    g0605(.A(G143), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n806), .B2(new_n774), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(G159), .B2(new_n771), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n308), .B1(new_n747), .B2(G132), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n811), .B1(new_n213), .B2(new_n754), .C1(new_n241), .C2(new_n760), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G50), .B2(new_n735), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n809), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G303), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n749), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G294), .ZN(new_n817));
  OAI22_X1  g0617(.A1(new_n774), .A2(new_n817), .B1(new_n754), .B2(new_n215), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n816), .B(new_n818), .C1(G87), .C2(new_n751), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n735), .A2(G107), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n771), .A2(G116), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n308), .B1(new_n746), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(new_n739), .B2(G283), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n814), .A2(new_n825), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n803), .B1(new_n804), .B2(new_n826), .C1(new_n798), .C2(new_n729), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n801), .A2(new_n827), .ZN(G384));
  XNOR2_X1  g0628(.A(new_n522), .B(KEYINPUT99), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(KEYINPUT35), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n830), .A2(new_n478), .A3(new_n225), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n832), .A2(KEYINPUT100), .B1(KEYINPUT35), .B2(new_n829), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(KEYINPUT100), .B2(new_n832), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT36), .Z(new_n835));
  OAI211_X1 g0635(.A(new_n682), .B(G77), .C1(new_n213), .C2(new_n241), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n250), .B(G13), .C1(new_n836), .C2(new_n240), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT103), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n359), .A2(new_n369), .A3(new_n363), .A4(new_n365), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT18), .B1(new_n339), .B2(new_n367), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n368), .A2(new_n369), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n649), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n316), .B1(new_n327), .B2(G68), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n273), .B1(new_n845), .B2(KEYINPUT16), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT102), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(KEYINPUT102), .B(new_n273), .C1(new_n845), .C2(KEYINPUT16), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n848), .A2(new_n331), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n304), .ZN(new_n851));
  INV_X1    g0651(.A(new_n662), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n839), .B1(new_n844), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n645), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n851), .A2(new_n367), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI211_X1 g0657(.A(KEYINPUT104), .B(KEYINPUT37), .C1(new_n855), .C2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT104), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n357), .A2(new_n358), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n662), .B1(new_n860), .B2(new_n304), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n371), .A2(new_n861), .A3(new_n647), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n662), .B1(new_n850), .B2(new_n304), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(new_n647), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n863), .B1(new_n866), .B2(new_n856), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n858), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n373), .A2(KEYINPUT103), .A3(new_n865), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n854), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n854), .A2(KEYINPUT38), .A3(new_n868), .A4(new_n869), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n872), .A2(KEYINPUT39), .A3(new_n873), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n359), .B(new_n662), .C1(new_n362), .C2(new_n653), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n862), .B(KEYINPUT37), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n459), .A2(new_n664), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n874), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n653), .A2(new_n852), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n872), .A2(new_n873), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n417), .A2(new_n418), .A3(new_n664), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT101), .Z(new_n886));
  NAND3_X1  g0686(.A1(new_n459), .A2(new_n463), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n457), .A2(new_n441), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(KEYINPUT77), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(new_n453), .A3(new_n463), .ZN(new_n890));
  INV_X1    g0690(.A(new_n885), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n719), .A2(new_n798), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n893), .B1(new_n797), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n883), .B1(new_n884), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n882), .A2(new_n896), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n465), .A2(new_n720), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n656), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n897), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n796), .A2(new_n797), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n620), .A2(new_n665), .B1(new_n706), .B2(new_n699), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n707), .A2(KEYINPUT31), .ZN(new_n903));
  AOI221_X4 g0703(.A(new_n901), .B1(new_n902), .B2(new_n903), .C1(new_n887), .C2(new_n892), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n878), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT40), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n887), .A2(new_n892), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT40), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n902), .A2(new_n903), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n907), .A2(new_n908), .A3(new_n798), .A4(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n884), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n465), .B1(new_n903), .B2(new_n902), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n668), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n914), .B2(new_n913), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n900), .A2(new_n916), .B1(new_n250), .B2(new_n725), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT105), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n900), .A2(new_n916), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n917), .B2(new_n918), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n838), .B1(new_n919), .B2(new_n921), .ZN(G367));
  NOR2_X1   g0722(.A1(new_n581), .A2(new_n665), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n624), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT106), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n714), .A2(new_n923), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n624), .A2(KEYINPUT106), .A3(new_n924), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n930), .A2(KEYINPUT107), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(KEYINPUT107), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n730), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n749), .A2(new_n806), .B1(new_n754), .B2(new_n241), .ZN(new_n935));
  INV_X1    g0735(.A(G137), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n762), .A2(new_n765), .B1(new_n936), .B2(new_n746), .ZN(new_n937));
  AOI211_X1 g0737(.A(new_n935), .B(new_n937), .C1(G150), .C2(new_n753), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n771), .A2(G50), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n308), .B1(new_n751), .B2(G77), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT109), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n735), .A2(G58), .B1(KEYINPUT109), .B2(new_n940), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n938), .A2(new_n939), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT46), .B1(new_n735), .B2(G116), .ZN(new_n944));
  XNOR2_X1  g0744(.A(KEYINPUT108), .B(G317), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n260), .B1(new_n747), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(G283), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n946), .B1(new_n817), .B2(new_n762), .C1(new_n770), .C2(new_n947), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n774), .A2(new_n815), .B1(new_n754), .B2(new_n376), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n760), .A2(new_n215), .B1(new_n822), .B2(new_n749), .ZN(new_n950));
  OR4_X1    g0750(.A1(new_n944), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n735), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT46), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n952), .A2(new_n953), .A3(new_n478), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n943), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT47), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n779), .ZN(new_n957));
  INV_X1    g0757(.A(new_n784), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n780), .B1(new_n209), .B2(new_n390), .C1(new_n958), .C2(new_n235), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n934), .A2(new_n793), .A3(new_n957), .A4(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT43), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n933), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n676), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n640), .A2(new_n664), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n528), .A2(new_n664), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n550), .A2(new_n553), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n627), .A2(new_n553), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n664), .B1(new_n972), .B2(new_n550), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n933), .A2(new_n962), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n963), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n968), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n674), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n974), .A2(new_n962), .A3(new_n933), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n980), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n982), .A2(new_n976), .B1(new_n674), .B2(new_n978), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n726), .A2(G1), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n676), .A2(new_n670), .A3(new_n968), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT45), .Z(new_n988));
  AOI21_X1  g0788(.A(new_n968), .B1(new_n676), .B2(new_n670), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT44), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n988), .A2(new_n674), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n674), .B1(new_n988), .B2(new_n990), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n675), .B1(new_n673), .B2(new_n670), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n964), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(new_n669), .Z(new_n996));
  AOI21_X1  g0796(.A(new_n721), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n679), .B(KEYINPUT41), .Z(new_n998));
  OAI21_X1  g0798(.A(new_n986), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n961), .B1(new_n984), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(G387));
  NAND2_X1  g0801(.A1(new_n996), .A2(new_n985), .ZN(new_n1002));
  AOI211_X1 g0802(.A(G20), .B(new_n729), .C1(new_n673), .C2(new_n670), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n750), .A2(G322), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n753), .A2(new_n945), .B1(new_n739), .B2(G311), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1004), .B(new_n1005), .C1(new_n770), .C2(new_n815), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT48), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n735), .A2(G294), .B1(G283), .B2(new_n755), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT49), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n760), .A2(new_n478), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n260), .B(new_n1015), .C1(G326), .C2(new_n747), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n735), .A2(G77), .ZN(new_n1018));
  INV_X1    g0818(.A(G150), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n746), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(KEYINPUT110), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(KEYINPUT110), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n774), .A2(new_n202), .B1(new_n754), .B2(new_n390), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n301), .B2(new_n739), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n260), .B1(new_n741), .B2(new_n241), .C1(new_n760), .C2(new_n215), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n749), .A2(KEYINPUT111), .A3(new_n765), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT111), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n750), .B2(G159), .ZN(new_n1028));
  NOR3_X1   g0828(.A1(new_n1025), .A2(new_n1026), .A3(new_n1028), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n804), .B1(new_n1017), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n681), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1032), .A2(new_n781), .B1(new_n376), .B2(new_n678), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n232), .A2(new_n508), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n392), .A2(G50), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT50), .Z(new_n1036));
  OAI211_X1 g0836(.A(new_n681), .B(new_n508), .C1(new_n241), .C2(new_n264), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n784), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1033), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n727), .B(new_n1031), .C1(new_n780), .C2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT112), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n722), .A2(new_n996), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n713), .A2(new_n996), .A3(new_n720), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n679), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1002), .B1(new_n1003), .B2(new_n1041), .C1(new_n1042), .C2(new_n1044), .ZN(G393));
  NAND2_X1  g0845(.A1(new_n993), .A2(new_n985), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n978), .A2(new_n730), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n774), .A2(new_n765), .B1(new_n749), .B2(new_n1019), .ZN(new_n1048));
  XOR2_X1   g0848(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n735), .A2(G68), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n260), .B1(new_n746), .B2(new_n806), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n739), .B2(G50), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n754), .A2(new_n264), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(G87), .B2(new_n751), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1054), .B(new_n1056), .C1(new_n770), .C2(new_n392), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n735), .A2(G283), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n260), .B1(new_n742), .B2(G294), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n739), .A2(G303), .B1(G322), .B2(new_n747), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n761), .B1(G116), .B2(new_n755), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n753), .A2(G311), .B1(new_n750), .B2(G317), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT52), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n1052), .A2(new_n1057), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n779), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n780), .B1(new_n215), .B2(new_n209), .C1(new_n958), .C2(new_n239), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1047), .A2(new_n793), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1046), .A2(new_n1068), .ZN(new_n1069));
  NOR3_X1   g0869(.A1(new_n1043), .A2(new_n991), .A3(new_n992), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n1070), .A2(G41), .A3(new_n678), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n993), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n1043), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1069), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(G390));
  NOR2_X1   g0875(.A1(new_n893), .A2(new_n901), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n668), .B1(new_n902), .B2(new_n903), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n717), .A2(new_n796), .A3(new_n665), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n797), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n881), .B1(new_n907), .B2(new_n1081), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n878), .A2(KEYINPUT114), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT114), .B1(new_n878), .B2(new_n1082), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n881), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n894), .A2(new_n797), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n907), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n874), .A2(new_n880), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1079), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n874), .A2(new_n880), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1088), .A2(new_n1086), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n878), .A2(new_n1082), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT114), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n878), .A2(new_n1082), .A3(KEYINPUT114), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n901), .B1(new_n711), .B2(new_n712), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n907), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1093), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1090), .A2(new_n1101), .A3(new_n985), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1091), .A2(new_n728), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n802), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n793), .B1(new_n301), .B2(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n774), .A2(new_n478), .B1(new_n749), .B2(new_n947), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1055), .B(new_n1106), .C1(G68), .C2(new_n751), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n771), .A2(G97), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n308), .B1(new_n746), .B2(new_n817), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n739), .B2(G107), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1107), .A2(new_n773), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(KEYINPUT53), .B1(new_n952), .B2(new_n1019), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n753), .A2(G132), .B1(G50), .B2(new_n751), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n750), .A2(G128), .B1(new_n755), .B2(G159), .ZN(new_n1114));
  INV_X1    g0914(.A(G125), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n260), .B1(new_n746), .B2(new_n1115), .C1(new_n762), .C2(new_n936), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT54), .B(G143), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1116), .B1(new_n771), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .A4(new_n1119), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n952), .A2(KEYINPUT53), .A3(new_n1019), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1111), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1105), .B1(new_n1122), .B2(new_n779), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1103), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1078), .B1(new_n1099), .B2(new_n907), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1077), .A2(new_n798), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1081), .B1(new_n1126), .B2(new_n893), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1125), .A2(new_n1087), .B1(new_n1100), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n466), .A2(new_n1077), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n898), .A3(new_n656), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT115), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1090), .A2(new_n1101), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1101), .B(new_n1090), .C1(new_n1131), .C2(KEYINPUT115), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n679), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1102), .B(new_n1124), .C1(new_n1136), .C2(new_n1138), .ZN(G378));
  NAND2_X1  g0939(.A1(new_n289), .A2(new_n852), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1140), .B(KEYINPUT55), .Z(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n296), .A2(new_n299), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  XOR2_X1   g0944(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1142), .B1(new_n296), .B2(new_n299), .ZN(new_n1147));
  OR3_X1    g0947(.A1(new_n1144), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n913), .B2(G330), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n908), .B1(new_n878), .B2(new_n904), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n910), .B1(new_n873), .B2(new_n872), .ZN(new_n1153));
  OAI211_X1 g0953(.A(G330), .B(new_n1150), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n897), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1150), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n668), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n897), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n1154), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1156), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1125), .A2(new_n1087), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1100), .A2(new_n1127), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1090), .A2(new_n1165), .A3(new_n1101), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1130), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1162), .A2(new_n1168), .A3(KEYINPUT57), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n897), .A2(KEYINPUT118), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT118), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n882), .A2(new_n896), .A3(new_n1171), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(new_n1151), .C2(new_n1155), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1173), .A2(new_n1161), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1169), .B(new_n679), .C1(KEYINPUT57), .C2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n793), .B1(G50), .B2(new_n1104), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1150), .A2(new_n729), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1178));
  INV_X1    g0978(.A(G41), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n308), .B2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n308), .B(new_n1179), .C1(new_n746), .C2(new_n947), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n741), .A2(new_n390), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(G97), .C2(new_n739), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n755), .A2(G68), .B1(new_n751), .B2(G58), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n753), .A2(G107), .B1(new_n750), .B2(G116), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1018), .A2(new_n1183), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT58), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1180), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n739), .A2(G132), .B1(new_n742), .B2(G137), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT116), .ZN(new_n1190));
  INV_X1    g0990(.A(G128), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n774), .A2(new_n1191), .B1(new_n749), .B2(new_n1115), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G150), .B2(new_n755), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1190), .B(new_n1193), .C1(new_n952), .C2(new_n1117), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n751), .A2(G159), .ZN(new_n1196));
  AOI211_X1 g0996(.A(G33), .B(G41), .C1(new_n747), .C2(G124), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1188), .B1(new_n1187), .B2(new_n1186), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n1176), .B(new_n1177), .C1(new_n779), .C2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1161), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1201), .B1(new_n1204), .B2(new_n985), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1175), .A2(new_n1205), .ZN(G375));
  INV_X1    g1006(.A(new_n998), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1132), .A2(new_n1207), .A3(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n893), .A2(new_n728), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n793), .B1(G68), .B2(new_n1104), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n762), .A2(new_n1117), .B1(new_n1191), .B2(new_n746), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n308), .B(new_n1212), .C1(G150), .C2(new_n742), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n735), .A2(G159), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n755), .A2(G50), .B1(new_n751), .B2(G58), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n753), .A2(G137), .B1(new_n750), .B2(G132), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n760), .A2(new_n264), .B1(new_n390), .B2(new_n754), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n770), .A2(new_n376), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n774), .A2(new_n947), .B1(new_n749), .B2(new_n817), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n308), .B1(new_n746), .B2(new_n815), .C1(new_n762), .C2(new_n478), .ZN(new_n1221));
  OR4_X1    g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n952), .A2(new_n215), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1217), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1211), .B1(new_n1224), .B2(new_n779), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1165), .A2(new_n985), .B1(new_n1210), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1209), .A2(new_n1226), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT119), .ZN(G381));
  OR2_X1    g1028(.A1(G393), .A2(G396), .ZN(new_n1229));
  INV_X1    g1029(.A(G384), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1074), .A2(new_n1230), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(G381), .A2(G387), .A3(new_n1229), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1102), .A2(new_n1124), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1138), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n1234), .B2(new_n1135), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1232), .A2(new_n1235), .A3(new_n1175), .A4(new_n1205), .ZN(G407));
  NAND2_X1  g1036(.A1(new_n663), .A2(G213), .ZN(new_n1237));
  OR3_X1    g1037(.A1(G375), .A2(G378), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G407), .A2(G213), .A3(new_n1238), .ZN(G409));
  INV_X1    g1039(.A(KEYINPUT125), .ZN(new_n1240));
  OAI21_X1  g1040(.A(G390), .B1(new_n1000), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n981), .A2(new_n983), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1207), .B1(new_n1070), .B2(new_n721), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n1243), .B2(new_n986), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1074), .B(KEYINPUT125), .C1(new_n1244), .C2(new_n961), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(G393), .B(G396), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1241), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT126), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT126), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1241), .A2(new_n1245), .A3(new_n1249), .A4(new_n1246), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  OR2_X1    g1051(.A1(new_n1246), .A2(KEYINPUT123), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G390), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1074), .A2(KEYINPUT124), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n1000), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(G387), .A2(new_n1253), .A3(G390), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1246), .A2(KEYINPUT123), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1252), .A2(new_n1256), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1251), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT60), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1208), .B1(new_n1131), .B2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1128), .A2(KEYINPUT60), .A3(new_n1130), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n679), .A3(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1264), .A2(new_n1226), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(G384), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n663), .A2(G213), .A3(G2897), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(new_n1266), .B(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1204), .A2(new_n1207), .A3(new_n1168), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT120), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT120), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1174), .A2(new_n1271), .A3(new_n1207), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1201), .B1(new_n1162), .B2(new_n985), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1235), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(G378), .A2(new_n1175), .A3(new_n1205), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1237), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT61), .B1(new_n1268), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(KEYINPUT62), .B1(new_n1278), .B2(new_n1266), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1277), .A2(KEYINPUT121), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT121), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1275), .A2(new_n1283), .A3(new_n1276), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1265), .B(new_n1230), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1282), .A2(new_n1237), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1286), .A2(KEYINPUT62), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1260), .B1(new_n1281), .B2(new_n1287), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1277), .A2(KEYINPUT63), .A3(new_n1237), .A4(new_n1285), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT61), .B1(new_n1251), .B2(new_n1259), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1292), .B2(new_n1286), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1284), .A2(new_n1237), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1283), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1295));
  OAI21_X1  g1095(.A(KEYINPUT122), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT122), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1282), .A2(new_n1297), .A3(new_n1237), .A4(new_n1284), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1268), .A3(new_n1298), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1293), .A2(KEYINPUT127), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT127), .B1(new_n1293), .B2(new_n1299), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1288), .B1(new_n1300), .B2(new_n1301), .ZN(G405));
  NAND2_X1  g1102(.A1(G375), .A2(new_n1235), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1276), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1304), .B(new_n1285), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(new_n1305), .B(new_n1260), .ZN(G402));
endmodule


