//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XOR2_X1   g002(.A(G197gat), .B(G204gat), .Z(new_n204));
  INV_X1    g003(.A(KEYINPUT75), .ZN(new_n205));
  INV_X1    g004(.A(G211gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT74), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n206), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n205), .B1(new_n211), .B2(KEYINPUT22), .ZN(new_n212));
  AND2_X1   g011(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT74), .A2(G218gat), .ZN(new_n214));
  OAI21_X1  g013(.A(G211gat), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT22), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(KEYINPUT75), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n204), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n203), .B1(new_n218), .B2(KEYINPUT76), .ZN(new_n219));
  INV_X1    g018(.A(new_n204), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n215), .A2(KEYINPUT75), .A3(new_n216), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT75), .B1(new_n215), .B2(new_n216), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT76), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(new_n202), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G226gat), .A2(G233gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G169gat), .ZN(new_n232));
  INV_X1    g031(.A(G176gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n233), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(KEYINPUT26), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(new_n232), .A3(new_n233), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT26), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n231), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n229), .A2(KEYINPUT27), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT27), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G183gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n245), .A3(new_n230), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT68), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT28), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n246), .A2(KEYINPUT69), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT28), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT69), .B1(new_n246), .B2(KEYINPUT68), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n242), .B(new_n250), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n229), .A2(new_n230), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT66), .B(KEYINPUT24), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(new_n231), .ZN(new_n257));
  NAND3_X1  g056(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n238), .A2(KEYINPUT23), .A3(new_n240), .ZN(new_n262));
  OAI21_X1  g061(.A(KEYINPUT23), .B1(new_n232), .B2(new_n233), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n235), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT25), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT25), .B1(new_n263), .B2(new_n235), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n258), .B(new_n255), .C1(new_n231), .C2(KEYINPUT24), .ZN(new_n268));
  OR2_X1    g067(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n269), .A2(KEYINPUT23), .A3(new_n233), .A4(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n267), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n254), .A2(new_n266), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n228), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n264), .B(new_n262), .C1(new_n257), .C2(new_n260), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n272), .B1(new_n277), .B2(KEYINPUT25), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n227), .B1(new_n278), .B2(new_n254), .ZN(new_n279));
  OAI211_X1 g078(.A(KEYINPUT77), .B(new_n226), .C1(new_n276), .C2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(new_n228), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT29), .B1(new_n278), .B2(new_n254), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(new_n228), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT77), .B1(new_n284), .B2(new_n226), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n226), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT78), .B1(new_n283), .B2(new_n228), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n274), .A2(new_n275), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n279), .B1(new_n289), .B2(new_n227), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n287), .B(new_n288), .C1(new_n290), .C2(KEYINPUT78), .ZN(new_n291));
  XNOR2_X1  g090(.A(G8gat), .B(G36gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(G64gat), .B(G92gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  NAND4_X1  g093(.A1(new_n286), .A2(KEYINPUT30), .A3(new_n291), .A4(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT77), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(new_n290), .B2(new_n287), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n291), .A2(new_n297), .A3(new_n280), .A4(new_n294), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT30), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n291), .A2(new_n280), .A3(new_n297), .ZN(new_n301));
  INV_X1    g100(.A(new_n294), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n295), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT87), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT87), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n295), .A2(new_n300), .A3(new_n306), .A4(new_n303), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G127gat), .B(G134gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G113gat), .B(G120gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(KEYINPUT1), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n311), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(new_n309), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G141gat), .B(G148gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT81), .ZN(new_n318));
  NAND2_X1  g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n318), .B1(new_n319), .B2(KEYINPUT2), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n318), .A3(KEYINPUT2), .ZN(new_n322));
  INV_X1    g121(.A(new_n319), .ZN(new_n323));
  NOR2_X1   g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT80), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n324), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT80), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(new_n327), .A3(new_n319), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n321), .A2(new_n322), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n317), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n319), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n319), .A2(KEYINPUT2), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n316), .A2(new_n329), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n320), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n330), .A2(new_n335), .A3(new_n322), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n328), .A2(new_n325), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n317), .B1(new_n319), .B2(new_n326), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n332), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n338), .A2(new_n340), .B1(new_n315), .B2(new_n312), .ZN(new_n341));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n334), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(KEYINPUT88), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n338), .A2(new_n340), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n346), .A2(new_n347), .A3(new_n316), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n329), .A2(new_n333), .ZN(new_n349));
  INV_X1    g148(.A(new_n316), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT4), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT3), .B1(new_n329), .B2(new_n333), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n340), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n355), .A3(new_n316), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n343), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n345), .A2(KEYINPUT39), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT0), .ZN(new_n361));
  XNOR2_X1  g160(.A(G57gat), .B(G85gat), .ZN(new_n362));
  XOR2_X1   g161(.A(new_n361), .B(new_n362), .Z(new_n363));
  OAI211_X1 g162(.A(new_n359), .B(new_n363), .C1(KEYINPUT39), .C2(new_n358), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT40), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n352), .A2(KEYINPUT5), .A3(new_n342), .A4(new_n356), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n343), .B1(new_n334), .B2(new_n341), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT5), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n347), .B1(new_n346), .B2(new_n316), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n349), .A2(new_n350), .A3(KEYINPUT4), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n356), .A2(new_n370), .A3(new_n371), .A4(new_n342), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n363), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n367), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(new_n364), .B2(new_n365), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n308), .A2(new_n366), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n219), .A2(new_n225), .A3(new_n275), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT83), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n219), .A2(new_n225), .A3(new_n381), .A4(new_n275), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(new_n354), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n346), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n355), .A2(new_n275), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n226), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(G228gat), .A3(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G22gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(G228gat), .A2(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n386), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n223), .A2(new_n202), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n218), .A2(new_n203), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(new_n275), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n349), .B1(new_n395), .B2(new_n354), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n391), .B1(new_n392), .B2(new_n396), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n389), .A2(KEYINPUT84), .A3(new_n390), .A4(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT3), .B1(new_n379), .B2(KEYINPUT83), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n349), .B1(new_n399), .B2(new_n382), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n390), .B(new_n397), .C1(new_n400), .C2(new_n387), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT84), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n397), .B1(new_n400), .B2(new_n387), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(G22gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n398), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G78gat), .B(G106gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(KEYINPUT31), .B(G50gat), .ZN(new_n408));
  XOR2_X1   g207(.A(new_n407), .B(new_n408), .Z(new_n409));
  NAND2_X1  g208(.A1(new_n406), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT85), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n389), .A2(KEYINPUT86), .A3(new_n390), .A4(new_n397), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n401), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n409), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n414), .A2(new_n416), .A3(new_n417), .A4(new_n405), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n411), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT90), .ZN(new_n420));
  XOR2_X1   g219(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n421));
  NAND4_X1  g220(.A1(new_n286), .A2(new_n420), .A3(new_n291), .A4(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n291), .A2(new_n297), .A3(new_n280), .A4(new_n421), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT90), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n301), .A2(KEYINPUT37), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n302), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT38), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n367), .A2(new_n373), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n363), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n375), .A3(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n367), .A2(new_n373), .A3(KEYINPUT6), .A4(new_n374), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n298), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n294), .B1(new_n422), .B2(new_n424), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n226), .B(new_n288), .C1(new_n290), .C2(KEYINPUT78), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT37), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n437), .B1(new_n284), .B2(new_n287), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT38), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n428), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n378), .A2(new_n419), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT79), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n295), .A2(new_n444), .A3(new_n303), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n432), .A2(new_n433), .B1(new_n298), .B2(new_n299), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n444), .B1(new_n295), .B2(new_n303), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n443), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n295), .A2(new_n303), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT79), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n451), .A2(KEYINPUT82), .A3(new_n445), .A4(new_n446), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n406), .A2(new_n412), .A3(new_n409), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n412), .B1(new_n406), .B2(new_n409), .ZN(new_n455));
  INV_X1    g254(.A(new_n418), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT34), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n274), .A2(KEYINPUT70), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT70), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n278), .A2(new_n461), .A3(new_n254), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n316), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n274), .A2(KEYINPUT70), .A3(new_n350), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(G227gat), .ZN(new_n466));
  INV_X1    g265(.A(G233gat), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n459), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  AOI211_X1 g269(.A(KEYINPUT34), .B(new_n468), .C1(new_n463), .C2(new_n464), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n463), .A2(new_n468), .A3(new_n464), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT32), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT33), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  XOR2_X1   g275(.A(G15gat), .B(G43gat), .Z(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT71), .ZN(new_n478));
  XOR2_X1   g277(.A(G71gat), .B(G99gat), .Z(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(KEYINPUT72), .ZN(new_n480));
  XOR2_X1   g279(.A(new_n478), .B(new_n480), .Z(new_n481));
  NAND3_X1  g280(.A1(new_n474), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n481), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n473), .B(KEYINPUT32), .C1(new_n475), .C2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n472), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n472), .B1(new_n482), .B2(new_n484), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n482), .A2(new_n484), .ZN(new_n492));
  INV_X1    g291(.A(new_n472), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(KEYINPUT73), .A3(new_n485), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT73), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n487), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n491), .B1(new_n499), .B2(new_n490), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n442), .A2(new_n458), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n419), .A2(new_n449), .A3(new_n452), .A4(new_n498), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n455), .A2(new_n456), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n308), .B1(new_n503), .B2(new_n413), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n432), .A2(new_n433), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n489), .A2(KEYINPUT35), .A3(new_n506), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n502), .A2(KEYINPUT35), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n390), .A2(G15gat), .ZN(new_n510));
  INV_X1    g309(.A(G15gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(G22gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT16), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n510), .B(new_n512), .C1(new_n513), .C2(G1gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(G1gat), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G8gat), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT95), .B1(new_n515), .B2(G1gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  OAI221_X1 g318(.A(new_n514), .B1(KEYINPUT95), .B2(G8gat), .C1(G1gat), .C2(new_n515), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT14), .ZN(new_n524));
  INV_X1    g323(.A(G29gat), .ZN(new_n525));
  INV_X1    g324(.A(G36gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n527), .A2(KEYINPUT93), .ZN(new_n528));
  NOR3_X1   g327(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT93), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n523), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G29gat), .A2(G36gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT15), .ZN(new_n534));
  XNOR2_X1  g333(.A(G43gat), .B(G50gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n535), .A2(new_n536), .A3(new_n534), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n532), .B(new_n533), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n535), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(new_n534), .ZN(new_n542));
  INV_X1    g341(.A(new_n523), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n533), .B1(new_n543), .B2(new_n529), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT96), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n522), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n527), .A2(KEYINPUT93), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n529), .A2(new_n530), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n551), .A2(new_n523), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n541), .A2(KEYINPUT92), .A3(KEYINPUT15), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n537), .ZN(new_n554));
  AOI22_X1  g353(.A1(new_n552), .A2(new_n554), .B1(new_n544), .B2(new_n542), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT96), .B1(new_n555), .B2(new_n521), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n540), .A2(KEYINPUT17), .A3(new_n545), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT94), .B(KEYINPUT17), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n559), .B(new_n521), .C1(new_n555), .C2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT97), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT99), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT18), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n557), .A2(KEYINPUT97), .A3(new_n558), .A4(new_n561), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n555), .A2(new_n521), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n547), .B1(new_n522), .B2(new_n546), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n555), .A2(new_n521), .A3(KEYINPUT96), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT98), .B(KEYINPUT13), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(new_n558), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n557), .A2(KEYINPUT18), .A3(new_n558), .A4(new_n561), .ZN(new_n577));
  XNOR2_X1  g376(.A(G113gat), .B(G141gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G169gat), .B(G197gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT12), .Z(new_n583));
  AND3_X1   g382(.A1(new_n576), .A2(new_n577), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT18), .B1(new_n562), .B2(new_n563), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n565), .B1(new_n586), .B2(new_n567), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n576), .A2(new_n577), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n588), .B1(new_n567), .B2(new_n586), .ZN(new_n589));
  OAI22_X1  g388(.A1(new_n585), .A2(new_n587), .B1(new_n589), .B2(new_n583), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT103), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n592));
  INV_X1    g391(.A(G155gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT101), .ZN(new_n599));
  OR2_X1    g398(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n600), .A2(G64gat), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G64gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(G57gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G71gat), .B(G78gat), .Z(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n604), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n603), .A2(G57gat), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT9), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(new_n606), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(G127gat), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n613), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT21), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n521), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n617), .B(G127gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(new_n624), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n597), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n621), .A2(new_n625), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n624), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n596), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G85gat), .ZN(new_n635));
  INV_X1    g434(.A(G92gat), .ZN(new_n636));
  OAI21_X1  g435(.A(KEYINPUT7), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT7), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(G85gat), .A3(G92gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G99gat), .B(G106gat), .Z(new_n641));
  NAND2_X1  g440(.A1(G99gat), .A2(G106gat), .ZN(new_n642));
  AOI22_X1  g441(.A1(KEYINPUT8), .A2(new_n642), .B1(new_n635), .B2(new_n636), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n640), .A2(new_n641), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n641), .B1(new_n640), .B2(new_n643), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n559), .B(new_n646), .C1(new_n555), .C2(new_n560), .ZN(new_n647));
  INV_X1    g446(.A(new_n646), .ZN(new_n648));
  INV_X1    g447(.A(G232gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n467), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n546), .A2(new_n648), .B1(KEYINPUT41), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G190gat), .B(G218gat), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G134gat), .B(G162gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(new_n654), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n650), .A2(KEYINPUT41), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  INV_X1    g461(.A(new_n658), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n652), .A2(new_n656), .A3(new_n663), .ZN(new_n664));
  AND3_X1   g463(.A1(new_n659), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n659), .B2(new_n664), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n591), .B1(new_n634), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n667), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n633), .A2(new_n669), .A3(KEYINPUT103), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT10), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n640), .A2(new_n643), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n641), .A2(KEYINPUT105), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n622), .A2(new_n674), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n613), .A2(new_n646), .A3(KEYINPUT104), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT104), .B1(new_n613), .B2(new_n646), .ZN(new_n677));
  OAI211_X1 g476(.A(new_n671), .B(new_n675), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n622), .A2(new_n648), .A3(KEYINPUT10), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(G230gat), .A2(G233gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT106), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n685));
  INV_X1    g484(.A(new_n681), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(G120gat), .B(G148gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(G176gat), .B(G204gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n689), .B(new_n690), .Z(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n686), .B1(new_n678), .B2(new_n679), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n687), .A3(new_n691), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AND4_X1   g497(.A1(new_n590), .A2(new_n668), .A3(new_n670), .A4(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n509), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n506), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g502(.A(new_n517), .B1(new_n701), .B2(new_n308), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n305), .A2(new_n307), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT16), .B(G8gat), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n700), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT42), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(KEYINPUT42), .B2(new_n707), .ZN(G1325gat));
  NOR2_X1   g508(.A1(new_n488), .A2(KEYINPUT36), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(KEYINPUT36), .B2(new_n498), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT107), .ZN(new_n712));
  OAI21_X1  g511(.A(G15gat), .B1(new_n700), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n488), .A2(new_n511), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n713), .B1(new_n700), .B2(new_n714), .ZN(G1326gat));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n419), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT43), .B(G22gat), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1327gat));
  OAI21_X1  g517(.A(new_n667), .B1(new_n501), .B2(new_n508), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n576), .A2(new_n577), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n583), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n568), .A2(new_n584), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(KEYINPUT99), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n726), .A2(new_n633), .A3(new_n697), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n720), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n505), .A2(G29gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(KEYINPUT45), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT44), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n719), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g532(.A(KEYINPUT44), .B(new_n667), .C1(new_n501), .C2(new_n508), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n727), .B(KEYINPUT108), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G29gat), .B1(new_n736), .B2(new_n505), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n738));
  INV_X1    g537(.A(new_n730), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n728), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n731), .A2(new_n737), .A3(new_n740), .ZN(G1328gat));
  XNOR2_X1  g540(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n705), .A2(G36gat), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n728), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G36gat), .B1(new_n736), .B2(new_n705), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n742), .B1(new_n728), .B2(new_n744), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(G1329gat));
  NOR3_X1   g547(.A1(new_n728), .A2(G43gat), .A3(new_n489), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G43gat), .B1(new_n736), .B2(new_n500), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n750), .A2(KEYINPUT47), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n500), .B(KEYINPUT107), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n733), .A2(new_n753), .A3(new_n734), .A4(new_n735), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n754), .A2(new_n755), .A3(G43gat), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n755), .B1(new_n754), .B2(G43gat), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n756), .A2(new_n757), .A3(new_n749), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n752), .B1(new_n758), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g558(.A1(new_n457), .A2(G50gat), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n736), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(G50gat), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n728), .B2(new_n419), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT48), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT48), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n766), .A3(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1331gat));
  AND4_X1   g567(.A1(new_n726), .A2(new_n668), .A3(new_n670), .A4(new_n697), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n509), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n506), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n600), .A2(new_n601), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1332gat));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n308), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT49), .B(G64gat), .Z(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(G1333gat));
  NAND3_X1  g576(.A1(new_n770), .A2(G71gat), .A3(new_n753), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n488), .B(KEYINPUT111), .Z(new_n780));
  AOI21_X1  g579(.A(G71gat), .B1(new_n770), .B2(new_n780), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n779), .A2(KEYINPUT50), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT50), .B1(new_n779), .B2(new_n781), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(G1334gat));
  NAND2_X1  g583(.A1(new_n770), .A2(new_n457), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g585(.A1(new_n633), .A2(new_n590), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n509), .A2(KEYINPUT51), .A3(new_n667), .A4(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  INV_X1    g588(.A(new_n787), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n719), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OAI211_X1 g592(.A(KEYINPUT112), .B(new_n789), .C1(new_n719), .C2(new_n790), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n698), .A2(new_n505), .A3(G85gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n790), .A2(new_n698), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n733), .A2(new_n734), .A3(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(G85gat), .B1(new_n798), .B2(new_n505), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n796), .A2(KEYINPUT113), .A3(new_n799), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(G1336gat));
  NOR3_X1   g603(.A1(new_n705), .A2(G92gat), .A3(new_n698), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n793), .A2(new_n794), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n733), .A2(new_n308), .A3(new_n734), .A4(new_n797), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G92gat), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT52), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n788), .A2(new_n791), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n811), .A2(new_n805), .B1(new_n807), .B2(G92gat), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n806), .A2(new_n810), .B1(new_n812), .B2(new_n809), .ZN(G1337gat));
  NOR3_X1   g612(.A1(new_n489), .A2(G99gat), .A3(new_n698), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n793), .A2(new_n794), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(G99gat), .B1(new_n798), .B2(new_n712), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1338gat));
  NOR3_X1   g616(.A1(new_n419), .A2(G106gat), .A3(new_n698), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n793), .A2(new_n794), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n733), .A2(new_n457), .A3(new_n734), .A4(new_n797), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G106gat), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n811), .A2(new_n818), .B1(new_n820), .B2(G106gat), .ZN(new_n824));
  OAI22_X1  g623(.A1(new_n819), .A2(new_n823), .B1(new_n824), .B2(new_n822), .ZN(G1339gat));
  AND4_X1   g624(.A1(new_n726), .A2(new_n668), .A3(new_n670), .A4(new_n698), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n725), .A2(new_n568), .A3(new_n584), .ZN(new_n827));
  INV_X1    g626(.A(new_n582), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n572), .A2(new_n575), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n558), .B1(new_n557), .B2(new_n561), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT116), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n833), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n827), .A2(new_n667), .A3(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n695), .B(KEYINPUT54), .C1(new_n683), .C2(new_n680), .ZN(new_n837));
  AOI211_X1 g636(.A(KEYINPUT54), .B(new_n682), .C1(new_n678), .C2(new_n679), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n838), .A2(new_n839), .A3(new_n691), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n680), .A2(new_n841), .A3(new_n683), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT114), .B1(new_n842), .B2(new_n692), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT55), .B(new_n837), .C1(new_n840), .C2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n696), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n836), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n678), .A2(new_n682), .A3(new_n679), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n847), .A2(new_n694), .A3(new_n841), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n839), .B1(new_n838), .B2(new_n691), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n842), .A2(KEYINPUT114), .A3(new_n692), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT115), .B1(new_n851), .B2(KEYINPUT55), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n837), .B1(new_n840), .B2(new_n843), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT115), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT55), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n846), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n827), .A2(new_n835), .A3(new_n697), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n726), .A2(new_n845), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n857), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n858), .B1(new_n862), .B2(new_n667), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n826), .B1(new_n863), .B2(new_n634), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(new_n505), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n865), .A2(new_n498), .A3(new_n504), .ZN(new_n866));
  AOI21_X1  g665(.A(G113gat), .B1(new_n866), .B2(new_n590), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n864), .A2(new_n457), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n868), .A2(new_n506), .A3(new_n488), .A4(new_n705), .ZN(new_n869));
  XNOR2_X1  g668(.A(new_n869), .B(KEYINPUT117), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n590), .A2(G113gat), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n867), .B1(new_n871), .B2(new_n872), .ZN(G1340gat));
  AOI21_X1  g672(.A(G120gat), .B1(new_n866), .B2(new_n697), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n697), .A2(G120gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n874), .B1(new_n871), .B2(new_n875), .ZN(G1341gat));
  OAI21_X1  g675(.A(G127gat), .B1(new_n870), .B2(new_n634), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n866), .A2(new_n618), .A3(new_n633), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1342gat));
  NOR2_X1   g678(.A1(new_n669), .A2(G134gat), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n866), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT118), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(G134gat), .B1(new_n870), .B2(new_n669), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n882), .A2(KEYINPUT56), .A3(new_n884), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G1343gat));
  NOR2_X1   g689(.A1(new_n753), .A2(new_n419), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n705), .A3(new_n865), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(G141gat), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n894), .A3(new_n590), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT119), .B1(new_n851), .B2(KEYINPUT55), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n853), .A2(new_n897), .A3(new_n855), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n590), .A2(new_n696), .A3(new_n844), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n859), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n669), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n633), .B1(new_n902), .B2(new_n858), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n457), .B1(new_n903), .B2(new_n826), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT57), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n711), .A2(new_n505), .A3(new_n308), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n864), .A2(KEYINPUT57), .A3(new_n419), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n907), .A2(new_n908), .A3(new_n726), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n895), .B1(new_n909), .B2(new_n894), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n911), .B1(new_n909), .B2(new_n894), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n910), .A2(KEYINPUT58), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n914));
  OAI221_X1 g713(.A(new_n895), .B1(new_n911), .B2(new_n914), .C1(new_n909), .C2(new_n894), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n913), .A2(new_n915), .ZN(G1344gat));
  INV_X1    g715(.A(G148gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n893), .A2(new_n917), .A3(new_n697), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n907), .A2(new_n908), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT59), .B(new_n917), .C1(new_n919), .C2(new_n697), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT57), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n864), .A2(new_n922), .A3(new_n419), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n668), .A2(new_n726), .A3(new_n670), .A4(new_n698), .ZN(new_n924));
  AOI22_X1  g723(.A1(new_n901), .A2(new_n669), .B1(new_n857), .B2(new_n846), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(new_n633), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n926), .B2(new_n457), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n697), .B(new_n906), .C1(new_n923), .C2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n921), .B1(new_n928), .B2(G148gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n918), .B1(new_n920), .B2(new_n929), .ZN(G1345gat));
  NAND3_X1  g729(.A1(new_n893), .A2(new_n593), .A3(new_n633), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n907), .A2(new_n634), .A3(new_n908), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n593), .B2(new_n932), .ZN(G1346gat));
  AOI21_X1  g732(.A(G162gat), .B1(new_n893), .B2(new_n667), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n667), .A2(G162gat), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n919), .B2(new_n935), .ZN(G1347gat));
  NOR3_X1   g735(.A1(new_n864), .A2(new_n506), .A3(new_n705), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n937), .A2(new_n498), .A3(new_n419), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n938), .A2(new_n269), .A3(new_n270), .A4(new_n590), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n705), .A2(new_n506), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(KEYINPUT122), .A3(new_n780), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n940), .A2(new_n941), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n705), .A2(KEYINPUT121), .A3(new_n506), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n780), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g747(.A1(new_n943), .A2(new_n868), .A3(new_n948), .A4(new_n590), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n949), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n950));
  AOI21_X1  g749(.A(KEYINPUT123), .B1(new_n949), .B2(G169gat), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n939), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT124), .ZN(G1348gat));
  NAND3_X1  g752(.A1(new_n938), .A2(new_n233), .A3(new_n697), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n943), .A2(new_n868), .A3(new_n948), .ZN(new_n955));
  OAI21_X1  g754(.A(G176gat), .B1(new_n955), .B2(new_n698), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1349gat));
  NAND4_X1  g756(.A1(new_n938), .A2(new_n243), .A3(new_n245), .A4(new_n633), .ZN(new_n958));
  OAI21_X1  g757(.A(G183gat), .B1(new_n955), .B2(new_n634), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n938), .A2(new_n230), .A3(new_n667), .ZN(new_n962));
  OAI21_X1  g761(.A(G190gat), .B1(new_n955), .B2(new_n669), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n966), .B(G190gat), .C1(new_n955), .C2(new_n669), .ZN(new_n967));
  AND3_X1   g766(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n965), .B1(new_n964), .B2(new_n967), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n962), .B1(new_n968), .B2(new_n969), .ZN(G1351gat));
  AND2_X1   g769(.A1(new_n891), .A2(new_n937), .ZN(new_n971));
  AOI21_X1  g770(.A(G197gat), .B1(new_n971), .B2(new_n590), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n712), .A2(new_n942), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n904), .A2(new_n922), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n900), .B1(new_n852), .B2(new_n856), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n669), .B1(new_n975), .B2(new_n860), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n633), .B1(new_n976), .B2(new_n858), .ZN(new_n977));
  OAI211_X1 g776(.A(KEYINPUT57), .B(new_n457), .C1(new_n977), .C2(new_n826), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n973), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n590), .A2(G197gat), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n972), .B1(new_n979), .B2(new_n980), .ZN(G1352gat));
  INV_X1    g780(.A(G204gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n971), .A2(new_n982), .A3(new_n697), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT62), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n982), .B1(new_n979), .B2(new_n697), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n984), .A2(new_n985), .ZN(G1353gat));
  INV_X1    g785(.A(KEYINPUT63), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n944), .A2(new_n945), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n753), .A2(new_n988), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n989), .B(new_n633), .C1(new_n923), .C2(new_n927), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n991));
  OAI21_X1  g790(.A(G211gat), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AOI21_X1  g791(.A(KEYINPUT126), .B1(new_n979), .B2(new_n633), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n979), .A2(KEYINPUT126), .A3(new_n633), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n990), .A2(new_n991), .ZN(new_n996));
  NAND4_X1  g795(.A1(new_n995), .A2(new_n996), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n994), .A2(KEYINPUT127), .A3(new_n997), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n999));
  OAI211_X1 g798(.A(new_n999), .B(new_n987), .C1(new_n992), .C2(new_n993), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n971), .A2(new_n206), .A3(new_n633), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .ZN(G1354gat));
  AOI21_X1  g801(.A(G218gat), .B1(new_n971), .B2(new_n667), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n669), .B1(new_n209), .B2(new_n210), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1003), .B1(new_n979), .B2(new_n1004), .ZN(G1355gat));
endmodule


