//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n583, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1236, new_n1237, new_n1238;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G218), .A2(G219), .A3(G220), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n454), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  XOR2_X1   g039(.A(new_n464), .B(KEYINPUT68), .Z(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT69), .B1(new_n468), .B2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n475));
  AND4_X1   g050(.A1(new_n472), .A2(new_n473), .A3(new_n475), .A4(new_n469), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G137), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n472), .A2(G101), .A3(G2104), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n471), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND4_X1  g055(.A1(new_n473), .A2(new_n475), .A3(G2105), .A4(new_n469), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n472), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI22_X1  g059(.A1(new_n481), .A2(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(G136), .B2(new_n476), .ZN(G162));
  NAND3_X1  g061(.A1(new_n473), .A2(new_n475), .A3(new_n469), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n472), .A2(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT4), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(new_n467), .A3(new_n469), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n472), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n494), .A2(KEYINPUT70), .A3(new_n496), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n492), .B1(new_n499), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT5), .B(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G62), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n504), .A2(new_n505), .B1(G75), .B2(G543), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n503), .A2(KEYINPUT72), .A3(G62), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n502), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(new_n503), .A3(KEYINPUT71), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n515), .A2(G88), .A3(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n521), .B1(new_n516), .B2(new_n517), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n508), .A2(new_n524), .ZN(G166));
  OAI211_X1 g100(.A(G51), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n527));
  NAND2_X1  g102(.A1(G76), .A2(G543), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(new_n502), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n510), .A2(new_n509), .ZN(new_n531));
  INV_X1    g106(.A(G63), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n531), .A2(new_n532), .B1(new_n527), .B2(new_n528), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n530), .B1(G651), .B2(new_n533), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT73), .B(G89), .Z(new_n535));
  NAND3_X1  g110(.A1(new_n515), .A2(new_n519), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  NAND3_X1  g113(.A1(new_n515), .A2(G90), .A3(new_n519), .ZN(new_n539));
  OAI21_X1  g114(.A(G64), .B1(new_n510), .B2(new_n509), .ZN(new_n540));
  NAND2_X1  g115(.A1(G77), .A2(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(G651), .B1(G52), .B2(new_n522), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(G171));
  AOI22_X1  g120(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n502), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n515), .A2(G81), .A3(new_n519), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT74), .B(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n522), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n548), .A2(KEYINPUT75), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(KEYINPUT75), .B1(new_n548), .B2(new_n550), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n547), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT76), .Z(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND3_X1  g135(.A1(new_n515), .A2(G91), .A3(new_n519), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n522), .A2(new_n562), .A3(G53), .ZN(new_n563));
  OAI211_X1 g138(.A(G53), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT9), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n531), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G651), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n561), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT77), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n573));
  NAND4_X1  g148(.A1(new_n561), .A2(new_n566), .A3(new_n573), .A4(new_n570), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n544), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n539), .A2(new_n543), .A3(KEYINPUT78), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G301));
  NAND2_X1  g156(.A1(new_n506), .A2(new_n507), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n583), .A2(new_n520), .A3(new_n523), .ZN(G303));
  NOR3_X1   g159(.A1(new_n510), .A2(new_n509), .A3(G74), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT79), .B1(new_n585), .B2(new_n502), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n587), .B(G651), .C1(new_n503), .C2(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n515), .A2(G87), .A3(new_n519), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n522), .A2(G49), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n531), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G48), .B2(new_n522), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n515), .A2(G86), .A3(new_n519), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G305));
  NAND3_X1  g173(.A1(new_n515), .A2(G85), .A3(new_n519), .ZN(new_n599));
  OAI21_X1  g174(.A(G60), .B1(new_n510), .B2(new_n509), .ZN(new_n600));
  NAND2_X1  g175(.A1(G72), .A2(G543), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G47), .B2(new_n522), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(G290));
  NAND3_X1  g179(.A1(new_n515), .A2(G92), .A3(new_n519), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n515), .A2(KEYINPUT10), .A3(G92), .A4(new_n519), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n531), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT80), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(G651), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n522), .A2(G54), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n609), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n580), .ZN(G284));
  AOI21_X1  g196(.A(new_n620), .B1(G868), .B2(new_n580), .ZN(G321));
  NAND2_X1  g197(.A1(G286), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n575), .B2(G868), .ZN(G297));
  OAI21_X1  g199(.A(new_n623), .B1(new_n575), .B2(G868), .ZN(G280));
  INV_X1    g200(.A(G860), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n619), .B1(G559), .B2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT81), .ZN(G148));
  INV_X1    g203(.A(G868), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n553), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n619), .A2(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(new_n629), .ZN(G323));
  XOR2_X1   g207(.A(KEYINPUT82), .B(KEYINPUT11), .Z(new_n633));
  XNOR2_X1  g208(.A(G323), .B(new_n633), .ZN(G282));
  AND2_X1   g209(.A1(new_n476), .A2(G135), .ZN(new_n635));
  INV_X1    g210(.A(G123), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n472), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  OAI22_X1  g213(.A1(new_n481), .A2(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g214(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n641), .A2(G2096), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n641), .A2(G2096), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n642), .A2(new_n646), .A3(new_n647), .ZN(G156));
  XNOR2_X1  g223(.A(G2427), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2430), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(KEYINPUT14), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT84), .B(KEYINPUT85), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2443), .B(G2446), .Z(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2451), .B(G2454), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n656), .A2(new_n661), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  INV_X1    g241(.A(new_n663), .ZN(new_n667));
  INV_X1    g242(.A(new_n664), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n656), .A2(new_n661), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(KEYINPUT86), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n672), .B(new_n667), .C1(new_n668), .C2(new_n669), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n666), .B1(new_n671), .B2(new_n673), .ZN(G401));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2072), .B(G2078), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT18), .Z(new_n679));
  INV_X1    g254(.A(KEYINPUT87), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n677), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(new_n680), .B2(new_n676), .ZN(new_n682));
  INV_X1    g257(.A(new_n675), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n676), .B(KEYINPUT17), .Z(new_n684));
  INV_X1    g259(.A(new_n677), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n682), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n684), .A2(new_n685), .A3(new_n675), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n679), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G2096), .B(G2100), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G227));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT19), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  AND2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT20), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n695), .A2(new_n696), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n694), .A2(new_n697), .A3(new_n700), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n699), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n698), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n702), .A2(new_n701), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(new_n704), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n691), .B1(new_n706), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1981), .B(G1986), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n703), .A2(new_n705), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n710), .A2(new_n704), .ZN(new_n715));
  INV_X1    g290(.A(new_n691), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AND3_X1   g292(.A1(new_n712), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n713), .B1(new_n712), .B2(new_n717), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n718), .A2(new_n719), .ZN(G229));
  INV_X1    g295(.A(G288), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n722), .B2(G23), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT33), .B(G1976), .ZN(new_n725));
  NAND2_X1  g300(.A1(G166), .A2(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G16), .B2(G22), .ZN(new_n727));
  INV_X1    g302(.A(G1971), .ZN(new_n728));
  OAI22_X1  g303(.A1(new_n724), .A2(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n728), .B2(new_n727), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n722), .A2(G6), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n596), .A2(new_n597), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n722), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT32), .B(G1981), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT90), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n733), .B(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n724), .B2(new_n725), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n730), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  NOR2_X1   g316(.A1(G25), .A2(G29), .ZN(new_n742));
  INV_X1    g317(.A(G119), .ZN(new_n743));
  OR3_X1    g318(.A1(new_n481), .A2(KEYINPUT88), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(KEYINPUT88), .B1(new_n481), .B2(new_n743), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n747));
  INV_X1    g322(.A(G107), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G2105), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n476), .B2(G131), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n742), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT35), .B(G1991), .Z(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  MUX2_X1   g331(.A(G24), .B(G290), .S(G16), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1986), .ZN(new_n758));
  INV_X1    g333(.A(new_n753), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n754), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n740), .A2(new_n741), .A3(new_n756), .A4(new_n760), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT36), .ZN(new_n762));
  INV_X1    g337(.A(G29), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G32), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT98), .B(KEYINPUT26), .ZN(new_n765));
  AND3_X1   g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n472), .A2(G105), .A3(G2104), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G129), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(new_n481), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n476), .A2(G141), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n764), .B1(new_n773), .B2(new_n763), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT27), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1996), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n722), .A2(G20), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT23), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(new_n575), .B2(new_n722), .ZN(new_n779));
  INV_X1    g354(.A(G1956), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n722), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n722), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT100), .ZN(new_n784));
  INV_X1    g359(.A(G1961), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n489), .A2(new_n491), .ZN(new_n787));
  AND3_X1   g362(.A1(new_n494), .A2(KEYINPUT70), .A3(new_n496), .ZN(new_n788));
  AOI21_X1  g363(.A(KEYINPUT70), .B1(new_n494), .B2(new_n496), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(G29), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n763), .A2(G27), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n786), .B1(G2078), .B2(new_n794), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n784), .A2(new_n785), .B1(new_n793), .B2(new_n443), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n776), .A2(new_n781), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n722), .A2(G21), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G286), .B2(G16), .ZN(new_n799));
  INV_X1    g374(.A(G1966), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT99), .ZN(new_n802));
  NAND2_X1  g377(.A1(G160), .A2(G29), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G34), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(new_n763), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n803), .A2(G2084), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT31), .B(G11), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT30), .B(G28), .Z(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(G29), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(new_n640), .B2(G29), .ZN(new_n811));
  AOI21_X1  g386(.A(G2084), .B1(new_n803), .B2(new_n806), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n800), .B2(new_n799), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n802), .A2(new_n807), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G16), .A2(G19), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n554), .B2(G16), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n816), .A2(G1341), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(G1341), .ZN(new_n818));
  NOR2_X1   g393(.A1(G29), .A2(G33), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT94), .ZN(new_n820));
  NAND2_X1  g395(.A1(G103), .A2(G2104), .ZN(new_n821));
  OAI21_X1  g396(.A(KEYINPUT95), .B1(new_n821), .B2(G2105), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT95), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n823), .A2(new_n472), .A3(G103), .A4(G2104), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(KEYINPUT25), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT25), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n822), .A2(new_n824), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n467), .A2(new_n469), .A3(G127), .ZN(new_n829));
  INV_X1    g404(.A(G115), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n466), .ZN(new_n831));
  AOI22_X1  g406(.A1(new_n826), .A2(new_n828), .B1(new_n831), .B2(G2105), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n476), .A2(G139), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n820), .B1(new_n834), .B2(new_n763), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT96), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(new_n442), .ZN(new_n837));
  NOR4_X1   g412(.A1(new_n814), .A2(new_n817), .A3(new_n818), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n763), .A2(G35), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(G162), .B2(new_n763), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT29), .Z(new_n841));
  INV_X1    g416(.A(G2090), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n841), .A2(new_n842), .B1(new_n836), .B2(new_n442), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n763), .A2(G26), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT28), .Z(new_n845));
  INV_X1    g420(.A(KEYINPUT92), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n476), .A2(new_n846), .A3(G140), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n473), .A2(new_n475), .A3(new_n472), .A4(new_n469), .ZN(new_n848));
  INV_X1    g423(.A(G140), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT92), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(new_n472), .B2(G116), .ZN(new_n852));
  OR3_X1    g427(.A1(KEYINPUT93), .A2(G104), .A3(G2105), .ZN(new_n853));
  OAI21_X1  g428(.A(KEYINPUT93), .B1(G104), .B2(G2105), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n481), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n856), .B2(G128), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n845), .B1(new_n858), .B2(G29), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(G2067), .ZN(new_n860));
  NOR2_X1   g435(.A1(G4), .A2(G16), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT91), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n619), .B2(new_n722), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(G1348), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n838), .A2(new_n843), .A3(new_n860), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n841), .A2(new_n842), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT101), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n797), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n762), .A2(new_n868), .ZN(G150));
  INV_X1    g444(.A(G150), .ZN(G311));
  AOI21_X1  g445(.A(new_n617), .B1(new_n607), .B2(new_n608), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(G559), .ZN(new_n872));
  XOR2_X1   g447(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(G80), .A2(G543), .ZN(new_n875));
  INV_X1    g450(.A(G67), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n531), .B2(new_n876), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n877), .A2(G651), .B1(G55), .B2(new_n522), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n515), .A2(G93), .A3(new_n519), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n553), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n547), .B(new_n880), .C1(new_n551), .C2(new_n552), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n874), .B(new_n884), .Z(new_n885));
  OR2_X1    g460(.A1(new_n885), .A2(KEYINPUT39), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(KEYINPUT39), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n626), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n880), .A2(new_n626), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(G145));
  XNOR2_X1  g466(.A(new_n640), .B(new_n479), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(G162), .Z(new_n893));
  INV_X1    g468(.A(new_n773), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n858), .A2(new_n834), .ZN(new_n895));
  INV_X1    g470(.A(new_n497), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n787), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n851), .A2(new_n832), .A3(new_n833), .A4(new_n857), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n895), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n897), .B1(new_n895), .B2(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n894), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OR2_X1    g476(.A1(G106), .A2(G2105), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n902), .B(G2104), .C1(G118), .C2(new_n472), .ZN(new_n903));
  INV_X1    g478(.A(G130), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(new_n481), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n905), .B1(G142), .B2(new_n476), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n746), .A2(new_n644), .A3(new_n750), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n644), .B1(new_n746), .B2(new_n750), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n644), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n751), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n746), .A2(new_n644), .A3(new_n750), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n906), .A3(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n897), .ZN(new_n916));
  INV_X1    g491(.A(new_n898), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n851), .A2(new_n857), .B1(new_n832), .B2(new_n833), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n895), .A2(new_n897), .A3(new_n898), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n773), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n901), .A2(new_n915), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n910), .A2(new_n914), .ZN(new_n927));
  INV_X1    g502(.A(new_n921), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n773), .B1(new_n919), .B2(new_n920), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n922), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n925), .B(new_n927), .C1(new_n928), .C2(new_n929), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n901), .A2(new_n915), .A3(KEYINPUT104), .A4(new_n921), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n893), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n930), .A2(KEYINPUT105), .A3(new_n893), .A4(new_n922), .ZN(new_n939));
  INV_X1    g514(.A(G37), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n943), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g519(.A1(new_n881), .A2(new_n629), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n884), .B(new_n631), .Z(new_n946));
  NAND3_X1  g521(.A1(new_n871), .A2(new_n572), .A3(new_n574), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n871), .B1(new_n572), .B2(new_n574), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n575), .A2(new_n619), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n952), .A2(KEYINPUT41), .A3(new_n947), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT41), .B1(new_n952), .B2(new_n947), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n951), .B1(new_n946), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n599), .A2(new_n603), .A3(KEYINPUT106), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT106), .B1(new_n599), .B2(new_n603), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n721), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  NAND2_X1  g536(.A1(G290), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n599), .A2(new_n603), .A3(KEYINPUT106), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(G288), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n732), .B1(new_n508), .B2(new_n524), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n583), .A2(new_n520), .A3(new_n523), .A4(G305), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n960), .A2(new_n964), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  AOI22_X1  g543(.A1(new_n960), .A2(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n957), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n960), .A2(new_n964), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n965), .A2(new_n966), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(KEYINPUT107), .A3(new_n967), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT42), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n967), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n976), .B1(KEYINPUT42), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n956), .B(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n945), .B1(new_n979), .B2(new_n629), .ZN(G295));
  OAI21_X1  g555(.A(new_n945), .B1(new_n979), .B2(new_n629), .ZN(G331));
  AND2_X1   g556(.A1(G286), .A2(new_n544), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n982), .B1(new_n580), .B2(G168), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n548), .A2(new_n550), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT75), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n548), .A2(KEYINPUT75), .A3(new_n550), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n880), .B1(new_n988), .B2(new_n547), .ZN(new_n989));
  INV_X1    g564(.A(new_n883), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n983), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n539), .A2(new_n543), .A3(KEYINPUT78), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT78), .B1(new_n539), .B2(new_n543), .ZN(new_n993));
  OAI21_X1  g568(.A(G168), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(G286), .A2(new_n544), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n996), .A2(new_n882), .A3(new_n883), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n950), .B1(new_n991), .B2(new_n997), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n996), .A2(new_n882), .A3(new_n883), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n996), .B1(new_n882), .B2(new_n883), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n998), .B1(new_n955), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n975), .ZN(new_n1003));
  AOI21_X1  g578(.A(G37), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT43), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n1006));
  INV_X1    g581(.A(new_n950), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n999), .B2(new_n1000), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n997), .B(new_n991), .C1(new_n953), .C2(new_n954), .ZN(new_n1009));
  AOI221_X4 g584(.A(new_n1006), .B1(new_n970), .B2(new_n974), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT108), .B1(new_n1011), .B2(new_n975), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1004), .B(new_n1005), .C1(new_n1010), .C2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT109), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1006), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(KEYINPUT108), .A3(new_n975), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT109), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n1005), .A4(new_n1004), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1011), .A2(new_n975), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1005), .B1(new_n1004), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1014), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1017), .A2(KEYINPUT43), .A3(new_n1004), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1020), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n940), .B1(new_n1011), .B2(new_n975), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1005), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  MUX2_X1   g603(.A(new_n1023), .B(new_n1028), .S(KEYINPUT44), .Z(G397));
  INV_X1    g604(.A(G1384), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n492), .B2(new_n497), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n471), .A2(G40), .A3(new_n477), .A4(new_n478), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT45), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n894), .A2(new_n1036), .A3(G1996), .ZN(new_n1037));
  XOR2_X1   g612(.A(new_n1037), .B(KEYINPUT110), .Z(new_n1038));
  INV_X1    g613(.A(G2067), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n858), .B(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n894), .B2(G1996), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1038), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n752), .A2(new_n754), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n751), .A2(new_n755), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1036), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(G290), .B(G1986), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(new_n1036), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n790), .A2(KEYINPUT45), .A3(new_n1030), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1032), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n800), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1384), .B1(new_n896), .B2(new_n787), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1055));
  AOI21_X1  g630(.A(new_n1032), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1052), .B(G168), .C1(G2084), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n1059));
  OAI21_X1  g634(.A(G8), .B1(new_n1059), .B2(KEYINPUT51), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(KEYINPUT51), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1058), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1057), .A2(G2084), .ZN(new_n1064));
  AOI21_X1  g639(.A(G1966), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1065));
  OAI211_X1 g640(.A(G8), .B(G286), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1062), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT62), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1068), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n1066), .A4(new_n1063), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT45), .B1(new_n790), .B2(new_n1030), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1033), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI22_X1  g650(.A1(new_n1075), .A2(G1971), .B1(new_n1057), .B2(G2090), .ZN(new_n1076));
  NAND2_X1  g651(.A1(G303), .A2(G8), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(KEYINPUT55), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1079), .A3(G8), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1054), .A2(new_n1033), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n721), .A2(G1976), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(G8), .A3(new_n1082), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1083), .A2(KEYINPUT112), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(KEYINPUT112), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(KEYINPUT52), .A3(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n721), .A2(G1976), .ZN(new_n1087));
  OR3_X1    g662(.A1(new_n1083), .A2(KEYINPUT52), .A3(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT113), .B(G1981), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n732), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G305), .A2(G1981), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1090), .A2(KEYINPUT49), .A3(new_n1091), .ZN(new_n1092));
  XOR2_X1   g667(.A(new_n1092), .B(KEYINPUT114), .Z(new_n1093));
  NAND2_X1  g668(.A1(new_n1081), .A2(G8), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT49), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1080), .A2(new_n1086), .A3(new_n1088), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT50), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n499), .A2(new_n500), .ZN(new_n1100));
  AOI21_X1  g675(.A(G1384), .B1(new_n1100), .B2(new_n787), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1055), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1032), .B1(new_n1031), .B2(new_n1102), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1099), .A2(new_n1101), .B1(new_n1103), .B2(KEYINPUT115), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1103), .A2(KEYINPUT115), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1104), .A2(new_n842), .A3(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(G1971), .B2(new_n1075), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1079), .B1(new_n1107), .B2(G8), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1098), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1074), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1110), .B(new_n443), .C1(new_n1101), .C2(KEYINPUT45), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1111), .A2(new_n1112), .B1(new_n1057), .B2(new_n785), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1049), .A2(new_n1050), .A3(KEYINPUT53), .A4(new_n443), .ZN(new_n1114));
  AOI21_X1  g689(.A(G301), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1069), .A2(new_n1072), .A3(new_n1109), .A4(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1097), .ZN(new_n1117));
  OR2_X1    g692(.A1(G288), .A2(G1976), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1090), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1094), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1097), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1080), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1119), .A2(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1101), .A2(new_n1099), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1103), .A2(KEYINPUT115), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1103), .A2(KEYINPUT115), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n780), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT56), .B(G2072), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1075), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n566), .B2(KEYINPUT118), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(new_n571), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1128), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(G1348), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1099), .B1(new_n790), .B2(new_n1030), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1033), .B1(new_n1031), .B2(new_n1102), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1054), .A2(new_n1039), .A3(new_n1033), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1133), .A2(new_n871), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1132), .ZN(new_n1141));
  AOI21_X1  g716(.A(G1956), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n1075), .A2(new_n1129), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1141), .B1(new_n1144), .B2(KEYINPUT119), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1128), .A2(KEYINPUT119), .A3(new_n1130), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1140), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n619), .A2(KEYINPUT121), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT60), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n1139), .B2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n871), .B(KEYINPUT121), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1137), .A2(KEYINPUT60), .A3(new_n1151), .A4(new_n1138), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1139), .A2(new_n1149), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1073), .A2(new_n1074), .A3(G1996), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT58), .B(G1341), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1156), .B1(new_n1054), .B2(new_n1033), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n554), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT59), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1160), .B(new_n554), .C1(new_n1155), .C2(new_n1157), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1159), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1154), .A2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1164));
  OAI21_X1  g739(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1165), .B2(new_n1133), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g742(.A(KEYINPUT61), .B(new_n1133), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1147), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT54), .ZN(new_n1170));
  OAI21_X1  g745(.A(KEYINPUT53), .B1(KEYINPUT124), .B2(G2078), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1032), .A2(KEYINPUT123), .ZN(new_n1172));
  AOI211_X1 g747(.A(new_n1171), .B(new_n1172), .C1(KEYINPUT124), .C2(G2078), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1054), .A2(KEYINPUT45), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1032), .A2(KEYINPUT123), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1113), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1178), .A2(new_n580), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1170), .B1(new_n1179), .B2(new_n1115), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1070), .A2(new_n1066), .A3(new_n1063), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1178), .A2(G171), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1113), .A2(G301), .A3(new_n1114), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1182), .A2(KEYINPUT54), .A3(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1180), .A2(new_n1109), .A3(new_n1181), .A4(new_n1184), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1116), .B(new_n1123), .C1(new_n1169), .C2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g761(.A(G8), .B(G168), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1076), .A2(G8), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1190), .A2(new_n1078), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g767(.A(KEYINPUT117), .B1(new_n1192), .B2(new_n1098), .ZN(new_n1193));
  AND4_X1   g768(.A1(new_n1080), .A2(new_n1086), .A3(new_n1088), .A4(new_n1097), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1079), .B1(new_n1076), .B2(G8), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n1195), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT117), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1194), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1193), .A2(new_n1198), .ZN(new_n1199));
  NOR3_X1   g774(.A1(new_n1098), .A2(new_n1108), .A3(new_n1187), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT116), .ZN(new_n1201));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1108), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1194), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(KEYINPUT116), .B1(new_n1204), .B2(new_n1187), .ZN(new_n1205));
  AOI21_X1  g780(.A(new_n1199), .B1(new_n1202), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1048), .B1(new_n1186), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n851), .A2(new_n1039), .A3(new_n857), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1035), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OR2_X1    g785(.A1(new_n1035), .A2(G1996), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT46), .ZN(new_n1212));
  NOR2_X1   g787(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  XOR2_X1   g788(.A(new_n1213), .B(KEYINPUT125), .Z(new_n1214));
  AOI21_X1  g789(.A(new_n1035), .B1(new_n1040), .B2(new_n773), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1215), .B1(new_n1212), .B2(new_n1211), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT47), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1217), .B(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1046), .ZN(new_n1220));
  NOR3_X1   g795(.A1(new_n1035), .A2(G1986), .A3(G290), .ZN(new_n1221));
  XOR2_X1   g796(.A(new_n1221), .B(KEYINPUT48), .Z(new_n1222));
  AOI211_X1 g797(.A(new_n1210), .B(new_n1219), .C1(new_n1220), .C2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1207), .A2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g799(.A1(G227), .A2(new_n462), .ZN(new_n1226));
  OAI21_X1  g800(.A(new_n1226), .B1(new_n718), .B2(new_n719), .ZN(new_n1227));
  NOR2_X1   g801(.A1(G401), .A2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g802(.A(new_n1228), .B1(new_n937), .B2(new_n941), .ZN(new_n1229));
  AOI21_X1  g803(.A(new_n1021), .B1(new_n1013), .B2(KEYINPUT109), .ZN(new_n1230));
  AOI211_X1 g804(.A(KEYINPUT126), .B(new_n1229), .C1(new_n1230), .C2(new_n1019), .ZN(new_n1231));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n1232));
  INV_X1    g806(.A(new_n1229), .ZN(new_n1233));
  AOI21_X1  g807(.A(new_n1232), .B1(new_n1023), .B2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g808(.A1(new_n1231), .A2(new_n1234), .ZN(G308));
  NAND2_X1  g809(.A1(new_n1023), .A2(new_n1233), .ZN(new_n1236));
  NAND2_X1  g810(.A1(new_n1236), .A2(KEYINPUT126), .ZN(new_n1237));
  NAND3_X1  g811(.A1(new_n1023), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1238));
  NAND2_X1  g812(.A1(new_n1237), .A2(new_n1238), .ZN(G225));
endmodule


