//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1129, new_n1130,
    new_n1131;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(KEYINPUT70), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n467), .B2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT69), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n468), .A2(G137), .A3(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT71), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n468), .A2(KEYINPUT71), .A3(G137), .A4(new_n473), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT70), .B(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n469), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G101), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(KEYINPUT3), .B(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G125), .ZN(new_n485));
  INV_X1    g060(.A(G113), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(new_n462), .ZN(new_n487));
  INV_X1    g062(.A(new_n473), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n483), .A2(new_n490), .ZN(G160));
  OAI221_X1 g066(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n473), .C2(G112), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n468), .A2(new_n469), .ZN(new_n493));
  INV_X1    g068(.A(G136), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n463), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT3), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n479), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(new_n473), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(G124), .B2(new_n499), .ZN(G162));
  NAND2_X1  g075(.A1(new_n473), .A2(G138), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT73), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n470), .B2(new_n472), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n468), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n502), .A2(new_n506), .A3(KEYINPUT4), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n484), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n508), .B1(new_n501), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n505), .A2(KEYINPUT74), .A3(new_n509), .A4(new_n484), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g089(.A(G126), .B(new_n496), .C1(new_n479), .C2(new_n497), .ZN(new_n515));
  NAND2_X1  g090(.A1(G114), .A2(G2104), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G2105), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n469), .A2(G102), .A3(G2104), .ZN(new_n519));
  AOI21_X1  g094(.A(KEYINPUT72), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n469), .B1(new_n515), .B2(new_n516), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  INV_X1    g097(.A(new_n519), .ZN(new_n523));
  NOR3_X1   g098(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n514), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(G164));
  XNOR2_X1  g101(.A(KEYINPUT6), .B(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G50), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT75), .ZN(new_n531));
  INV_X1    g106(.A(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT5), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT5), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G543), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n536), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n527), .ZN(new_n539));
  INV_X1    g114(.A(G88), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n537), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n531), .A2(new_n541), .ZN(G303));
  INV_X1    g117(.A(G303), .ZN(G166));
  XNOR2_X1  g118(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT77), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n536), .A2(G63), .A3(G651), .ZN(new_n548));
  INV_X1    g123(.A(G51), .ZN(new_n549));
  INV_X1    g124(.A(G89), .ZN(new_n550));
  OAI221_X1 g125(.A(new_n548), .B1(new_n528), .B2(new_n549), .C1(new_n539), .C2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n547), .A2(new_n551), .ZN(G168));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n533), .A2(new_n535), .ZN(new_n554));
  INV_X1    g129(.A(G64), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G651), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT78), .ZN(new_n558));
  INV_X1    g133(.A(G90), .ZN(new_n559));
  INV_X1    g134(.A(G52), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n539), .A2(new_n559), .B1(new_n560), .B2(new_n528), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G301));
  INV_X1    g138(.A(G301), .ZN(G171));
  INV_X1    g139(.A(G81), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n539), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n536), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n567), .A2(new_n538), .ZN(new_n568));
  AOI211_X1 g143(.A(new_n566), .B(new_n568), .C1(G43), .C2(new_n529), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G188));
  NAND2_X1  g150(.A1(new_n529), .A2(G53), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT9), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n536), .A2(G65), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT79), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n538), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n539), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n581), .B1(G91), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n577), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G168), .ZN(G286));
  OAI21_X1  g160(.A(G651), .B1(new_n536), .B2(G74), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT80), .ZN(new_n587));
  INV_X1    g162(.A(G87), .ZN(new_n588));
  INV_X1    g163(.A(G49), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n539), .A2(new_n588), .B1(new_n589), .B2(new_n528), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G288));
  AOI22_X1  g168(.A1(new_n536), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n538), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  INV_X1    g171(.A(G48), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n539), .A2(new_n596), .B1(new_n597), .B2(new_n528), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n595), .A2(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n536), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n539), .A2(new_n604), .B1(new_n605), .B2(new_n528), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G290));
  NAND2_X1  g183(.A1(G301), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OR3_X1    g185(.A1(new_n539), .A2(KEYINPUT10), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT10), .B1(new_n539), .B2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n536), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G54), .ZN(new_n615));
  OAI22_X1  g190(.A1(new_n614), .A2(new_n538), .B1(new_n528), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n609), .B1(G868), .B2(new_n617), .ZN(G284));
  XNOR2_X1  g193(.A(G284), .B(KEYINPUT82), .ZN(G321));
  NAND2_X1  g194(.A1(G286), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(G299), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(G868), .B2(new_n621), .ZN(G297));
  OAI21_X1  g197(.A(new_n620), .B1(G868), .B2(new_n621), .ZN(G280));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n617), .B1(new_n624), .B2(G860), .ZN(G148));
  INV_X1    g200(.A(new_n617), .ZN(new_n626));
  OAI21_X1  g201(.A(G868), .B1(new_n626), .B2(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g204(.A1(new_n481), .A2(new_n484), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n633), .A2(KEYINPUT83), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n632), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n499), .A2(G123), .ZN(new_n636));
  OAI221_X1 g211(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n473), .C2(G111), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n493), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n633), .A2(KEYINPUT83), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n635), .A2(new_n640), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2435), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2438), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2451), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n653), .B(new_n654), .Z(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(G14), .ZN(G401));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2096), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n633), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n659), .A2(new_n660), .ZN(new_n666));
  AOI21_X1  g241(.A(KEYINPUT18), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n664), .B(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT85), .ZN(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n670), .A2(new_n671), .ZN(new_n677));
  AOI22_X1  g252(.A1(new_n675), .A2(new_n676), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  OR3_X1    g253(.A1(new_n672), .A2(new_n677), .A3(new_n674), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n678), .B(new_n679), .C1(new_n676), .C2(new_n675), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(G1986), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT22), .B(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G229));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT99), .B(G28), .Z(new_n688));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT100), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n689), .B2(new_n688), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n481), .A2(G105), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT98), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n499), .A2(G129), .ZN(new_n695));
  NAND3_X1  g270(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT26), .Z(new_n697));
  INV_X1    g272(.A(new_n493), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G141), .ZN(new_n699));
  NAND4_X1  g274(.A1(new_n694), .A2(new_n695), .A3(new_n697), .A4(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G32), .B(new_n700), .S(G29), .Z(new_n701));
  XOR2_X1   g276(.A(KEYINPUT27), .B(G1996), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(G16), .A2(G19), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n569), .B2(G16), .ZN(new_n705));
  AOI211_X1 g280(.A(new_n692), .B(new_n703), .C1(G1341), .C2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT31), .B(G11), .Z(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G21), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G168), .B2(G16), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n707), .B1(new_n709), .B2(G1966), .ZN(new_n710));
  OAI221_X1 g285(.A(new_n710), .B1(G1341), .B2(new_n705), .C1(G1966), .C2(new_n709), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n639), .A2(new_n687), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G4), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n617), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT93), .B(G1348), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT94), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n715), .B(new_n717), .ZN(new_n718));
  NOR3_X1   g293(.A1(new_n711), .A2(new_n712), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n713), .A2(KEYINPUT23), .A3(G20), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT23), .ZN(new_n721));
  INV_X1    g296(.A(G20), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G16), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n723), .C1(new_n621), .C2(new_n713), .ZN(new_n724));
  INV_X1    g299(.A(G1956), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(KEYINPUT24), .A2(G34), .ZN(new_n727));
  NOR2_X1   g302(.A1(KEYINPUT24), .A2(G34), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n727), .A2(new_n728), .A3(G29), .ZN(new_n729));
  INV_X1    g304(.A(G160), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G29), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n687), .A2(G27), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G164), .B2(new_n687), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2078), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT96), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n687), .A2(G26), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n738), .B(new_n739), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n499), .A2(G128), .ZN(new_n741));
  OAI221_X1 g316(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n473), .C2(G116), .ZN(new_n742));
  INV_X1    g317(.A(G140), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n493), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n740), .B1(new_n745), .B2(new_n687), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2067), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n733), .A2(new_n736), .A3(new_n747), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n706), .A2(new_n719), .A3(new_n726), .A4(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n713), .A2(G23), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n592), .B2(new_n713), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT91), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT33), .B(G1976), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n713), .A2(G22), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G166), .B2(new_n713), .ZN(new_n757));
  INV_X1    g332(.A(G1971), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(G305), .A2(G16), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n713), .A2(G6), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n762), .B(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT32), .B(G1981), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n755), .A2(new_n759), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n750), .B1(new_n769), .B2(KEYINPUT34), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n769), .A2(new_n750), .A3(KEYINPUT34), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT34), .ZN(new_n773));
  INV_X1    g348(.A(new_n769), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n771), .A2(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT36), .ZN(new_n776));
  NOR2_X1   g351(.A1(G25), .A2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G131), .ZN(new_n778));
  OAI21_X1  g353(.A(G2104), .B1(new_n473), .B2(G107), .ZN(new_n779));
  NOR2_X1   g354(.A1(G95), .A2(G2105), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT86), .ZN(new_n781));
  OAI22_X1  g356(.A1(new_n493), .A2(new_n778), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G119), .B2(new_n499), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT87), .Z(new_n784));
  AOI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT88), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT35), .B(G1991), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G24), .B(G290), .S(G16), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1986), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n775), .A2(new_n776), .A3(new_n788), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n774), .A2(new_n773), .ZN(new_n793));
  INV_X1    g368(.A(new_n772), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n793), .B(new_n788), .C1(new_n794), .C2(new_n770), .ZN(new_n795));
  OAI21_X1  g370(.A(KEYINPUT36), .B1(new_n795), .B2(new_n790), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n749), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT25), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n698), .A2(G139), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n484), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT97), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n799), .B(new_n800), .C1(new_n802), .C2(new_n473), .ZN(new_n803));
  MUX2_X1   g378(.A(G33), .B(new_n803), .S(G29), .Z(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G2072), .Z(new_n805));
  INV_X1    g380(.A(KEYINPUT101), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G5), .B2(G16), .ZN(new_n807));
  OR3_X1    g382(.A1(new_n806), .A2(G5), .A3(G16), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n807), .B(new_n808), .C1(G301), .C2(new_n713), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT102), .B(G1961), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G29), .A2(G35), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G162), .B2(G29), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT29), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(G2090), .Z(new_n815));
  NAND4_X1  g390(.A1(new_n797), .A2(new_n805), .A3(new_n811), .A4(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  XOR2_X1   g392(.A(KEYINPUT104), .B(G860), .Z(new_n818));
  INV_X1    g393(.A(G93), .ZN(new_n819));
  INV_X1    g394(.A(G55), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n539), .A2(new_n819), .B1(new_n820), .B2(new_n528), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n536), .A2(G67), .ZN(new_n822));
  NAND2_X1  g397(.A1(G80), .A2(G543), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n538), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n818), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  NOR2_X1   g401(.A1(new_n821), .A2(new_n824), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT103), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n569), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n617), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n829), .B(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n826), .B1(new_n833), .B2(new_n818), .ZN(G145));
  NOR2_X1   g409(.A1(new_n521), .A2(new_n523), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT106), .ZN(new_n836));
  AND3_X1   g411(.A1(new_n507), .A2(new_n836), .A3(new_n513), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n507), .B2(new_n513), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n744), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n700), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(new_n803), .ZN(new_n842));
  INV_X1    g417(.A(G142), .ZN(new_n843));
  OR3_X1    g418(.A1(new_n493), .A2(KEYINPUT107), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n499), .A2(G130), .ZN(new_n845));
  OAI221_X1 g420(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n473), .C2(G118), .ZN(new_n846));
  OAI21_X1  g421(.A(KEYINPUT107), .B1(new_n493), .B2(new_n843), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n844), .A2(new_n845), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(new_n631), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n783), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT108), .B1(new_n842), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n842), .B(new_n850), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(KEYINPUT108), .ZN(new_n853));
  XNOR2_X1  g428(.A(G162), .B(KEYINPUT105), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G160), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n639), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n856), .ZN(new_n858));
  AOI21_X1  g433(.A(G37), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT40), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n857), .A2(new_n862), .A3(new_n859), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(G395));
  INV_X1    g439(.A(G305), .ZN(new_n865));
  XNOR2_X1  g440(.A(G290), .B(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G166), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n592), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT42), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n617), .B1(G299), .B2(KEYINPUT109), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(KEYINPUT109), .B2(G299), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n626), .A2(G299), .A3(KEYINPUT109), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT41), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n626), .A2(G559), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n829), .B(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n873), .B(KEYINPUT110), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n869), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(G868), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(G868), .B2(new_n827), .ZN(G295));
  OAI21_X1  g457(.A(new_n881), .B1(G868), .B2(new_n827), .ZN(G331));
  XNOR2_X1  g458(.A(G168), .B(G301), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n829), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n874), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT111), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n867), .B(G288), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n874), .A2(KEYINPUT111), .A3(new_n885), .ZN(new_n890));
  INV_X1    g465(.A(new_n885), .ZN(new_n891));
  INV_X1    g466(.A(new_n873), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n888), .A2(new_n889), .A3(new_n890), .A4(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n886), .B1(new_n878), .B2(new_n885), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n868), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT112), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n894), .A2(new_n897), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n886), .A2(new_n887), .B1(new_n892), .B2(new_n891), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n889), .B1(new_n902), .B2(new_n890), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT44), .B1(new_n904), .B2(KEYINPUT43), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT43), .B1(new_n901), .B2(new_n903), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n894), .A2(new_n896), .A3(new_n907), .A4(new_n897), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  OAI22_X1  g484(.A1(new_n900), .A2(new_n905), .B1(KEYINPUT44), .B2(new_n909), .ZN(G397));
  INV_X1    g485(.A(KEYINPUT45), .ZN(new_n911));
  INV_X1    g486(.A(new_n835), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n514), .A2(KEYINPUT106), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n507), .A2(new_n836), .A3(new_n513), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n911), .B1(new_n915), .B2(G1384), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n478), .A2(G40), .A3(new_n489), .A4(new_n482), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n700), .A2(G1996), .ZN(new_n919));
  INV_X1    g494(.A(G2067), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n744), .B(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n700), .A2(G1996), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n918), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n783), .B(new_n787), .Z(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(G290), .B(G1986), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n927), .B1(new_n918), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G1384), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n525), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n917), .B1(new_n931), .B2(KEYINPUT50), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT50), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n839), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  AOI21_X1  g509(.A(G1961), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G40), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n483), .A2(KEYINPUT123), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT123), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n478), .A2(new_n938), .A3(new_n482), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n916), .A2(new_n489), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT124), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n839), .A2(KEYINPUT45), .A3(new_n930), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT53), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n945), .A2(G2078), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n916), .A2(KEYINPUT124), .A3(new_n940), .A4(new_n489), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n943), .A2(new_n944), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT125), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n935), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n931), .A2(new_n911), .ZN(new_n952));
  INV_X1    g527(.A(new_n917), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n944), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G2078), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT53), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n948), .B2(KEYINPUT125), .ZN(new_n957));
  AOI21_X1  g532(.A(G301), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n944), .A2(new_n952), .A3(new_n953), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n945), .B1(new_n959), .B2(G2078), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n518), .A2(KEYINPUT72), .A3(new_n519), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n522), .B1(new_n521), .B2(new_n523), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n963), .B2(new_n514), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n917), .B1(new_n964), .B2(KEYINPUT45), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n916), .A2(new_n965), .A3(new_n946), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n966), .A2(new_n935), .A3(KEYINPUT121), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT121), .ZN(new_n968));
  INV_X1    g543(.A(G1961), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n915), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n953), .B1(new_n964), .B2(new_n933), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n916), .A2(new_n965), .A3(new_n946), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(G301), .B(new_n960), .C1(new_n967), .C2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT126), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT121), .B1(new_n966), .B2(new_n935), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n972), .A2(new_n968), .A3(new_n973), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n956), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n980), .A2(KEYINPUT126), .A3(G301), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT54), .B1(new_n958), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n951), .A2(G301), .A3(new_n957), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n960), .B1(new_n967), .B2(new_n974), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(KEYINPUT122), .A3(G171), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT122), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n988), .B1(new_n980), .B2(G301), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n984), .A2(new_n985), .A3(new_n987), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n983), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n839), .A2(new_n953), .A3(new_n930), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n592), .A2(G1976), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n992), .A2(G8), .A3(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n592), .A2(G1976), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n994), .A2(KEYINPUT52), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n994), .B2(KEYINPUT52), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NOR4_X1   g574(.A1(new_n994), .A2(new_n997), .A3(KEYINPUT52), .A4(new_n995), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(G303), .A2(G8), .ZN(new_n1002));
  XOR2_X1   g577(.A(new_n1002), .B(KEYINPUT55), .Z(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n953), .B1(new_n931), .B2(KEYINPUT50), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n933), .B1(new_n839), .B2(new_n930), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT113), .B(G2090), .Z(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1007), .A2(new_n1009), .B1(new_n959), .B2(new_n758), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1004), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n932), .A2(new_n1009), .A3(new_n934), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n954), .B2(G1971), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(G8), .A3(new_n1003), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n992), .A2(G8), .ZN(new_n1016));
  XNOR2_X1  g591(.A(G305), .B(G1981), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT49), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1001), .A2(new_n1012), .A3(new_n1015), .A4(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(G1348), .B1(new_n932), .B2(new_n934), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT60), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n992), .A2(G2067), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT119), .B1(new_n1026), .B2(new_n626), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1026), .A2(KEYINPUT118), .A3(new_n626), .ZN(new_n1028));
  INV_X1    g603(.A(G1348), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n970), .B2(new_n971), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1025), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(KEYINPUT60), .A4(new_n626), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1031), .A3(KEYINPUT60), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n617), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1027), .A2(new_n1028), .A3(new_n1034), .A4(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1024), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n725), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1041));
  XOR2_X1   g616(.A(G299), .B(KEYINPUT57), .Z(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT56), .B(G2072), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n944), .A2(new_n952), .A3(new_n953), .A4(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT61), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1041), .A2(KEYINPUT117), .A3(new_n1042), .A4(new_n1044), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1041), .A2(new_n1044), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1042), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(KEYINPUT61), .A3(new_n1045), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT58), .B(G1341), .Z(new_n1056));
  NAND2_X1  g631(.A1(new_n992), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n959), .B2(G1996), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n569), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n1059), .B(KEYINPUT59), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1040), .A2(new_n1055), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n617), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1053), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1022), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n970), .A2(new_n971), .A3(G2084), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1966), .B1(new_n916), .B2(new_n965), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G286), .A2(G8), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(KEYINPUT51), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  INV_X1    g647(.A(G1966), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n953), .B1(new_n931), .B2(new_n911), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT45), .B1(new_n839), .B2(new_n930), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1073), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n932), .A2(new_n732), .A3(new_n934), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1072), .B(G8), .C1(new_n1078), .C2(G286), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1070), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  AOI211_X1 g657(.A(KEYINPUT120), .B(new_n1070), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1071), .B(new_n1079), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n991), .A2(new_n1066), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT63), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1078), .A2(G8), .A3(G168), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1022), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1000), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(new_n1021), .C1(new_n998), .C2(new_n996), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1003), .B1(new_n1014), .B2(G8), .ZN(new_n1094));
  OR3_X1    g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1015), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1096), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1093), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1095), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT115), .B(new_n1086), .C1(new_n1022), .C2(new_n1087), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1090), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1084), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1022), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n987), .A2(new_n989), .B1(new_n1084), .B2(KEYINPUT62), .ZN(new_n1105));
  INV_X1    g680(.A(G1976), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1021), .A2(new_n1106), .A3(new_n592), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(G1981), .B2(G305), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1104), .A2(new_n1105), .B1(new_n1016), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1001), .A2(new_n1096), .A3(new_n1021), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1101), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n929), .B1(new_n1085), .B2(new_n1111), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n925), .A2(G1986), .A3(G290), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(KEYINPUT48), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n927), .B(KEYINPUT127), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT46), .ZN(new_n1117));
  OR3_X1    g692(.A1(new_n925), .A2(new_n1117), .A3(G1996), .ZN(new_n1118));
  INV_X1    g693(.A(new_n921), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n918), .B1(new_n700), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1117), .B1(new_n925), .B2(G1996), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  XOR2_X1   g697(.A(new_n1122), .B(KEYINPUT47), .Z(new_n1123));
  NAND3_X1  g698(.A1(new_n924), .A2(new_n787), .A3(new_n784), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(G2067), .B2(new_n744), .ZN(new_n1125));
  AOI211_X1 g700(.A(new_n1116), .B(new_n1123), .C1(new_n918), .C2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1112), .A2(new_n1126), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g702(.A1(G401), .A2(G227), .ZN(new_n1129));
  INV_X1    g703(.A(G319), .ZN(new_n1130));
  AOI211_X1 g704(.A(new_n1130), .B(G229), .C1(new_n906), .C2(new_n908), .ZN(new_n1131));
  NAND3_X1  g705(.A1(new_n860), .A2(new_n1129), .A3(new_n1131), .ZN(G225));
  INV_X1    g706(.A(G225), .ZN(G308));
endmodule


