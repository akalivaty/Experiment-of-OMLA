//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT84), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT85), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n190), .A2(G952), .ZN(new_n191));
  INV_X1    g005(.A(G234), .ZN(new_n192));
  INV_X1    g006(.A(G237), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n191), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G902), .ZN(new_n196));
  AOI211_X1 g010(.A(new_n196), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT21), .B(G898), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n195), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(G210), .B1(G237), .B2(G902), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G224), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(G953), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT7), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G125), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  OAI22_X1  g027(.A1(new_n209), .A2(new_n211), .B1(new_n213), .B2(G128), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  AOI21_X1  g030(.A(KEYINPUT66), .B1(new_n216), .B2(new_n209), .ZN(new_n217));
  AND4_X1   g031(.A1(KEYINPUT66), .A2(new_n209), .A3(new_n211), .A4(new_n213), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n207), .B(new_n215), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT90), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n211), .A2(new_n213), .ZN(new_n221));
  NAND2_X1  g035(.A1(KEYINPUT0), .A2(G128), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(KEYINPUT0), .B2(G128), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT0), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(new_n208), .A3(KEYINPUT65), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n221), .A2(new_n222), .A3(new_n224), .A4(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n222), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n216), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n219), .A2(new_n220), .B1(G125), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n209), .A2(new_n211), .A3(new_n213), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n216), .A2(KEYINPUT66), .A3(new_n209), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n214), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT90), .A3(new_n207), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n206), .B1(new_n231), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT91), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT89), .ZN(new_n241));
  XNOR2_X1  g055(.A(G110), .B(G122), .ZN(new_n242));
  XOR2_X1   g056(.A(new_n242), .B(KEYINPUT8), .Z(new_n243));
  INV_X1    g057(.A(G113), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT86), .A2(KEYINPUT5), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT86), .A2(KEYINPUT5), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G119), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n244), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT68), .B1(new_n248), .B2(G119), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n252));
  INV_X1    g066(.A(G119), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G116), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n248), .A2(G119), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n251), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n250), .B1(new_n256), .B2(new_n247), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT2), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n258), .A2(G113), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n244), .A2(KEYINPUT2), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n255), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n251), .A2(new_n254), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT69), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n251), .A2(new_n254), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n244), .A2(KEYINPUT2), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n258), .A2(G113), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n266), .A2(new_n267), .B1(new_n248), .B2(G119), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n264), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n257), .B1(new_n263), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT81), .ZN(new_n271));
  INV_X1    g085(.A(G107), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G104), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n271), .A2(new_n272), .A3(KEYINPUT3), .A4(G104), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G104), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G107), .ZN(new_n279));
  INV_X1    g093(.A(G101), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n272), .A2(G104), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n280), .B1(new_n284), .B2(new_n279), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n270), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n285), .B1(new_n277), .B2(new_n282), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n251), .A2(new_n254), .A3(KEYINPUT5), .A4(new_n255), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n250), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n289), .B(new_n291), .C1(new_n263), .C2(new_n269), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n241), .B(new_n243), .C1(new_n288), .C2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT69), .B1(new_n261), .B2(new_n262), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n265), .A2(new_n264), .A3(new_n268), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n245), .A2(new_n246), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n296), .A2(new_n255), .A3(new_n251), .A4(new_n254), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n294), .A2(new_n295), .B1(new_n297), .B2(new_n250), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n292), .B1(new_n289), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n243), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT89), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n240), .B1(new_n293), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n294), .A2(new_n295), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n257), .A3(new_n289), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n278), .A2(G107), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT3), .B1(new_n305), .B2(new_n271), .ZN(new_n306));
  INV_X1    g120(.A(new_n276), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n279), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT4), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(new_n309), .A3(G101), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n283), .A2(KEYINPUT4), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n280), .B1(new_n277), .B2(new_n279), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n259), .A2(new_n260), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n294), .A2(new_n295), .B1(new_n256), .B2(new_n314), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n304), .B(new_n242), .C1(new_n313), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n230), .A2(G125), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT88), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n317), .A2(new_n318), .B1(new_n207), .B2(new_n236), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n230), .A2(KEYINPUT88), .A3(G125), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(new_n206), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n316), .B(new_n321), .C1(new_n238), .C2(new_n239), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n196), .B1(new_n302), .B2(new_n322), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n319), .A2(new_n204), .A3(new_n320), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n204), .B1(new_n319), .B2(new_n320), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n316), .A2(KEYINPUT6), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n304), .B1(new_n313), .B2(new_n315), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n242), .A2(KEYINPUT87), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(KEYINPUT6), .A3(new_n329), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n326), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n201), .B1(new_n323), .B2(new_n333), .ZN(new_n334));
  AOI211_X1 g148(.A(KEYINPUT91), .B(new_n206), .C1(new_n231), .C2(new_n237), .ZN(new_n335));
  INV_X1    g149(.A(new_n292), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n289), .B1(new_n303), .B2(new_n257), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n300), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n241), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n299), .A2(KEYINPUT89), .A3(new_n300), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n335), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n322), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n316), .A2(KEYINPUT6), .B1(new_n328), .B2(new_n329), .ZN(new_n344));
  INV_X1    g158(.A(new_n332), .ZN(new_n345));
  OAI22_X1  g159(.A1(new_n344), .A2(new_n345), .B1(new_n325), .B2(new_n324), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n343), .A2(new_n346), .A3(new_n196), .A4(new_n200), .ZN(new_n347));
  AOI211_X1 g161(.A(new_n189), .B(new_n199), .C1(new_n334), .C2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT9), .B(G234), .ZN(new_n350));
  OAI21_X1  g164(.A(G221), .B1(new_n350), .B2(G902), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n351), .B(KEYINPUT78), .Z(new_n352));
  INV_X1    g166(.A(G469), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n353), .A2(new_n196), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n190), .A2(G227), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT79), .ZN(new_n356));
  XNOR2_X1  g170(.A(G110), .B(G140), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT11), .ZN(new_n360));
  INV_X1    g174(.A(G134), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n360), .B1(new_n361), .B2(G137), .ZN(new_n362));
  INV_X1    g176(.A(G137), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT11), .A3(G134), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n361), .A2(G137), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G131), .ZN(new_n367));
  INV_X1    g181(.A(G131), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n362), .A2(new_n364), .A3(new_n368), .A4(new_n365), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n371));
  NOR3_X1   g185(.A1(new_n287), .A2(new_n236), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n215), .B1(new_n217), .B2(new_n218), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT10), .B1(new_n373), .B2(new_n289), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n228), .A2(new_n211), .A3(new_n213), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n216), .A2(new_n228), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n226), .A2(new_n224), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n310), .B(new_n379), .C1(new_n311), .C2(new_n312), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n370), .B1(new_n375), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n371), .B1(new_n287), .B2(new_n236), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n373), .A2(KEYINPUT10), .A3(new_n289), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n380), .A2(new_n382), .A3(new_n370), .A4(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n359), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n373), .A2(new_n289), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n234), .A2(new_n235), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n281), .B1(new_n275), .B2(new_n276), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n388), .B(new_n215), .C1(new_n389), .C2(new_n285), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n367), .A2(new_n369), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(KEYINPUT12), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n370), .B1(new_n387), .B2(new_n390), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n384), .A3(new_n358), .ZN(new_n400));
  AOI21_X1  g214(.A(G902), .B1(new_n386), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n354), .B1(new_n401), .B2(new_n353), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT83), .ZN(new_n403));
  XOR2_X1   g217(.A(new_n358), .B(KEYINPUT80), .Z(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n399), .B2(new_n384), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n384), .A2(new_n358), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n381), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n403), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n398), .B1(new_n391), .B2(new_n392), .ZN(new_n409));
  AOI211_X1 g223(.A(new_n370), .B(new_n394), .C1(new_n387), .C2(new_n390), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n384), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n404), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n384), .A2(new_n358), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n392), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n413), .A2(KEYINPUT83), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n408), .A2(new_n418), .A3(G469), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n352), .B1(new_n402), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n193), .A2(new_n190), .A3(G214), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(new_n210), .ZN(new_n423));
  NOR2_X1   g237(.A1(G237), .A2(G953), .ZN(new_n424));
  AOI21_X1  g238(.A(G143), .B1(new_n424), .B2(G214), .ZN(new_n425));
  OAI21_X1  g239(.A(G131), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT93), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n210), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n424), .A2(G143), .A3(G214), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT93), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n431), .A3(G131), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT17), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT97), .ZN(new_n435));
  INV_X1    g249(.A(G140), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G125), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n207), .A2(G140), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT16), .ZN(new_n439));
  OR3_X1    g253(.A1(new_n207), .A2(KEYINPUT16), .A3(G140), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(G146), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(G146), .B1(new_n439), .B2(new_n440), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n435), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n439), .A2(new_n440), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n212), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT97), .A3(new_n441), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n423), .A2(new_n425), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n368), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT17), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n427), .A2(new_n450), .A3(new_n451), .A4(new_n432), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n434), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT18), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n449), .B1(new_n454), .B2(new_n368), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n430), .A2(KEYINPUT18), .A3(G131), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n437), .A2(new_n438), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G146), .ZN(new_n458));
  XNOR2_X1  g272(.A(G125), .B(G140), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n212), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n458), .A2(new_n460), .A3(KEYINPUT92), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT92), .B1(new_n458), .B2(new_n460), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n455), .B(new_n456), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n453), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G113), .B(G122), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT96), .B(G104), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n453), .A2(new_n463), .A3(new_n467), .ZN(new_n470));
  AOI21_X1  g284(.A(G902), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G475), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT20), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n427), .A2(new_n450), .A3(new_n432), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT95), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(new_n459), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT95), .B1(new_n457), .B2(new_n476), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n457), .A2(KEYINPUT19), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n212), .A4(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT74), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n441), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n439), .A2(new_n440), .A3(KEYINPUT74), .A4(G146), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n463), .B1(new_n475), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n468), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n470), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(G475), .A2(G902), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n474), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n474), .A3(new_n490), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(KEYINPUT98), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT98), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n489), .A2(new_n494), .A3(new_n474), .A4(new_n490), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n473), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G122), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(G116), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n248), .A2(G122), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT99), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(G116), .B(G122), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(KEYINPUT99), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n272), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n501), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(KEYINPUT99), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n507), .A3(G107), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n208), .A2(G143), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT13), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n210), .A2(G128), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT100), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(new_n512), .B2(new_n511), .ZN(new_n514));
  AOI211_X1 g328(.A(KEYINPUT100), .B(KEYINPUT13), .C1(new_n210), .C2(G128), .ZN(new_n515));
  OAI221_X1 g329(.A(new_n510), .B1(new_n511), .B2(new_n512), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G134), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n510), .A3(new_n361), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n509), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n505), .A2(KEYINPUT101), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT101), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n521), .B(new_n272), .C1(new_n502), .C2(new_n504), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n500), .A2(KEYINPUT14), .ZN(new_n523));
  INV_X1    g337(.A(new_n499), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n272), .B1(new_n524), .B2(KEYINPUT14), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n512), .A2(new_n510), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G134), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n523), .A2(new_n525), .B1(new_n527), .B2(new_n518), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n520), .A2(new_n522), .A3(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G217), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n350), .A2(new_n530), .A3(G953), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n519), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(new_n519), .B2(new_n529), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n196), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT15), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n535), .A3(G478), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(G478), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n196), .B(new_n537), .C1(new_n532), .C2(new_n533), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n496), .A2(new_n539), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n349), .A2(new_n421), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n530), .B1(G234), .B2(new_n196), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n196), .A2(KEYINPUT25), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT24), .B(G110), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n253), .A2(G128), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n208), .A2(G119), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT73), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n545), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT23), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n253), .B2(G128), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n208), .A2(KEYINPUT23), .A3(G119), .ZN(new_n555));
  INV_X1    g369(.A(G110), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .A4(new_n546), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n460), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n484), .A2(new_n485), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT75), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n460), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n546), .A2(new_n547), .A3(new_n550), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n550), .B1(new_n546), .B2(new_n547), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n544), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n562), .B1(new_n565), .B2(new_n557), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT75), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n484), .A4(new_n485), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n442), .A2(new_n443), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n549), .A2(new_n551), .A3(new_n545), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n554), .A2(new_n546), .A3(new_n555), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G110), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT22), .B(G137), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n543), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n575), .B1(new_n561), .B2(new_n568), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n583), .A2(KEYINPUT76), .A3(new_n580), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT76), .B1(new_n583), .B2(new_n580), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT77), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT77), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n582), .B(new_n588), .C1(new_n584), .C2(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n583), .A2(new_n580), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT76), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n577), .B2(new_n581), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n583), .A2(KEYINPUT76), .A3(new_n580), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT25), .B1(new_n595), .B2(new_n196), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n542), .B1(new_n590), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n542), .A2(G902), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(G472), .A2(G902), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT31), .ZN(new_n602));
  INV_X1    g416(.A(new_n365), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n361), .A2(G137), .ZN(new_n604));
  OAI21_X1  g418(.A(G131), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n369), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n373), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n379), .A2(new_n392), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n608), .A2(new_n315), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT26), .B(G101), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n424), .A2(G210), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n373), .A2(new_n607), .B1(new_n379), .B2(new_n392), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n315), .B1(new_n617), .B2(KEYINPUT30), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT67), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  OAI22_X1  g435(.A1(new_n370), .A2(new_n230), .B1(new_n236), .B2(new_n606), .ZN(new_n622));
  INV_X1    g436(.A(new_n620), .ZN(new_n623));
  AOI21_X1  g437(.A(KEYINPUT67), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI211_X1 g438(.A(KEYINPUT70), .B(new_n618), .C1(new_n621), .C2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n619), .B1(new_n617), .B2(new_n620), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n622), .A2(KEYINPUT67), .A3(new_n623), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT70), .B1(new_n629), .B2(new_n618), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n602), .B(new_n616), .C1(new_n626), .C2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n615), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n315), .B1(new_n608), .B2(new_n609), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT28), .B1(new_n610), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(KEYINPUT28), .B1(new_n617), .B2(new_n315), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n632), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n618), .B1(new_n621), .B2(new_n624), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT70), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n625), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n602), .B1(new_n643), .B2(new_n616), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n601), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT32), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n634), .A2(new_n632), .A3(new_n636), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT29), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n610), .B1(new_n642), .B2(new_n625), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n651), .B1(new_n652), .B2(new_n632), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT28), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n256), .A2(new_n314), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n303), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n622), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n608), .A2(new_n315), .A3(new_n609), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n659), .A2(new_n615), .A3(new_n635), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT72), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n661), .A3(KEYINPUT29), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n634), .A2(KEYINPUT29), .A3(new_n632), .A4(new_n636), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT72), .ZN(new_n664));
  AOI21_X1  g478(.A(G902), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n653), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n616), .B1(new_n626), .B2(new_n630), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT31), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(new_n638), .A3(new_n631), .ZN(new_n669));
  INV_X1    g483(.A(new_n601), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n646), .ZN(new_n671));
  AOI22_X1  g485(.A1(G472), .A2(new_n666), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n600), .B1(new_n647), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n541), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G101), .ZN(G3));
  INV_X1    g489(.A(new_n616), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n676), .B1(new_n642), .B2(new_n625), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n637), .B1(new_n677), .B2(new_n602), .ZN(new_n678));
  AOI21_X1  g492(.A(G902), .B1(new_n678), .B2(new_n668), .ZN(new_n679));
  INV_X1    g493(.A(G472), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n645), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n600), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n420), .ZN(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT102), .Z(new_n684));
  OAI21_X1  g498(.A(KEYINPUT33), .B1(new_n532), .B2(new_n533), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n519), .A2(new_n529), .ZN(new_n686));
  INV_X1    g500(.A(new_n531), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT33), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n519), .A2(new_n529), .A3(new_n531), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n685), .A2(new_n691), .A3(G478), .ZN(new_n692));
  NAND2_X1  g506(.A1(G478), .A2(G902), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n692), .B(new_n693), .C1(G478), .C2(new_n534), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n492), .A2(KEYINPUT98), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n489), .A2(new_n490), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(KEYINPUT20), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n695), .A2(new_n495), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n473), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n694), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n199), .B1(new_n334), .B2(new_n347), .ZN(new_n701));
  INV_X1    g515(.A(new_n188), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n684), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT103), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT34), .B(G104), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G6));
  AND3_X1   g521(.A1(new_n489), .A2(new_n474), .A3(new_n490), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n491), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n709), .A2(new_n539), .A3(new_n473), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n701), .A2(new_n710), .A3(new_n702), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n684), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT104), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT35), .B(G107), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G9));
  INV_X1    g529(.A(KEYINPUT25), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n577), .A2(new_n581), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n717), .B1(new_n584), .B2(new_n585), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n716), .B1(new_n718), .B2(G902), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n587), .A3(new_n589), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n577), .B(KEYINPUT105), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n581), .A2(KEYINPUT36), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n720), .A2(new_n542), .B1(new_n723), .B2(new_n598), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n681), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n541), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT37), .B(G110), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G12));
  AOI21_X1  g542(.A(new_n724), .B1(new_n672), .B2(new_n647), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n188), .B1(new_n334), .B2(new_n347), .ZN(new_n730));
  INV_X1    g544(.A(G900), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n197), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n194), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(new_n471), .B2(new_n472), .ZN(new_n734));
  NOR3_X1   g548(.A1(new_n709), .A2(new_n539), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n420), .A2(new_n730), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT106), .B1(new_n729), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n658), .B1(new_n626), .B2(new_n630), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n650), .B1(new_n738), .B2(new_n615), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n661), .B1(new_n660), .B2(KEYINPUT29), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n663), .A2(KEYINPUT72), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n196), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(G472), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n671), .B1(new_n639), .B2(new_n644), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n670), .B1(new_n678), .B2(new_n668), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n743), .B(new_n744), .C1(new_n745), .C2(KEYINPUT32), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n723), .A2(new_n598), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n597), .A2(new_n747), .ZN(new_n748));
  AND4_X1   g562(.A1(KEYINPUT106), .A2(new_n736), .A3(new_n746), .A4(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n737), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G128), .ZN(G30));
  NAND2_X1  g565(.A1(new_n334), .A2(new_n347), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT38), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n536), .A2(new_n538), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n698), .A2(new_n699), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n756), .A2(new_n188), .A3(new_n748), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n733), .B(KEYINPUT39), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n420), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n759), .B(KEYINPUT40), .Z(new_n760));
  NOR2_X1   g574(.A1(new_n652), .A2(new_n615), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n657), .A2(new_n658), .A3(new_n615), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n196), .ZN(new_n763));
  OAI21_X1  g577(.A(G472), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n744), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n647), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n757), .A2(new_n760), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G143), .ZN(G45));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n700), .A2(new_n733), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n769), .B1(new_n771), .B2(new_n730), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n700), .A2(new_n730), .A3(new_n769), .A4(new_n733), .ZN(new_n774));
  AND4_X1   g588(.A1(new_n746), .A2(new_n774), .A3(new_n420), .A4(new_n748), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G146), .ZN(G48));
  AOI21_X1  g591(.A(new_n358), .B1(new_n416), .B2(new_n384), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(new_n414), .B2(new_n399), .ZN(new_n779));
  OAI21_X1  g593(.A(G469), .B1(new_n779), .B2(G902), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n401), .A2(new_n353), .ZN(new_n781));
  INV_X1    g595(.A(new_n352), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n673), .A2(new_n703), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT41), .B(G113), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT108), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n784), .B(new_n786), .ZN(G15));
  AOI22_X1  g601(.A1(new_n720), .A2(new_n542), .B1(new_n595), .B2(new_n598), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n746), .A2(new_n711), .A3(new_n788), .A4(new_n783), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G116), .ZN(G18));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n323), .A2(new_n201), .A3(new_n333), .ZN(new_n792));
  AOI21_X1  g606(.A(G902), .B1(new_n341), .B2(new_n342), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n200), .B1(new_n793), .B2(new_n346), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n702), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n783), .A2(new_n730), .A3(KEYINPUT109), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n540), .ZN(new_n800));
  INV_X1    g614(.A(new_n199), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n729), .A2(new_n799), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G119), .ZN(G21));
  NOR3_X1   g617(.A1(new_n795), .A2(new_n539), .A3(new_n496), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n682), .A2(new_n801), .A3(new_n783), .A4(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G122), .ZN(G24));
  OAI21_X1  g620(.A(KEYINPUT110), .B1(new_n681), .B2(new_n724), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n196), .B1(new_n639), .B2(new_n644), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(G472), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n748), .A2(new_n808), .A3(new_n645), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n807), .A2(new_n799), .A3(new_n811), .A4(new_n771), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G125), .ZN(G27));
  INV_X1    g627(.A(KEYINPUT42), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n746), .A2(new_n788), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n334), .A2(new_n347), .A3(new_n702), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n413), .A2(G469), .A3(new_n417), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n352), .B1(new_n402), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n817), .A2(new_n700), .A3(new_n733), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n814), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n820), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n673), .A2(KEYINPUT42), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G131), .ZN(G33));
  AND3_X1   g639(.A1(new_n817), .A2(new_n735), .A3(new_n819), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n673), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(G134), .ZN(G36));
  INV_X1    g642(.A(KEYINPUT43), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n693), .B1(new_n534), .B2(G478), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n685), .A2(new_n691), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(G478), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n829), .B1(new_n496), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n698), .A2(new_n832), .A3(new_n699), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(KEYINPUT43), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT112), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n810), .A2(new_n645), .B1(new_n597), .B2(new_n747), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n496), .A2(new_n829), .A3(new_n832), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n834), .A2(KEYINPUT43), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n836), .A2(new_n837), .A3(KEYINPUT44), .A4(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT113), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n836), .A2(new_n841), .A3(new_n837), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT44), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n354), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT45), .B1(new_n408), .B2(new_n418), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n413), .A2(KEYINPUT45), .A3(new_n417), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(G469), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n847), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT46), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(KEYINPUT46), .B(new_n847), .C1(new_n848), .C2(new_n850), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n781), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n782), .A3(new_n758), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT111), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT111), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n855), .A2(new_n858), .A3(new_n782), .A4(new_n758), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n843), .A2(new_n817), .A3(new_n846), .A4(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(G137), .ZN(G39));
  NAND2_X1  g676(.A1(new_n855), .A2(new_n782), .ZN(new_n863));
  XNOR2_X1  g677(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n855), .A2(new_n782), .A3(new_n864), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OR4_X1    g682(.A1(new_n746), .A2(new_n788), .A3(new_n770), .A4(new_n816), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(new_n436), .ZN(G42));
  NAND3_X1  g685(.A1(new_n838), .A2(new_n839), .A3(new_n195), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT121), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n753), .A2(new_n702), .A3(new_n796), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n682), .A3(new_n874), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n875), .B(KEYINPUT50), .Z(new_n876));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n817), .A2(new_n783), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n873), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n877), .B1(new_n873), .B2(new_n879), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n807), .B(new_n811), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n780), .A2(new_n781), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n868), .B1(new_n782), .B2(new_n883), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n873), .A2(new_n682), .A3(new_n817), .ZN(new_n885));
  INV_X1    g699(.A(new_n766), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n886), .A2(new_n788), .A3(new_n195), .A4(new_n879), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n755), .A2(new_n832), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  OR3_X1    g703(.A1(new_n887), .A2(KEYINPUT123), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT123), .B1(new_n887), .B2(new_n889), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n884), .A2(new_n885), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n876), .A2(new_n882), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT51), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n873), .A2(new_n682), .A3(new_n799), .ZN(new_n897));
  INV_X1    g711(.A(new_n700), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n897), .B(new_n191), .C1(new_n887), .C2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n673), .B1(new_n880), .B2(new_n881), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n900), .A2(KEYINPUT48), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(KEYINPUT48), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n895), .A2(new_n896), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n812), .B1(new_n737), .B2(new_n749), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT118), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n733), .B(KEYINPUT119), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n724), .A2(new_n819), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(new_n766), .A3(new_n804), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT118), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n812), .B(new_n911), .C1(new_n737), .C2(new_n749), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n906), .A2(new_n776), .A3(new_n910), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT52), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n776), .A2(new_n910), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT52), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n917), .A2(new_n750), .A3(new_n918), .A4(new_n812), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n802), .A2(new_n784), .A3(new_n805), .A4(new_n789), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n821), .A2(new_n823), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n189), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT115), .A4(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT116), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n754), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n536), .A2(KEYINPUT116), .A3(new_n538), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n929), .A2(new_n701), .A3(new_n496), .A4(new_n923), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n924), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT115), .B1(new_n348), .B2(new_n700), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n682), .B(new_n420), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(new_n674), .A3(new_n726), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT117), .ZN(new_n935));
  INV_X1    g749(.A(new_n709), .ZN(new_n936));
  INV_X1    g750(.A(new_n734), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n935), .B1(new_n929), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n928), .A2(KEYINPUT117), .A3(new_n936), .A4(new_n937), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n940), .A2(new_n817), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n729), .A2(new_n420), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n807), .A2(new_n811), .A3(new_n822), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n943), .A3(new_n827), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n934), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n922), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n914), .A2(new_n915), .A3(new_n919), .A4(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT52), .B1(new_n916), .B2(new_n905), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n919), .A2(new_n922), .A3(new_n945), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(KEYINPUT53), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n947), .A2(new_n950), .A3(KEYINPUT54), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n934), .A2(new_n944), .A3(new_n915), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT120), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n920), .B2(new_n921), .ZN(new_n954));
  INV_X1    g768(.A(new_n799), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n746), .A2(new_n800), .A3(new_n801), .A4(new_n748), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n789), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n784), .A2(new_n805), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n958), .A2(new_n959), .A3(KEYINPUT120), .A4(new_n824), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n952), .A2(new_n954), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n961), .A2(new_n914), .A3(new_n919), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n949), .A2(new_n915), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n951), .B1(new_n964), .B2(KEYINPUT54), .ZN(new_n965));
  OAI22_X1  g779(.A1(new_n904), .A2(new_n965), .B1(G952), .B2(G953), .ZN(new_n966));
  AOI211_X1 g780(.A(new_n189), .B(new_n352), .C1(new_n883), .C2(KEYINPUT49), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(KEYINPUT49), .B2(new_n883), .ZN(new_n968));
  OR4_X1    g782(.A1(new_n600), .A2(new_n968), .A3(new_n753), .A4(new_n834), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n966), .B1(new_n766), .B2(new_n969), .ZN(G75));
  NOR2_X1   g784(.A1(new_n344), .A2(new_n345), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n326), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n346), .ZN(new_n973));
  XNOR2_X1  g787(.A(KEYINPUT124), .B(KEYINPUT55), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(G210), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n977), .B(new_n196), .C1(new_n962), .C2(new_n963), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n976), .B1(new_n978), .B2(KEYINPUT56), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT56), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n964), .A2(G902), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n980), .B(new_n975), .C1(new_n981), .C2(new_n977), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n190), .A2(G952), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n979), .A2(new_n982), .A3(new_n984), .ZN(G51));
  XNOR2_X1  g799(.A(new_n354), .B(KEYINPUT57), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT54), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n962), .A2(new_n963), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n987), .B1(new_n962), .B2(new_n963), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n986), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n779), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OR3_X1    g806(.A1(new_n981), .A2(new_n848), .A3(new_n850), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n983), .B1(new_n992), .B2(new_n993), .ZN(G54));
  AOI21_X1  g808(.A(new_n196), .B1(new_n962), .B2(new_n963), .ZN(new_n995));
  NAND2_X1  g809(.A1(KEYINPUT58), .A2(G475), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n995), .A2(new_n489), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n489), .B1(new_n995), .B2(new_n997), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n998), .A2(new_n999), .A3(new_n983), .ZN(G60));
  XNOR2_X1  g814(.A(new_n831), .B(KEYINPUT125), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n693), .B(KEYINPUT59), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n1001), .B(new_n1002), .C1(new_n988), .C2(new_n989), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n984), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1001), .B1(new_n965), .B2(new_n1002), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1004), .A2(new_n1005), .ZN(G63));
  INV_X1    g820(.A(KEYINPUT61), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G217), .A2(G902), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT60), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(new_n962), .B2(new_n963), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n723), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n984), .B1(new_n1010), .B2(new_n595), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1007), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n1010), .A2(new_n595), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n1015), .A2(KEYINPUT61), .A3(new_n984), .A4(new_n1011), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1014), .A2(new_n1016), .ZN(G66));
  OAI21_X1  g831(.A(G953), .B1(new_n198), .B2(new_n202), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n920), .A2(new_n934), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n1019), .B2(G953), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n971), .B1(G898), .B2(new_n190), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1020), .B(new_n1021), .ZN(G69));
  AOI21_X1  g836(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT127), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT30), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n629), .B1(new_n1027), .B2(new_n622), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n729), .A2(new_n420), .A3(new_n774), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1031), .A2(new_n772), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1032), .B1(new_n905), .B2(KEYINPUT118), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT62), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1033), .A2(new_n1034), .A3(new_n767), .A4(new_n912), .ZN(new_n1035));
  INV_X1    g849(.A(new_n870), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n700), .B1(new_n496), .B2(new_n929), .ZN(new_n1037));
  OR4_X1    g851(.A1(new_n815), .A2(new_n759), .A3(new_n816), .A4(new_n1037), .ZN(new_n1038));
  AND3_X1   g852(.A1(new_n861), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n906), .A2(new_n767), .A3(new_n776), .A4(new_n912), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT126), .ZN(new_n1041));
  AND3_X1   g855(.A1(new_n1040), .A2(new_n1041), .A3(KEYINPUT62), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1041), .B1(new_n1040), .B2(KEYINPUT62), .ZN(new_n1043));
  OAI211_X1 g857(.A(new_n1035), .B(new_n1039), .C1(new_n1042), .C2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1030), .B1(new_n1044), .B2(new_n190), .ZN(new_n1045));
  INV_X1    g859(.A(new_n1030), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1046), .B1(G900), .B2(G953), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n861), .A2(new_n1036), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n826), .B1(new_n860), .B2(new_n804), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n1050), .A2(new_n815), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1033), .A2(new_n824), .A3(new_n912), .ZN(new_n1052));
  NOR3_X1   g866(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1048), .B1(new_n1053), .B2(new_n190), .ZN(new_n1054));
  OAI211_X1 g868(.A(new_n1025), .B(new_n1026), .C1(new_n1045), .C2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g869(.A1(new_n1035), .A2(new_n861), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1056));
  INV_X1    g870(.A(new_n1043), .ZN(new_n1057));
  NAND3_X1  g871(.A1(new_n1040), .A2(new_n1041), .A3(KEYINPUT62), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g873(.A(new_n1046), .B1(new_n1059), .B2(G953), .ZN(new_n1060));
  INV_X1    g874(.A(new_n1054), .ZN(new_n1061));
  NAND4_X1  g875(.A1(new_n1060), .A2(new_n1024), .A3(new_n1023), .A4(new_n1061), .ZN(new_n1062));
  AND2_X1   g876(.A1(new_n1055), .A2(new_n1062), .ZN(G72));
  NAND2_X1  g877(.A1(new_n947), .A2(new_n950), .ZN(new_n1064));
  NOR2_X1   g878(.A1(new_n738), .A2(new_n632), .ZN(new_n1065));
  NAND2_X1  g879(.A1(G472), .A2(G902), .ZN(new_n1066));
  XOR2_X1   g880(.A(new_n1066), .B(KEYINPUT63), .Z(new_n1067));
  INV_X1    g881(.A(new_n1067), .ZN(new_n1068));
  OR3_X1    g882(.A1(new_n1065), .A2(new_n761), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g883(.A(new_n1068), .B1(new_n1053), .B2(new_n1019), .ZN(new_n1070));
  INV_X1    g884(.A(new_n1065), .ZN(new_n1071));
  OAI221_X1 g885(.A(new_n984), .B1(new_n1064), .B2(new_n1069), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  INV_X1    g886(.A(new_n1019), .ZN(new_n1073));
  OAI21_X1  g887(.A(new_n1067), .B1(new_n1044), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g888(.A(new_n1072), .B1(new_n761), .B2(new_n1074), .ZN(G57));
endmodule


