

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U553 ( .A1(n762), .A2(n973), .ZN(n757) );
  NOR2_X1 U554 ( .A1(n831), .A2(n830), .ZN(n839) );
  OR2_X1 U555 ( .A1(n531), .A2(G164), .ZN(n797) );
  OR2_X1 U556 ( .A1(n842), .A2(n523), .ZN(n550) );
  INV_X1 U557 ( .A(KEYINPUT40), .ZN(n546) );
  NOR2_X1 U558 ( .A1(n534), .A2(n1025), .ZN(n533) );
  INV_X1 U559 ( .A(n535), .ZN(n534) );
  NOR2_X1 U560 ( .A1(n549), .A2(KEYINPUT40), .ZN(n548) );
  NAND2_X1 U561 ( .A1(n522), .A2(n544), .ZN(n543) );
  NAND2_X1 U562 ( .A1(n858), .A2(n545), .ZN(n544) );
  NAND2_X1 U563 ( .A1(n550), .A2(n546), .ZN(n545) );
  NOR2_X1 U564 ( .A1(G164), .A2(n532), .ZN(n538) );
  NAND2_X1 U565 ( .A1(n533), .A2(n536), .ZN(n532) );
  INV_X1 U566 ( .A(KEYINPUT92), .ZN(n756) );
  NOR2_X1 U567 ( .A1(n560), .A2(n519), .ZN(n535) );
  INV_X1 U568 ( .A(n561), .ZN(n536) );
  INV_X1 U569 ( .A(G2104), .ZN(n530) );
  AND2_X1 U570 ( .A1(n553), .A2(G2104), .ZN(n923) );
  NOR2_X1 U571 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U572 ( .A(n584), .B(n583), .ZN(n679) );
  NOR2_X1 U573 ( .A1(G2104), .A2(n553), .ZN(n920) );
  NAND2_X1 U574 ( .A1(n541), .A2(n540), .ZN(n539) );
  AND2_X1 U575 ( .A1(n547), .A2(n543), .ZN(n542) );
  NOR2_X1 U576 ( .A1(n550), .A2(n546), .ZN(n540) );
  NOR2_X1 U577 ( .A1(n561), .A2(n560), .ZN(G160) );
  OR2_X1 U578 ( .A1(G1384), .A2(n749), .ZN(n519) );
  NAND2_X1 U579 ( .A1(n771), .A2(n770), .ZN(n520) );
  NAND2_X1 U580 ( .A1(G160), .A2(G40), .ZN(n521) );
  OR2_X1 U581 ( .A1(n858), .A2(KEYINPUT40), .ZN(n522) );
  AND2_X1 U582 ( .A1(n975), .A2(n856), .ZN(n523) );
  XNOR2_X1 U583 ( .A(n524), .B(n774), .ZN(n779) );
  NAND2_X1 U584 ( .A1(n525), .A2(n773), .ZN(n524) );
  NAND2_X1 U585 ( .A1(n526), .A2(n520), .ZN(n525) );
  XNOR2_X1 U586 ( .A(n765), .B(n527), .ZN(n526) );
  INV_X1 U587 ( .A(KEYINPUT93), .ZN(n527) );
  NAND2_X1 U588 ( .A1(n573), .A2(n528), .ZN(n574) );
  NAND2_X1 U589 ( .A1(n925), .A2(G138), .ZN(n528) );
  XNOR2_X2 U590 ( .A(n529), .B(KEYINPUT17), .ZN(n925) );
  NAND2_X1 U591 ( .A1(n553), .A2(n530), .ZN(n529) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n531) );
  XNOR2_X1 U593 ( .A(n538), .B(n537), .ZN(n752) );
  INV_X1 U594 ( .A(KEYINPUT26), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n542), .A2(n539), .ZN(G329) );
  INV_X1 U596 ( .A(n841), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n841), .A2(n548), .ZN(n547) );
  INV_X1 U598 ( .A(n858), .ZN(n549) );
  INV_X1 U599 ( .A(KEYINPUT64), .ZN(n754) );
  NAND2_X1 U600 ( .A1(n679), .A2(G81), .ZN(n617) );
  XNOR2_X1 U601 ( .A(KEYINPUT73), .B(KEYINPUT13), .ZN(n621) );
  XNOR2_X1 U602 ( .A(n622), .B(n621), .ZN(n623) );
  INV_X1 U603 ( .A(KEYINPUT65), .ZN(n583) );
  NOR2_X1 U604 ( .A1(G651), .A2(n691), .ZN(n686) );
  NAND2_X1 U605 ( .A1(G137), .A2(n925), .ZN(n551) );
  XNOR2_X1 U606 ( .A(n551), .B(KEYINPUT68), .ZN(n557) );
  INV_X1 U607 ( .A(G2105), .ZN(n553) );
  NAND2_X1 U608 ( .A1(G101), .A2(n923), .ZN(n552) );
  XOR2_X1 U609 ( .A(KEYINPUT23), .B(n552), .Z(n555) );
  NAND2_X1 U610 ( .A1(n920), .A2(G125), .ZN(n554) );
  AND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U613 ( .A1(G2104), .A2(G2105), .ZN(n558) );
  XOR2_X1 U614 ( .A(KEYINPUT66), .B(n558), .Z(n575) );
  BUF_X1 U615 ( .A(n575), .Z(n905) );
  NAND2_X1 U616 ( .A1(G113), .A2(n905), .ZN(n559) );
  XNOR2_X1 U617 ( .A(KEYINPUT67), .B(n559), .ZN(n560) );
  XNOR2_X1 U618 ( .A(G2451), .B(G2443), .ZN(n571) );
  XOR2_X1 U619 ( .A(G2446), .B(G2454), .Z(n563) );
  XNOR2_X1 U620 ( .A(KEYINPUT105), .B(G2435), .ZN(n562) );
  XNOR2_X1 U621 ( .A(n563), .B(n562), .ZN(n567) );
  XOR2_X1 U622 ( .A(KEYINPUT106), .B(G2438), .Z(n565) );
  XNOR2_X1 U623 ( .A(G1341), .B(G1348), .ZN(n564) );
  XNOR2_X1 U624 ( .A(n565), .B(n564), .ZN(n566) );
  XOR2_X1 U625 ( .A(n567), .B(n566), .Z(n569) );
  XNOR2_X1 U626 ( .A(G2430), .B(G2427), .ZN(n568) );
  XNOR2_X1 U627 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U628 ( .A(n571), .B(n570), .ZN(n572) );
  AND2_X1 U629 ( .A1(n572), .A2(G14), .ZN(G401) );
  NAND2_X1 U630 ( .A1(G102), .A2(n923), .ZN(n573) );
  XOR2_X1 U631 ( .A(KEYINPUT86), .B(n574), .Z(n579) );
  NAND2_X1 U632 ( .A1(n920), .A2(G126), .ZN(n577) );
  NAND2_X1 U633 ( .A1(G114), .A2(n905), .ZN(n576) );
  AND2_X1 U634 ( .A1(n577), .A2(n576), .ZN(n578) );
  AND2_X1 U635 ( .A1(n579), .A2(n578), .ZN(G164) );
  XOR2_X1 U636 ( .A(G543), .B(KEYINPUT0), .Z(n691) );
  NAND2_X1 U637 ( .A1(n686), .A2(G52), .ZN(n582) );
  INV_X1 U638 ( .A(G651), .ZN(n585) );
  NOR2_X1 U639 ( .A1(G543), .A2(n585), .ZN(n580) );
  XOR2_X1 U640 ( .A(KEYINPUT1), .B(n580), .Z(n613) );
  NAND2_X1 U641 ( .A1(G64), .A2(n613), .ZN(n581) );
  AND2_X1 U642 ( .A1(n582), .A2(n581), .ZN(n591) );
  XNOR2_X1 U643 ( .A(KEYINPUT70), .B(KEYINPUT9), .ZN(n589) );
  NOR2_X1 U644 ( .A1(G651), .A2(G543), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G90), .A2(n679), .ZN(n587) );
  NOR2_X1 U646 ( .A1(n691), .A2(n585), .ZN(n618) );
  NAND2_X1 U647 ( .A1(G77), .A2(n618), .ZN(n586) );
  NAND2_X1 U648 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U649 ( .A(n589), .B(n588), .ZN(n590) );
  NAND2_X1 U650 ( .A1(n591), .A2(n590), .ZN(G301) );
  INV_X1 U651 ( .A(G301), .ZN(G171) );
  AND2_X1 U652 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U653 ( .A1(G135), .A2(n925), .ZN(n593) );
  NAND2_X1 U654 ( .A1(G111), .A2(n905), .ZN(n592) );
  NAND2_X1 U655 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U656 ( .A1(n920), .A2(G123), .ZN(n594) );
  XOR2_X1 U657 ( .A(KEYINPUT18), .B(n594), .Z(n595) );
  NOR2_X1 U658 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U659 ( .A1(n923), .A2(G99), .ZN(n597) );
  NAND2_X1 U660 ( .A1(n598), .A2(n597), .ZN(n954) );
  XNOR2_X1 U661 ( .A(G2096), .B(n954), .ZN(n599) );
  OR2_X1 U662 ( .A1(G2100), .A2(n599), .ZN(G156) );
  INV_X1 U663 ( .A(G57), .ZN(G237) );
  INV_X1 U664 ( .A(G132), .ZN(G219) );
  INV_X1 U665 ( .A(G82), .ZN(G220) );
  NAND2_X1 U666 ( .A1(n679), .A2(G89), .ZN(n600) );
  XNOR2_X1 U667 ( .A(n600), .B(KEYINPUT4), .ZN(n602) );
  NAND2_X1 U668 ( .A1(G76), .A2(n618), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U670 ( .A(n603), .B(KEYINPUT5), .ZN(n609) );
  NAND2_X1 U671 ( .A1(n686), .A2(G51), .ZN(n604) );
  XNOR2_X1 U672 ( .A(n604), .B(KEYINPUT78), .ZN(n606) );
  NAND2_X1 U673 ( .A1(G63), .A2(n613), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U675 ( .A(KEYINPUT6), .B(n607), .Z(n608) );
  NAND2_X1 U676 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U677 ( .A(n610), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U678 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U679 ( .A1(G7), .A2(G661), .ZN(n611) );
  XNOR2_X1 U680 ( .A(n611), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U681 ( .A(G223), .ZN(n859) );
  NAND2_X1 U682 ( .A1(n859), .A2(G567), .ZN(n612) );
  XOR2_X1 U683 ( .A(KEYINPUT11), .B(n612), .Z(G234) );
  XOR2_X1 U684 ( .A(G860), .B(KEYINPUT75), .Z(n650) );
  NAND2_X1 U685 ( .A1(n613), .A2(G56), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n614), .B(KEYINPUT14), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G43), .A2(n686), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n624) );
  XNOR2_X1 U689 ( .A(n617), .B(KEYINPUT12), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G68), .A2(n618), .ZN(n619) );
  NAND2_X1 U691 ( .A1(n620), .A2(n619), .ZN(n622) );
  XOR2_X2 U692 ( .A(KEYINPUT74), .B(n625), .Z(n978) );
  INV_X1 U693 ( .A(n978), .ZN(n626) );
  NAND2_X1 U694 ( .A1(n650), .A2(n626), .ZN(G153) );
  NAND2_X1 U695 ( .A1(G301), .A2(G868), .ZN(n627) );
  XNOR2_X1 U696 ( .A(n627), .B(KEYINPUT76), .ZN(n637) );
  INV_X1 U697 ( .A(G868), .ZN(n703) );
  NAND2_X1 U698 ( .A1(n618), .A2(G79), .ZN(n634) );
  NAND2_X1 U699 ( .A1(G54), .A2(n686), .ZN(n629) );
  NAND2_X1 U700 ( .A1(G66), .A2(n613), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U702 ( .A1(G92), .A2(n679), .ZN(n630) );
  XNOR2_X1 U703 ( .A(KEYINPUT77), .B(n630), .ZN(n631) );
  NOR2_X1 U704 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U706 ( .A(KEYINPUT15), .B(n635), .Z(n973) );
  NAND2_X1 U707 ( .A1(n703), .A2(n973), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n637), .A2(n636), .ZN(G284) );
  NAND2_X1 U709 ( .A1(G65), .A2(n613), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n638), .B(KEYINPUT72), .ZN(n645) );
  NAND2_X1 U711 ( .A1(G91), .A2(n679), .ZN(n640) );
  NAND2_X1 U712 ( .A1(G53), .A2(n686), .ZN(n639) );
  NAND2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U714 ( .A1(G78), .A2(n618), .ZN(n641) );
  XNOR2_X1 U715 ( .A(KEYINPUT71), .B(n641), .ZN(n642) );
  NOR2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(G299) );
  XNOR2_X1 U718 ( .A(KEYINPUT79), .B(G868), .ZN(n646) );
  NOR2_X1 U719 ( .A1(G286), .A2(n646), .ZN(n648) );
  NOR2_X1 U720 ( .A1(G868), .A2(G299), .ZN(n647) );
  NOR2_X1 U721 ( .A1(n648), .A2(n647), .ZN(G297) );
  INV_X1 U722 ( .A(G559), .ZN(n649) );
  NOR2_X1 U723 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U724 ( .A1(n973), .A2(n651), .ZN(n652) );
  XOR2_X1 U725 ( .A(KEYINPUT16), .B(n652), .Z(G148) );
  NOR2_X1 U726 ( .A1(n978), .A2(G868), .ZN(n655) );
  INV_X1 U727 ( .A(n973), .ZN(n866) );
  NAND2_X1 U728 ( .A1(G868), .A2(n866), .ZN(n653) );
  NOR2_X1 U729 ( .A1(G559), .A2(n653), .ZN(n654) );
  NOR2_X1 U730 ( .A1(n655), .A2(n654), .ZN(G282) );
  NAND2_X1 U731 ( .A1(G559), .A2(n866), .ZN(n656) );
  XNOR2_X1 U732 ( .A(n978), .B(n656), .ZN(n699) );
  NOR2_X1 U733 ( .A1(G860), .A2(n699), .ZN(n664) );
  NAND2_X1 U734 ( .A1(G55), .A2(n686), .ZN(n658) );
  NAND2_X1 U735 ( .A1(G67), .A2(n613), .ZN(n657) );
  NAND2_X1 U736 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U737 ( .A(KEYINPUT80), .B(n659), .ZN(n663) );
  NAND2_X1 U738 ( .A1(G93), .A2(n679), .ZN(n661) );
  NAND2_X1 U739 ( .A1(G80), .A2(n618), .ZN(n660) );
  NAND2_X1 U740 ( .A1(n661), .A2(n660), .ZN(n662) );
  OR2_X1 U741 ( .A1(n663), .A2(n662), .ZN(n702) );
  XOR2_X1 U742 ( .A(n664), .B(n702), .Z(G145) );
  NAND2_X1 U743 ( .A1(G85), .A2(n679), .ZN(n666) );
  NAND2_X1 U744 ( .A1(G72), .A2(n618), .ZN(n665) );
  NAND2_X1 U745 ( .A1(n666), .A2(n665), .ZN(n669) );
  NAND2_X1 U746 ( .A1(G60), .A2(n613), .ZN(n667) );
  XNOR2_X1 U747 ( .A(KEYINPUT69), .B(n667), .ZN(n668) );
  NOR2_X1 U748 ( .A1(n669), .A2(n668), .ZN(n671) );
  NAND2_X1 U749 ( .A1(n686), .A2(G47), .ZN(n670) );
  NAND2_X1 U750 ( .A1(n671), .A2(n670), .ZN(G290) );
  NAND2_X1 U751 ( .A1(G48), .A2(n686), .ZN(n673) );
  NAND2_X1 U752 ( .A1(G61), .A2(n613), .ZN(n672) );
  NAND2_X1 U753 ( .A1(n673), .A2(n672), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n618), .A2(G73), .ZN(n674) );
  XOR2_X1 U755 ( .A(KEYINPUT2), .B(n674), .Z(n675) );
  NOR2_X1 U756 ( .A1(n676), .A2(n675), .ZN(n678) );
  NAND2_X1 U757 ( .A1(n679), .A2(G86), .ZN(n677) );
  NAND2_X1 U758 ( .A1(n678), .A2(n677), .ZN(G305) );
  NAND2_X1 U759 ( .A1(G88), .A2(n679), .ZN(n681) );
  NAND2_X1 U760 ( .A1(G75), .A2(n618), .ZN(n680) );
  NAND2_X1 U761 ( .A1(n681), .A2(n680), .ZN(n685) );
  NAND2_X1 U762 ( .A1(G50), .A2(n686), .ZN(n683) );
  NAND2_X1 U763 ( .A1(G62), .A2(n613), .ZN(n682) );
  NAND2_X1 U764 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U765 ( .A1(n685), .A2(n684), .ZN(G166) );
  NAND2_X1 U766 ( .A1(G49), .A2(n686), .ZN(n688) );
  NAND2_X1 U767 ( .A1(G74), .A2(G651), .ZN(n687) );
  NAND2_X1 U768 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U769 ( .A(KEYINPUT81), .B(n689), .Z(n690) );
  NOR2_X1 U770 ( .A1(n613), .A2(n690), .ZN(n693) );
  NAND2_X1 U771 ( .A1(n691), .A2(G87), .ZN(n692) );
  NAND2_X1 U772 ( .A1(n693), .A2(n692), .ZN(G288) );
  XOR2_X1 U773 ( .A(n702), .B(G290), .Z(n694) );
  XNOR2_X1 U774 ( .A(n694), .B(G305), .ZN(n695) );
  XOR2_X1 U775 ( .A(n695), .B(KEYINPUT19), .Z(n697) );
  INV_X1 U776 ( .A(G299), .ZN(n771) );
  XNOR2_X1 U777 ( .A(n771), .B(G166), .ZN(n696) );
  XNOR2_X1 U778 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U779 ( .A(n698), .B(G288), .ZN(n865) );
  XOR2_X1 U780 ( .A(n865), .B(n699), .Z(n700) );
  NAND2_X1 U781 ( .A1(n700), .A2(G868), .ZN(n701) );
  XNOR2_X1 U782 ( .A(n701), .B(KEYINPUT82), .ZN(n705) );
  NAND2_X1 U783 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U784 ( .A1(n705), .A2(n704), .ZN(G295) );
  NAND2_X1 U785 ( .A1(G2084), .A2(G2078), .ZN(n706) );
  XNOR2_X1 U786 ( .A(n706), .B(KEYINPUT83), .ZN(n707) );
  XNOR2_X1 U787 ( .A(n707), .B(KEYINPUT20), .ZN(n708) );
  NAND2_X1 U788 ( .A1(n708), .A2(G2090), .ZN(n709) );
  XNOR2_X1 U789 ( .A(KEYINPUT21), .B(n709), .ZN(n710) );
  NAND2_X1 U790 ( .A1(n710), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U791 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U792 ( .A1(G220), .A2(G219), .ZN(n711) );
  XOR2_X1 U793 ( .A(KEYINPUT22), .B(n711), .Z(n712) );
  NOR2_X1 U794 ( .A1(G218), .A2(n712), .ZN(n713) );
  NAND2_X1 U795 ( .A1(G96), .A2(n713), .ZN(n864) );
  AND2_X1 U796 ( .A1(G2106), .A2(n864), .ZN(n718) );
  NAND2_X1 U797 ( .A1(G120), .A2(G108), .ZN(n714) );
  NOR2_X1 U798 ( .A1(G237), .A2(n714), .ZN(n715) );
  NAND2_X1 U799 ( .A1(G69), .A2(n715), .ZN(n863) );
  NAND2_X1 U800 ( .A1(G567), .A2(n863), .ZN(n716) );
  XOR2_X1 U801 ( .A(KEYINPUT84), .B(n716), .Z(n717) );
  NOR2_X1 U802 ( .A1(n718), .A2(n717), .ZN(G319) );
  INV_X1 U803 ( .A(G319), .ZN(n941) );
  NAND2_X1 U804 ( .A1(G483), .A2(G661), .ZN(n719) );
  NOR2_X1 U805 ( .A1(n941), .A2(n719), .ZN(n720) );
  XOR2_X1 U806 ( .A(KEYINPUT85), .B(n720), .Z(n862) );
  NAND2_X1 U807 ( .A1(n862), .A2(G36), .ZN(G176) );
  INV_X1 U808 ( .A(G166), .ZN(G303) );
  NOR2_X1 U809 ( .A1(G164), .A2(G1384), .ZN(n721) );
  NOR2_X1 U810 ( .A1(n721), .A2(n521), .ZN(n856) );
  NAND2_X1 U811 ( .A1(n925), .A2(G140), .ZN(n722) );
  XOR2_X1 U812 ( .A(KEYINPUT87), .B(n722), .Z(n724) );
  NAND2_X1 U813 ( .A1(n923), .A2(G104), .ZN(n723) );
  NAND2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U815 ( .A(KEYINPUT34), .B(n725), .ZN(n730) );
  NAND2_X1 U816 ( .A1(n920), .A2(G128), .ZN(n727) );
  NAND2_X1 U817 ( .A1(G116), .A2(n575), .ZN(n726) );
  NAND2_X1 U818 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U819 ( .A(KEYINPUT35), .B(n728), .Z(n729) );
  NOR2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U821 ( .A(KEYINPUT36), .B(n731), .ZN(n936) );
  XNOR2_X1 U822 ( .A(G2067), .B(KEYINPUT37), .ZN(n854) );
  NOR2_X1 U823 ( .A1(n936), .A2(n854), .ZN(n953) );
  NAND2_X1 U824 ( .A1(n856), .A2(n953), .ZN(n852) );
  NAND2_X1 U825 ( .A1(G131), .A2(n925), .ZN(n733) );
  NAND2_X1 U826 ( .A1(G95), .A2(n923), .ZN(n732) );
  NAND2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n737) );
  NAND2_X1 U828 ( .A1(n920), .A2(G119), .ZN(n735) );
  NAND2_X1 U829 ( .A1(G107), .A2(n905), .ZN(n734) );
  NAND2_X1 U830 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U831 ( .A1(n737), .A2(n736), .ZN(n914) );
  INV_X1 U832 ( .A(G1991), .ZN(n844) );
  NOR2_X1 U833 ( .A1(n914), .A2(n844), .ZN(n746) );
  NAND2_X1 U834 ( .A1(G141), .A2(n925), .ZN(n739) );
  NAND2_X1 U835 ( .A1(G117), .A2(n575), .ZN(n738) );
  NAND2_X1 U836 ( .A1(n739), .A2(n738), .ZN(n742) );
  NAND2_X1 U837 ( .A1(n923), .A2(G105), .ZN(n740) );
  XOR2_X1 U838 ( .A(KEYINPUT38), .B(n740), .Z(n741) );
  NOR2_X1 U839 ( .A1(n742), .A2(n741), .ZN(n744) );
  NAND2_X1 U840 ( .A1(n920), .A2(G129), .ZN(n743) );
  NAND2_X1 U841 ( .A1(n744), .A2(n743), .ZN(n915) );
  AND2_X1 U842 ( .A1(G1996), .A2(n915), .ZN(n745) );
  NOR2_X1 U843 ( .A1(n746), .A2(n745), .ZN(n955) );
  INV_X1 U844 ( .A(n856), .ZN(n747) );
  NOR2_X1 U845 ( .A1(n955), .A2(n747), .ZN(n848) );
  INV_X1 U846 ( .A(n848), .ZN(n748) );
  NAND2_X1 U847 ( .A1(n852), .A2(n748), .ZN(n842) );
  INV_X1 U848 ( .A(KEYINPUT97), .ZN(n790) );
  INV_X1 U849 ( .A(G40), .ZN(n749) );
  XNOR2_X1 U850 ( .A(G1996), .B(KEYINPUT91), .ZN(n1025) );
  NAND2_X1 U851 ( .A1(n797), .A2(G1341), .ZN(n751) );
  NAND2_X1 U852 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U853 ( .A1(n753), .A2(n978), .ZN(n755) );
  XNOR2_X1 U854 ( .A(n755), .B(n754), .ZN(n762) );
  XNOR2_X1 U855 ( .A(n757), .B(n756), .ZN(n761) );
  INV_X1 U856 ( .A(n797), .ZN(n775) );
  NOR2_X1 U857 ( .A1(n775), .A2(G1348), .ZN(n759) );
  NOR2_X1 U858 ( .A1(G2067), .A2(n797), .ZN(n758) );
  NOR2_X1 U859 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U860 ( .A1(n761), .A2(n760), .ZN(n764) );
  NAND2_X1 U861 ( .A1(n762), .A2(n973), .ZN(n763) );
  NAND2_X1 U862 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U863 ( .A1(G1956), .A2(n797), .ZN(n768) );
  NAND2_X1 U864 ( .A1(n775), .A2(G2072), .ZN(n766) );
  XOR2_X1 U865 ( .A(KEYINPUT27), .B(n766), .Z(n767) );
  NAND2_X1 U866 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U867 ( .A(KEYINPUT90), .B(n769), .Z(n770) );
  NOR2_X1 U868 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U869 ( .A(n772), .B(KEYINPUT28), .Z(n773) );
  XOR2_X1 U870 ( .A(KEYINPUT94), .B(KEYINPUT29), .Z(n774) );
  XNOR2_X1 U871 ( .A(G1961), .B(KEYINPUT89), .ZN(n998) );
  NAND2_X1 U872 ( .A1(n797), .A2(n998), .ZN(n777) );
  XNOR2_X1 U873 ( .A(KEYINPUT25), .B(G2078), .ZN(n1026) );
  NAND2_X1 U874 ( .A1(n775), .A2(n1026), .ZN(n776) );
  NAND2_X1 U875 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U876 ( .A1(n780), .A2(G171), .ZN(n778) );
  NAND2_X1 U877 ( .A1(n779), .A2(n778), .ZN(n806) );
  NOR2_X1 U878 ( .A1(G171), .A2(n780), .ZN(n786) );
  NAND2_X1 U879 ( .A1(G8), .A2(n797), .ZN(n835) );
  NOR2_X1 U880 ( .A1(G1966), .A2(n835), .ZN(n794) );
  NOR2_X1 U881 ( .A1(G2084), .A2(n797), .ZN(n791) );
  NOR2_X1 U882 ( .A1(n794), .A2(n791), .ZN(n781) );
  NAND2_X1 U883 ( .A1(G8), .A2(n781), .ZN(n782) );
  XNOR2_X1 U884 ( .A(KEYINPUT30), .B(n782), .ZN(n783) );
  XOR2_X1 U885 ( .A(KEYINPUT95), .B(n783), .Z(n784) );
  NOR2_X1 U886 ( .A1(G168), .A2(n784), .ZN(n785) );
  NOR2_X1 U887 ( .A1(n786), .A2(n785), .ZN(n788) );
  XOR2_X1 U888 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n787) );
  XNOR2_X1 U889 ( .A(n788), .B(n787), .ZN(n804) );
  NAND2_X1 U890 ( .A1(n806), .A2(n804), .ZN(n789) );
  XNOR2_X1 U891 ( .A(n790), .B(n789), .ZN(n796) );
  NAND2_X1 U892 ( .A1(n791), .A2(G8), .ZN(n792) );
  XOR2_X1 U893 ( .A(KEYINPUT88), .B(n792), .Z(n793) );
  NOR2_X1 U894 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U895 ( .A1(n796), .A2(n795), .ZN(n814) );
  INV_X1 U896 ( .A(G8), .ZN(n803) );
  NOR2_X1 U897 ( .A1(G1971), .A2(n835), .ZN(n799) );
  NOR2_X1 U898 ( .A1(G2090), .A2(n797), .ZN(n798) );
  NOR2_X1 U899 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U900 ( .A(n800), .B(KEYINPUT98), .ZN(n801) );
  NAND2_X1 U901 ( .A1(n801), .A2(G303), .ZN(n802) );
  OR2_X1 U902 ( .A1(n803), .A2(n802), .ZN(n807) );
  AND2_X1 U903 ( .A1(n804), .A2(n807), .ZN(n805) );
  NAND2_X1 U904 ( .A1(n806), .A2(n805), .ZN(n811) );
  INV_X1 U905 ( .A(n807), .ZN(n809) );
  AND2_X1 U906 ( .A1(G286), .A2(G8), .ZN(n808) );
  OR2_X1 U907 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U909 ( .A(n812), .B(KEYINPUT32), .ZN(n813) );
  NAND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n834) );
  NOR2_X1 U911 ( .A1(G1976), .A2(G288), .ZN(n820) );
  NOR2_X1 U912 ( .A1(G1971), .A2(G303), .ZN(n815) );
  NOR2_X1 U913 ( .A1(n820), .A2(n815), .ZN(n981) );
  INV_X1 U914 ( .A(KEYINPUT33), .ZN(n816) );
  AND2_X1 U915 ( .A1(n981), .A2(n816), .ZN(n817) );
  NAND2_X1 U916 ( .A1(n834), .A2(n817), .ZN(n826) );
  XOR2_X1 U917 ( .A(G1981), .B(G305), .Z(n987) );
  INV_X1 U918 ( .A(n835), .ZN(n818) );
  NAND2_X1 U919 ( .A1(G1976), .A2(G288), .ZN(n985) );
  AND2_X1 U920 ( .A1(n818), .A2(n985), .ZN(n819) );
  NOR2_X1 U921 ( .A1(KEYINPUT33), .A2(n819), .ZN(n823) );
  NAND2_X1 U922 ( .A1(n820), .A2(KEYINPUT33), .ZN(n821) );
  NOR2_X1 U923 ( .A1(n821), .A2(n835), .ZN(n822) );
  NOR2_X1 U924 ( .A1(n823), .A2(n822), .ZN(n824) );
  AND2_X1 U925 ( .A1(n987), .A2(n824), .ZN(n825) );
  NAND2_X1 U926 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U927 ( .A(n827), .B(KEYINPUT99), .ZN(n831) );
  NOR2_X1 U928 ( .A1(G1981), .A2(G305), .ZN(n828) );
  XOR2_X1 U929 ( .A(n828), .B(KEYINPUT24), .Z(n829) );
  NOR2_X1 U930 ( .A1(n835), .A2(n829), .ZN(n830) );
  NOR2_X1 U931 ( .A1(G2090), .A2(G303), .ZN(n832) );
  NAND2_X1 U932 ( .A1(G8), .A2(n832), .ZN(n833) );
  NAND2_X1 U933 ( .A1(n834), .A2(n833), .ZN(n836) );
  NAND2_X1 U934 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n837), .B(KEYINPUT100), .ZN(n838) );
  NAND2_X1 U936 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U937 ( .A(KEYINPUT101), .B(n840), .ZN(n841) );
  XNOR2_X1 U938 ( .A(G1986), .B(G290), .ZN(n975) );
  XOR2_X1 U939 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n843) );
  XNOR2_X1 U940 ( .A(KEYINPUT103), .B(n843), .ZN(n851) );
  NOR2_X1 U941 ( .A1(G1996), .A2(n915), .ZN(n957) );
  AND2_X1 U942 ( .A1(n844), .A2(n914), .ZN(n845) );
  XNOR2_X1 U943 ( .A(KEYINPUT102), .B(n845), .ZN(n965) );
  NOR2_X1 U944 ( .A1(G1986), .A2(G290), .ZN(n846) );
  NOR2_X1 U945 ( .A1(n965), .A2(n846), .ZN(n847) );
  NOR2_X1 U946 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U947 ( .A1(n957), .A2(n849), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n853) );
  NAND2_X1 U949 ( .A1(n853), .A2(n852), .ZN(n855) );
  NAND2_X1 U950 ( .A1(n936), .A2(n854), .ZN(n950) );
  NAND2_X1 U951 ( .A1(n855), .A2(n950), .ZN(n857) );
  NAND2_X1 U952 ( .A1(n857), .A2(n856), .ZN(n858) );
  NAND2_X1 U953 ( .A1(G2106), .A2(n859), .ZN(G217) );
  AND2_X1 U954 ( .A1(G15), .A2(G2), .ZN(n860) );
  NAND2_X1 U955 ( .A1(G661), .A2(n860), .ZN(G259) );
  NAND2_X1 U956 ( .A1(G3), .A2(G1), .ZN(n861) );
  NAND2_X1 U957 ( .A1(n862), .A2(n861), .ZN(G188) );
  XOR2_X1 U958 ( .A(G108), .B(KEYINPUT120), .Z(G238) );
  INV_X1 U960 ( .A(G120), .ZN(G236) );
  INV_X1 U961 ( .A(G96), .ZN(G221) );
  NOR2_X1 U962 ( .A1(n864), .A2(n863), .ZN(G325) );
  INV_X1 U963 ( .A(G325), .ZN(G261) );
  XOR2_X1 U964 ( .A(n865), .B(G286), .Z(n868) );
  XNOR2_X1 U965 ( .A(G171), .B(n866), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U967 ( .A(n978), .B(n869), .Z(n870) );
  NOR2_X1 U968 ( .A1(G37), .A2(n870), .ZN(G397) );
  XOR2_X1 U969 ( .A(G1976), .B(G1971), .Z(n872) );
  XNOR2_X1 U970 ( .A(G1986), .B(G1966), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n882) );
  XOR2_X1 U972 ( .A(G2474), .B(KEYINPUT41), .Z(n874) );
  XNOR2_X1 U973 ( .A(G1991), .B(KEYINPUT110), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U975 ( .A(G1956), .B(G1961), .Z(n876) );
  XNOR2_X1 U976 ( .A(G1996), .B(G1981), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U978 ( .A(n878), .B(n877), .Z(n880) );
  XNOR2_X1 U979 ( .A(KEYINPUT111), .B(KEYINPUT109), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n881) );
  XOR2_X1 U981 ( .A(n882), .B(n881), .Z(G229) );
  XOR2_X1 U982 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n884) );
  XNOR2_X1 U983 ( .A(KEYINPUT42), .B(G2678), .ZN(n883) );
  XNOR2_X1 U984 ( .A(n884), .B(n883), .ZN(n888) );
  XOR2_X1 U985 ( .A(KEYINPUT107), .B(G2090), .Z(n886) );
  XNOR2_X1 U986 ( .A(G2067), .B(G2072), .ZN(n885) );
  XNOR2_X1 U987 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U988 ( .A(n888), .B(n887), .Z(n890) );
  XNOR2_X1 U989 ( .A(G2096), .B(G2100), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n892) );
  XOR2_X1 U991 ( .A(G2084), .B(G2078), .Z(n891) );
  XNOR2_X1 U992 ( .A(n892), .B(n891), .ZN(G227) );
  NAND2_X1 U993 ( .A1(G124), .A2(n920), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n893), .B(KEYINPUT112), .ZN(n894) );
  XNOR2_X1 U995 ( .A(n894), .B(KEYINPUT44), .ZN(n896) );
  NAND2_X1 U996 ( .A1(G136), .A2(n925), .ZN(n895) );
  NAND2_X1 U997 ( .A1(n896), .A2(n895), .ZN(n900) );
  NAND2_X1 U998 ( .A1(G100), .A2(n923), .ZN(n898) );
  NAND2_X1 U999 ( .A1(G112), .A2(n905), .ZN(n897) );
  NAND2_X1 U1000 ( .A1(n898), .A2(n897), .ZN(n899) );
  NOR2_X1 U1001 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1002 ( .A(KEYINPUT113), .B(n901), .Z(G162) );
  NAND2_X1 U1003 ( .A1(G139), .A2(n925), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(G103), .A2(n923), .ZN(n902) );
  NAND2_X1 U1005 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1006 ( .A(KEYINPUT117), .B(n904), .Z(n910) );
  NAND2_X1 U1007 ( .A1(n920), .A2(G127), .ZN(n907) );
  NAND2_X1 U1008 ( .A1(G115), .A2(n905), .ZN(n906) );
  NAND2_X1 U1009 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U1010 ( .A(KEYINPUT47), .B(n908), .Z(n909) );
  NOR2_X1 U1011 ( .A1(n910), .A2(n909), .ZN(n946) );
  XNOR2_X1 U1012 ( .A(G164), .B(n946), .ZN(n919) );
  XOR2_X1 U1013 ( .A(KEYINPUT48), .B(KEYINPUT116), .Z(n912) );
  XNOR2_X1 U1014 ( .A(KEYINPUT46), .B(KEYINPUT118), .ZN(n911) );
  XNOR2_X1 U1015 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1016 ( .A(n954), .B(n913), .ZN(n917) );
  XOR2_X1 U1017 ( .A(n915), .B(n914), .Z(n916) );
  XNOR2_X1 U1018 ( .A(n917), .B(n916), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(n919), .B(n918), .ZN(n933) );
  NAND2_X1 U1020 ( .A1(n920), .A2(G130), .ZN(n922) );
  NAND2_X1 U1021 ( .A1(G118), .A2(n575), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n931) );
  NAND2_X1 U1023 ( .A1(n923), .A2(G106), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(n924), .B(KEYINPUT114), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(G142), .A2(n925), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(KEYINPUT45), .B(n928), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(KEYINPUT115), .B(n929), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1030 ( .A(n933), .B(n932), .Z(n935) );
  XNOR2_X1 U1031 ( .A(G160), .B(G162), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(n935), .B(n934), .ZN(n937) );
  XOR2_X1 U1033 ( .A(n937), .B(n936), .Z(n938) );
  NOR2_X1 U1034 ( .A1(G37), .A2(n938), .ZN(G395) );
  NOR2_X1 U1035 ( .A1(G229), .A2(G227), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(KEYINPUT49), .B(n939), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(G397), .A2(n940), .ZN(n945) );
  NOR2_X1 U1038 ( .A1(G401), .A2(n941), .ZN(n942) );
  XNOR2_X1 U1039 ( .A(KEYINPUT119), .B(n942), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(G395), .A2(n943), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(G225) );
  INV_X1 U1042 ( .A(G225), .ZN(G308) );
  INV_X1 U1043 ( .A(G69), .ZN(G235) );
  INV_X1 U1044 ( .A(KEYINPUT55), .ZN(n971) );
  XOR2_X1 U1045 ( .A(G2072), .B(n946), .Z(n948) );
  XOR2_X1 U1046 ( .A(G164), .B(G2078), .Z(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(n949), .B(KEYINPUT50), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n967) );
  XNOR2_X1 U1051 ( .A(G160), .B(G2084), .ZN(n963) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(G2090), .B(G162), .ZN(n956) );
  XNOR2_X1 U1054 ( .A(n956), .B(KEYINPUT121), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(KEYINPUT51), .B(n959), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT52), .B(n968), .ZN(n969) );
  XOR2_X1 U1062 ( .A(KEYINPUT122), .B(n969), .Z(n970) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n972), .A2(G29), .ZN(n997) );
  XNOR2_X1 U1065 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XNOR2_X1 U1066 ( .A(G1348), .B(n973), .ZN(n974) );
  NOR2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(G1971), .A2(G303), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(G1341), .B(n978), .ZN(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n993) );
  XNOR2_X1 U1072 ( .A(G171), .B(G1961), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(G1956), .B(G299), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n991) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G168), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n989), .Z(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n1051) );
  XOR2_X1 U1084 ( .A(G16), .B(KEYINPUT125), .Z(n1022) );
  XNOR2_X1 U1085 ( .A(G5), .B(n998), .ZN(n1019) );
  XOR2_X1 U1086 ( .A(G1966), .B(G21), .Z(n1010) );
  XOR2_X1 U1087 ( .A(G1348), .B(KEYINPUT59), .Z(n999) );
  XNOR2_X1 U1088 ( .A(G4), .B(n999), .ZN(n1007) );
  XOR2_X1 U1089 ( .A(G1956), .B(G20), .Z(n1002) );
  XOR2_X1 U1090 ( .A(G6), .B(KEYINPUT126), .Z(n1000) );
  XNOR2_X1 U1091 ( .A(n1000), .B(G1981), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G19), .B(G1341), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(n1005), .B(KEYINPUT127), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1017) );
  XNOR2_X1 U1099 ( .A(G1971), .B(G22), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(G23), .B(G1976), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(G1986), .B(G24), .Z(n1013) );
  NAND2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(KEYINPUT58), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(n1020), .B(KEYINPUT61), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1044) );
  XNOR2_X1 U1109 ( .A(G2084), .B(G34), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(n1023), .B(KEYINPUT54), .ZN(n1041) );
  XNOR2_X1 U1111 ( .A(G2090), .B(G35), .ZN(n1038) );
  XOR2_X1 U1112 ( .A(G2072), .B(G33), .Z(n1024) );
  NAND2_X1 U1113 ( .A1(n1024), .A2(G28), .ZN(n1035) );
  XNOR2_X1 U1114 ( .A(n1025), .B(G32), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(n1026), .B(G27), .ZN(n1027) );
  NAND2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1117 ( .A(KEYINPUT123), .B(n1029), .ZN(n1033) );
  XNOR2_X1 U1118 ( .A(G2067), .B(G26), .ZN(n1031) );
  XNOR2_X1 U1119 ( .A(G1991), .B(G25), .ZN(n1030) );
  NOR2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1121 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XNOR2_X1 U1123 ( .A(KEYINPUT53), .B(n1036), .ZN(n1037) );
  NOR2_X1 U1124 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  XOR2_X1 U1125 ( .A(KEYINPUT124), .B(n1039), .Z(n1040) );
  NOR2_X1 U1126 ( .A1(n1041), .A2(n1040), .ZN(n1045) );
  NAND2_X1 U1127 ( .A1(KEYINPUT55), .A2(n1045), .ZN(n1042) );
  NAND2_X1 U1128 ( .A1(G11), .A2(n1042), .ZN(n1043) );
  NOR2_X1 U1129 ( .A1(n1044), .A2(n1043), .ZN(n1049) );
  INV_X1 U1130 ( .A(n1045), .ZN(n1047) );
  NOR2_X1 U1131 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1046) );
  NAND2_X1 U1132 ( .A1(n1047), .A2(n1046), .ZN(n1048) );
  NAND2_X1 U1133 ( .A1(n1049), .A2(n1048), .ZN(n1050) );
  NOR2_X1 U1134 ( .A1(n1051), .A2(n1050), .ZN(n1052) );
  XNOR2_X1 U1135 ( .A(n1052), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1136 ( .A(G311), .ZN(G150) );
endmodule

