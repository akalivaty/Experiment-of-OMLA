//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(G77), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(G244), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G68), .A2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n216), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n208), .B1(new_n211), .B2(new_n212), .C1(new_n223), .C2(KEYINPUT1), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n229), .B(new_n232), .Z(G358));
  XOR2_X1   g0033(.A(G87), .B(G97), .Z(new_n234));
  XOR2_X1   g0034(.A(G107), .B(G116), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G50), .B(G68), .Z(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G351));
  INV_X1    g0040(.A(KEYINPUT74), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT3), .B(G33), .ZN(new_n242));
  NOR2_X1   g0042(.A1(G222), .A2(G1698), .ZN(new_n243));
  INV_X1    g0043(.A(G1698), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n244), .A2(G223), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n242), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g0046(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n247));
  OAI211_X1 g0047(.A(new_n246), .B(new_n247), .C1(new_n217), .C2(new_n242), .ZN(new_n248));
  INV_X1    g0048(.A(G274), .ZN(new_n249));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n249), .B1(new_n210), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G226), .ZN(new_n256));
  INV_X1    g0056(.A(G1), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT66), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G1), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n258), .B(new_n260), .C1(G41), .C2(G45), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n210), .A2(new_n250), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n248), .B(new_n255), .C1(new_n256), .C2(new_n263), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n264), .A2(G179), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n209), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  INV_X1    g0068(.A(G20), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G150), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n268), .A2(new_n270), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G50), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n269), .B1(new_n201), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n267), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n258), .A2(new_n260), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G20), .ZN(new_n279));
  INV_X1    g0079(.A(new_n267), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n258), .A2(new_n260), .A3(G13), .A4(G20), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n279), .A2(G50), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n277), .B(new_n282), .C1(G50), .C2(new_n281), .ZN(new_n283));
  INV_X1    g0083(.A(G169), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n264), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n265), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G190), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n264), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(G200), .B2(new_n264), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n283), .B(KEYINPUT9), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT10), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n290), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n287), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n256), .A2(new_n244), .ZN(new_n297));
  INV_X1    g0097(.A(G232), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G1698), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n242), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G97), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT68), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n300), .A2(KEYINPUT68), .A3(new_n301), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n247), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT13), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n261), .A2(new_n262), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n308), .A2(G238), .B1(new_n251), .B2(new_n254), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n307), .B1(new_n306), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g0111(.A(G169), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT14), .ZN(new_n313));
  INV_X1    g0113(.A(new_n311), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(G179), .A3(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT14), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(G169), .C1(new_n310), .C2(new_n311), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n313), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G68), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G20), .ZN(new_n321));
  INV_X1    g0121(.A(G77), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n321), .B1(new_n270), .B2(new_n322), .C1(new_n273), .C2(new_n275), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n323), .A2(KEYINPUT69), .A3(new_n267), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT69), .B1(new_n323), .B2(new_n267), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT11), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT11), .B1(new_n324), .B2(new_n325), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT12), .B1(new_n281), .B2(G68), .ZN(new_n330));
  OR3_X1    g0130(.A1(new_n281), .A2(KEYINPUT12), .A3(G68), .ZN(new_n331));
  INV_X1    g0131(.A(new_n281), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(new_n267), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n320), .B1(new_n278), .B2(G20), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n330), .A2(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n328), .A2(new_n329), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n319), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n314), .A2(G190), .A3(new_n315), .ZN(new_n338));
  INV_X1    g0138(.A(new_n336), .ZN(new_n339));
  OAI21_X1  g0139(.A(G200), .B1(new_n310), .B2(new_n311), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n242), .A2(G238), .A3(G1698), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n242), .A2(G232), .A3(new_n244), .ZN(new_n343));
  INV_X1    g0143(.A(G107), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(new_n343), .C1(new_n344), .C2(new_n242), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n247), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n308), .A2(G244), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n346), .A2(new_n255), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(G179), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n284), .B2(new_n348), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n217), .A2(G20), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT15), .B(G87), .ZN(new_n352));
  OAI221_X1 g0152(.A(new_n351), .B1(new_n273), .B2(new_n268), .C1(new_n270), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n267), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n333), .A2(G77), .A3(new_n279), .ZN(new_n355));
  INV_X1    g0155(.A(new_n217), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n332), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(new_n355), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT67), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n359), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n350), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n348), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G190), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n348), .A2(G200), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n360), .A2(new_n365), .A3(new_n361), .A4(new_n366), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n296), .A2(new_n337), .A3(new_n341), .A4(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n268), .A2(new_n267), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n279), .A2(new_n370), .B1(new_n332), .B2(new_n268), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G58), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(new_n320), .ZN(new_n374));
  OAI21_X1  g0174(.A(G20), .B1(new_n374), .B2(new_n201), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n272), .A2(G159), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(G33), .ZN(new_n380));
  INV_X1    g0180(.A(G33), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT3), .ZN(new_n382));
  AOI21_X1  g0182(.A(G20), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(KEYINPUT7), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n381), .B2(KEYINPUT3), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n379), .A2(KEYINPUT71), .A3(G33), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n382), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(G20), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT72), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(KEYINPUT72), .A3(new_n390), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n384), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n378), .B1(new_n395), .B2(new_n320), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT16), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT70), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n383), .B2(KEYINPUT7), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n380), .A2(new_n382), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n390), .ZN(new_n402));
  OAI211_X1 g0202(.A(KEYINPUT70), .B(new_n389), .C1(new_n242), .C2(G20), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n377), .B1(new_n404), .B2(G68), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n280), .B1(new_n405), .B2(KEYINPUT16), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n372), .B1(new_n398), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT73), .ZN(new_n408));
  NOR2_X1   g0208(.A1(G223), .A2(G1698), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n256), .B2(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n242), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G33), .A2(G87), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n408), .B1(new_n413), .B2(new_n262), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n262), .B1(new_n411), .B2(new_n412), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT73), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n255), .B1(new_n263), .B2(new_n298), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(G179), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n418), .A2(new_n415), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n284), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT18), .B1(new_n407), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n418), .A2(G190), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n414), .A2(new_n425), .A3(new_n416), .ZN(new_n426));
  INV_X1    g0226(.A(G200), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n418), .B2(new_n415), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n384), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n388), .A2(KEYINPUT72), .A3(new_n390), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT72), .B1(new_n388), .B2(new_n390), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G68), .ZN(new_n434));
  AOI21_X1  g0234(.A(KEYINPUT16), .B1(new_n434), .B2(new_n378), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n403), .A2(new_n402), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n381), .A2(KEYINPUT3), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n379), .A2(G33), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n269), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT70), .B1(new_n439), .B2(new_n389), .ZN(new_n440));
  OAI21_X1  g0240(.A(G68), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(KEYINPUT16), .A3(new_n378), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n267), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n371), .B(new_n429), .C1(new_n435), .C2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT17), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n371), .B1(new_n435), .B2(new_n443), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT18), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n417), .A2(new_n419), .B1(new_n284), .B2(new_n421), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n398), .A2(new_n406), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n451), .A2(KEYINPUT17), .A3(new_n371), .A4(new_n429), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n424), .A2(new_n446), .A3(new_n450), .A4(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n241), .B1(new_n369), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n296), .A2(new_n368), .ZN(new_n455));
  INV_X1    g0255(.A(new_n341), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n319), .B2(new_n336), .ZN(new_n457));
  AND4_X1   g0257(.A1(new_n424), .A2(new_n446), .A3(new_n450), .A4(new_n452), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n455), .A2(new_n457), .A3(KEYINPUT74), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n258), .A2(new_n260), .A3(G33), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n281), .A2(new_n280), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G116), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n281), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  INV_X1    g0267(.A(G97), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n467), .B(new_n269), .C1(G33), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n464), .A2(G20), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(new_n267), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT20), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n469), .A2(new_n267), .A3(KEYINPUT20), .A4(new_n470), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(KEYINPUT78), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT78), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n471), .A2(new_n476), .A3(new_n472), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n466), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n258), .A2(new_n260), .A3(G45), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n251), .A3(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(G270), .B(new_n262), .C1(new_n479), .C2(new_n483), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n242), .A2(G264), .A3(G1698), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n242), .A2(G257), .A3(new_n244), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n401), .A2(G303), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n247), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n478), .A2(new_n493), .A3(KEYINPUT21), .A4(G169), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT79), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n284), .B1(new_n487), .B2(new_n492), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n497), .A2(new_n478), .A3(KEYINPUT79), .A4(KEYINPUT21), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n478), .ZN(new_n500));
  XOR2_X1   g0300(.A(KEYINPUT80), .B(KEYINPUT21), .Z(new_n501));
  INV_X1    g0301(.A(G179), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n500), .A2(new_n501), .B1(new_n503), .B2(new_n478), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n493), .A2(G200), .ZN(new_n505));
  INV_X1    g0305(.A(new_n478), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n505), .B(new_n506), .C1(new_n288), .C2(new_n493), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n499), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  XOR2_X1   g0308(.A(KEYINPUT84), .B(G294), .Z(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G33), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n242), .A2(G257), .A3(G1698), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n242), .A2(G250), .A3(new_n244), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n247), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n247), .B1(new_n480), .B2(new_n484), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G264), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n516), .A3(new_n485), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n284), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n514), .A2(new_n516), .A3(new_n502), .A4(new_n485), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n380), .A2(new_n382), .A3(new_n269), .A4(G87), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT81), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT81), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n242), .A2(new_n523), .A3(new_n269), .A4(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n522), .A2(new_n524), .A3(KEYINPUT22), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT23), .B1(new_n269), .B2(G107), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT23), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(new_n344), .A3(G20), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n269), .A2(G33), .A3(G116), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT82), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n529), .A2(new_n531), .A3(new_n532), .A4(KEYINPUT82), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n527), .A2(new_n528), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT24), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n525), .A2(new_n526), .B1(new_n535), .B2(new_n536), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(new_n541), .A3(new_n528), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n280), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n462), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G107), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT83), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n546), .B(KEYINPUT25), .C1(new_n281), .C2(G107), .ZN(new_n547));
  XNOR2_X1  g0347(.A(KEYINPUT83), .B(KEYINPUT25), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n332), .A2(new_n344), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n545), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n520), .B1(new_n543), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n538), .A2(KEYINPUT24), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n541), .B1(new_n540), .B2(new_n528), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n267), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n550), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n517), .A2(new_n427), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G190), .B2(new_n517), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT76), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n380), .A2(new_n382), .A3(G244), .A4(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n380), .A2(new_n382), .A3(G238), .A4(new_n244), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G116), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(G250), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n247), .B1(new_n479), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n278), .A2(G45), .A3(new_n249), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n247), .A2(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n560), .B1(new_n568), .B2(new_n502), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n564), .A2(new_n247), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n566), .A2(new_n567), .ZN(new_n571));
  AND4_X1   g0371(.A1(new_n560), .A2(new_n570), .A3(new_n571), .A4(new_n502), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n380), .A2(new_n382), .A3(new_n269), .A4(G68), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n270), .B2(new_n468), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n269), .B1(new_n301), .B2(new_n575), .ZN(new_n577));
  NOR2_X1   g0377(.A1(G97), .A2(G107), .ZN(new_n578));
  INV_X1    g0378(.A(G87), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n577), .A2(KEYINPUT77), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT77), .B1(new_n577), .B2(new_n580), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n574), .B(new_n576), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(new_n267), .B1(new_n332), .B2(new_n352), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n462), .A2(new_n352), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n570), .A2(new_n571), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n584), .A2(new_n586), .B1(new_n284), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n574), .A2(new_n576), .ZN(new_n589));
  INV_X1    g0389(.A(new_n582), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n577), .A2(new_n580), .A3(KEYINPUT77), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n352), .ZN(new_n593));
  OAI22_X1  g0393(.A1(new_n592), .A2(new_n280), .B1(new_n281), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n462), .A2(new_n579), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n570), .A2(new_n571), .A3(G190), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n427), .B1(new_n570), .B2(new_n571), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n573), .A2(new_n588), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n380), .A2(new_n382), .A3(G250), .A4(G1698), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT75), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n242), .A2(KEYINPUT75), .A3(G250), .A4(G1698), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n380), .A2(new_n382), .A3(G244), .A4(new_n244), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT4), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n242), .A2(KEYINPUT4), .A3(G244), .A4(new_n244), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n610), .A3(new_n467), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n247), .B1(new_n606), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(G257), .B(new_n262), .C1(new_n479), .C2(new_n483), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n485), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n612), .A2(new_n288), .A3(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n609), .A2(new_n610), .A3(new_n467), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n605), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n614), .B1(new_n618), .B2(new_n247), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n616), .B1(new_n619), .B2(G200), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n332), .A2(new_n468), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n468), .B2(new_n462), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n344), .A2(KEYINPUT6), .A3(G97), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n468), .A2(new_n344), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n624), .A2(new_n578), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n623), .B1(new_n625), .B2(KEYINPUT6), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n626), .A2(G20), .B1(G77), .B2(new_n272), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n395), .B2(new_n344), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n622), .B1(new_n628), .B2(new_n267), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n620), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n612), .A2(new_n502), .A3(new_n615), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n262), .B1(new_n617), .B2(new_n605), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n284), .B1(new_n632), .B2(new_n614), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n433), .A2(G107), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n280), .B1(new_n634), .B2(new_n627), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n631), .B(new_n633), .C1(new_n635), .C2(new_n622), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n600), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n460), .A2(new_n508), .A3(new_n559), .A4(new_n637), .ZN(G372));
  NAND3_X1  g0438(.A1(new_n551), .A2(new_n499), .A3(new_n504), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT85), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n587), .A2(new_n284), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n568), .A2(new_n502), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n641), .B(new_n642), .C1(new_n594), .C2(new_n585), .ZN(new_n643));
  INV_X1    g0443(.A(new_n598), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n568), .A2(G190), .ZN(new_n645));
  INV_X1    g0445(.A(new_n595), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n644), .A2(new_n584), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  AND4_X1   g0448(.A1(new_n558), .A2(new_n636), .A3(new_n630), .A4(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT85), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n551), .A2(new_n650), .A3(new_n499), .A4(new_n504), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n640), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n633), .A2(new_n631), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(new_n629), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n653), .B1(new_n655), .B2(new_n600), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n643), .A2(new_n647), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n636), .A2(new_n657), .A3(KEYINPUT26), .ZN(new_n658));
  INV_X1    g0458(.A(new_n643), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n460), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n424), .A2(new_n450), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n337), .A2(new_n363), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n446), .A2(new_n452), .A3(new_n341), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n295), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n294), .B1(new_n290), .B2(new_n291), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n286), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n662), .A2(new_n670), .ZN(G369));
  INV_X1    g0471(.A(G13), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(G20), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n278), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT86), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT27), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n677), .A2(new_n678), .A3(G213), .A4(G343), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n478), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n508), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n499), .A2(new_n504), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n681), .ZN(new_n685));
  OAI21_X1  g0485(.A(G330), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT87), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n682), .B1(new_n684), .B2(new_n681), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(KEYINPUT87), .A3(G330), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n543), .A2(new_n550), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n559), .B1(new_n693), .B2(new_n679), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n551), .A2(new_n679), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n551), .A2(new_n680), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n499), .A2(new_n504), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n679), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT88), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n701), .A2(KEYINPUT88), .A3(new_n679), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n700), .B1(new_n696), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n699), .A2(new_n707), .ZN(G399));
  INV_X1    g0508(.A(new_n206), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G41), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n580), .A2(G116), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(G1), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n212), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g0514(.A(new_n714), .B(KEYINPUT28), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n630), .A2(new_n636), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT89), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n657), .B1(new_n693), .B2(new_n557), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT89), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n630), .A2(new_n636), .A3(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n717), .A2(new_n639), .A3(new_n718), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n655), .A2(new_n600), .A3(new_n653), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT26), .B1(new_n636), .B2(new_n657), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n722), .A2(new_n723), .A3(new_n643), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n721), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT29), .B1(new_n725), .B2(new_n680), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n661), .A2(new_n679), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(KEYINPUT29), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G330), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n568), .A2(new_n516), .A3(new_n514), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n503), .A2(new_n730), .A3(new_n619), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT30), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n503), .A2(new_n619), .A3(new_n730), .A4(KEYINPUT30), .ZN(new_n734));
  INV_X1    g0534(.A(new_n619), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n568), .A2(G179), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n493), .A3(new_n517), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n733), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n680), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT31), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n508), .A2(new_n559), .A3(new_n637), .A4(new_n679), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n729), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n728), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n715), .B1(new_n743), .B2(G1), .ZN(G364));
  AOI21_X1  g0544(.A(new_n257), .B1(new_n673), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n710), .A2(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n692), .B(new_n748), .C1(G330), .C2(new_n689), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n209), .B1(G20), .B2(new_n284), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n269), .A2(G190), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT94), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n754), .A2(G179), .A3(new_n427), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n755), .A2(KEYINPUT95), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(KEYINPUT95), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n754), .A2(G179), .A3(G200), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT97), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(KEYINPUT97), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(G283), .A2(new_n759), .B1(new_n764), .B2(G329), .ZN(new_n765));
  NAND3_X1  g0565(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT93), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n288), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G326), .ZN(new_n769));
  INV_X1    g0569(.A(new_n509), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G179), .A2(G200), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n269), .B1(new_n771), .B2(G190), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n502), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n752), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n242), .B1(new_n776), .B2(G311), .ZN(new_n777));
  INV_X1    g0577(.A(G303), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n269), .A2(new_n288), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(new_n502), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n779), .A2(new_n774), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n777), .B1(new_n778), .B2(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n767), .A2(G190), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT33), .B(G317), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n773), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n765), .A2(new_n769), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n759), .A2(G107), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n242), .B1(new_n782), .B2(new_n373), .C1(new_n579), .C2(new_n780), .ZN(new_n789));
  INV_X1    g0589(.A(new_n768), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n275), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n776), .A2(KEYINPUT92), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n776), .A2(KEYINPUT92), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n789), .B(new_n791), .C1(new_n217), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n760), .A2(G159), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT32), .Z(new_n798));
  XOR2_X1   g0598(.A(new_n772), .B(KEYINPUT96), .Z(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n468), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G68), .B2(new_n784), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n788), .A2(new_n796), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n751), .B1(new_n787), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G13), .A2(G33), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G20), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n750), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n239), .A2(new_n253), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n401), .A2(new_n206), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT90), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(G45), .B2(new_n212), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n810), .B1(new_n814), .B2(KEYINPUT91), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(KEYINPUT91), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n709), .A2(new_n401), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G355), .B1(new_n464), .B2(new_n709), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n809), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n804), .A2(new_n748), .A3(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n807), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n820), .B1(new_n689), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n749), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  INV_X1    g0624(.A(new_n367), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n679), .B1(new_n360), .B2(new_n361), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n363), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n350), .A2(new_n362), .A3(new_n679), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n727), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n829), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n661), .A2(new_n679), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n742), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n711), .B2(new_n745), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n830), .A2(new_n742), .A3(new_n832), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(G294), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n401), .B1(new_n782), .B2(new_n837), .C1(new_n344), .C2(new_n780), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n838), .B(new_n801), .C1(G116), .C2(new_n795), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n759), .A2(G87), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n764), .A2(G311), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G283), .A2(new_n784), .B1(new_n768), .B2(G303), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(new_n782), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n795), .A2(G159), .B1(G143), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  INV_X1    g0646(.A(new_n784), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n845), .B1(new_n846), .B2(new_n790), .C1(new_n271), .C2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT98), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n242), .B1(new_n772), .B2(new_n373), .C1(new_n780), .C2(new_n275), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n758), .A2(new_n320), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n851), .B(new_n852), .C1(G132), .C2(new_n764), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n843), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n750), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n750), .A2(new_n805), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n748), .B1(new_n322), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n857), .B(new_n859), .C1(new_n806), .C2(new_n831), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n836), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(G384));
  INV_X1    g0662(.A(KEYINPUT100), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n441), .A2(new_n378), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n397), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n372), .B1(new_n406), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n677), .A2(new_n678), .A3(G213), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n405), .A2(KEYINPUT16), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n371), .B1(new_n443), .B2(new_n869), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n677), .A2(new_n678), .A3(G213), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(KEYINPUT100), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n453), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT101), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT101), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n453), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n444), .B1(new_n423), .B2(new_n866), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT37), .B1(new_n873), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n447), .A2(new_n449), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n447), .A2(new_n871), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT37), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .A4(new_n444), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n878), .B2(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n453), .A2(new_n876), .A3(new_n873), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n876), .B1(new_n453), .B2(new_n873), .ZN(new_n888));
  OAI211_X1 g0688(.A(KEYINPUT38), .B(new_n885), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT103), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(KEYINPUT31), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n739), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n893), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n738), .A2(new_n680), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n741), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n680), .A2(new_n336), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n337), .A2(new_n341), .A3(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n336), .B(new_n680), .C1(new_n319), .C2(new_n456), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n897), .A2(new_n901), .A3(new_n902), .A4(new_n831), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n897), .A2(new_n901), .A3(new_n831), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n881), .A2(new_n882), .A3(new_n444), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(new_n883), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n458), .A2(new_n882), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n904), .B1(new_n889), .B2(new_n909), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n891), .A2(new_n903), .B1(new_n910), .B2(new_n902), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n460), .A2(new_n897), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n729), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n912), .B2(new_n911), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT104), .ZN(new_n915));
  INV_X1    g0715(.A(new_n901), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n832), .B2(new_n828), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n886), .B2(new_n890), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n663), .A2(new_n867), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT102), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n919), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n905), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n889), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n923), .B1(new_n926), .B2(new_n917), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT102), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n889), .A2(new_n909), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT39), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n925), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n319), .A2(new_n336), .A3(new_n679), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n922), .A2(new_n928), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n670), .B1(new_n728), .B2(new_n460), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n915), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n915), .A2(new_n938), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n939), .B(new_n940), .C1(new_n278), .C2(new_n673), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n464), .B(new_n211), .C1(new_n626), .C2(KEYINPUT35), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(KEYINPUT35), .B2(new_n626), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT36), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n212), .A2(new_n374), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n945), .A2(new_n356), .B1(G50), .B2(new_n320), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n278), .A2(G13), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT99), .Z(new_n950));
  NAND2_X1  g0750(.A1(new_n941), .A2(new_n950), .ZN(G367));
  OAI211_X1 g0751(.A(new_n717), .B(new_n720), .C1(new_n629), .C2(new_n679), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n952), .A2(new_n551), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n680), .B1(new_n953), .B2(new_n636), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n655), .A2(new_n680), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n956), .A2(new_n696), .A3(new_n706), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n954), .B1(KEYINPUT42), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n957), .A2(KEYINPUT42), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n648), .B1(new_n596), .B2(new_n679), .ZN(new_n961));
  OR3_X1    g0761(.A1(new_n679), .A2(new_n596), .A3(new_n643), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n960), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n958), .A2(new_n965), .A3(new_n964), .A4(new_n959), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n698), .A2(new_n956), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n970), .A2(new_n971), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n710), .B(KEYINPUT41), .Z(new_n975));
  INV_X1    g0775(.A(KEYINPUT106), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n689), .A2(KEYINPUT87), .A3(G330), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT87), .B1(new_n689), .B2(G330), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n688), .A2(KEYINPUT106), .A3(new_n690), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n696), .A2(new_n706), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n694), .A2(new_n704), .A3(new_n695), .A4(new_n705), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n979), .A2(new_n980), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n691), .A2(new_n983), .A3(new_n976), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n743), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT107), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT107), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n990), .A3(new_n743), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n691), .A2(KEYINPUT105), .A3(new_n696), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n707), .A2(new_n956), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT45), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT44), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n707), .A2(new_n996), .A3(new_n956), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n707), .B2(new_n956), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n992), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  AND3_X1   g0800(.A1(new_n995), .A2(new_n992), .A3(new_n999), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n989), .B(new_n991), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n975), .B1(new_n1002), .B2(new_n743), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n974), .B1(new_n1003), .B2(new_n746), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n812), .A2(new_n232), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n809), .B1(new_n709), .B2(new_n593), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n748), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(G159), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n800), .A2(new_n320), .B1(new_n1008), .B2(new_n847), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n242), .B1(new_n782), .B2(new_n271), .C1(new_n373), .C2(new_n780), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n760), .B2(G137), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n795), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1011), .B1(new_n275), .B2(new_n1012), .C1(new_n758), .C2(new_n356), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1009), .B(new_n1013), .C1(G143), .C2(new_n768), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT110), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n759), .A2(G97), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n784), .A2(new_n509), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n401), .B1(new_n772), .B2(new_n344), .ZN(new_n1018));
  OR3_X1    g0818(.A1(new_n780), .A2(KEYINPUT46), .A3(new_n464), .ZN(new_n1019));
  OAI21_X1  g0819(.A(KEYINPUT46), .B1(new_n780), .B2(new_n464), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n795), .A2(G283), .B1(G317), .B2(new_n760), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1016), .A2(new_n1017), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n768), .A2(G311), .B1(G303), .B2(new_n844), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT108), .Z(new_n1025));
  NOR2_X1   g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1015), .B1(KEYINPUT109), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(KEYINPUT109), .B2(new_n1026), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT47), .Z(new_n1029));
  OAI221_X1 g0829(.A(new_n1007), .B1(new_n821), .B2(new_n963), .C1(new_n1029), .C2(new_n751), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1004), .A2(new_n1030), .ZN(G387));
  NAND2_X1  g0831(.A1(new_n989), .A2(new_n991), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n710), .B(KEYINPUT113), .Z(new_n1033));
  OAI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n743), .C2(new_n987), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n799), .A2(new_n593), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G50), .A2(new_n844), .B1(new_n776), .B2(G68), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n780), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n217), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n242), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G150), .B2(new_n760), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n268), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G159), .A2(new_n768), .B1(new_n784), .B2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1016), .A2(new_n1035), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n242), .B1(new_n760), .B2(G326), .ZN(new_n1044));
  INV_X1    g0844(.A(G283), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n770), .A2(new_n780), .B1(new_n1045), .B2(new_n772), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n795), .A2(G303), .B1(G317), .B2(new_n844), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n784), .A2(G311), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(new_n781), .C2(new_n790), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n1050), .B2(new_n1049), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1044), .B1(new_n464), .B2(new_n758), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1043), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n751), .B1(new_n1056), .B2(KEYINPUT112), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(KEYINPUT112), .B2(new_n1056), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n696), .A2(new_n821), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n712), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1060), .A2(new_n817), .B1(new_n344), .B2(new_n709), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT111), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n229), .A2(new_n253), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1041), .A2(new_n275), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT50), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n712), .B(new_n253), .C1(new_n320), .C2(new_n322), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n812), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1062), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n748), .B(new_n1059), .C1(new_n808), .C2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n987), .A2(new_n746), .B1(new_n1058), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1034), .A2(new_n1070), .ZN(G393));
  INV_X1    g0871(.A(new_n1032), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n995), .A2(new_n999), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(new_n699), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1002), .B(new_n1033), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n847), .A2(new_n778), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n242), .B1(new_n1037), .B2(G283), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n464), .B2(new_n772), .C1(new_n837), .C2(new_n775), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1076), .B(new_n1078), .C1(G322), .C2(new_n760), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n768), .A2(G317), .B1(G311), .B2(new_n844), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1081));
  XNOR2_X1  g0881(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n788), .A3(new_n1082), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n242), .B1(new_n320), .B2(new_n780), .C1(new_n1012), .C2(new_n268), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G143), .B2(new_n760), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n800), .A2(new_n322), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G50), .B2(new_n784), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1085), .A2(new_n840), .A3(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n768), .A2(G150), .B1(G159), .B2(new_n844), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT51), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1083), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n750), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n812), .A2(new_n236), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n809), .B1(G97), .B2(new_n709), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n748), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1092), .B(new_n1095), .C1(new_n956), .C2(new_n821), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1074), .B2(new_n746), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1075), .A2(new_n1098), .ZN(G390));
  AOI211_X1 g0899(.A(new_n680), .B(new_n829), .C1(new_n652), .C2(new_n660), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n828), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n901), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n933), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n925), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT39), .B1(new_n889), .B2(new_n909), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1103), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n362), .A2(new_n680), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1107), .A2(new_n367), .B1(new_n350), .B2(new_n362), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n680), .B(new_n1108), .C1(new_n721), .C2(new_n724), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n901), .B1(new_n1109), .B2(new_n1101), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n929), .A2(new_n1110), .A3(new_n933), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n740), .A2(new_n741), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n829), .A2(new_n729), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1112), .A2(new_n901), .A3(new_n1113), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1106), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n931), .A2(new_n932), .B1(new_n1102), .B2(new_n933), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT115), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n897), .A2(new_n1113), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1122), .A2(new_n916), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1117), .A2(new_n1120), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n746), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n805), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n858), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n747), .B1(new_n1041), .B2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1012), .A2(new_n468), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n401), .B1(new_n782), .B2(new_n464), .C1(new_n579), .C2(new_n780), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1129), .A2(new_n1086), .A3(new_n1130), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n344), .B2(new_n847), .C1(new_n1045), .C2(new_n790), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n320), .A2(new_n758), .B1(new_n763), .B2(new_n837), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n764), .A2(G125), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n780), .A2(new_n271), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  INV_X1    g0936(.A(G132), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1136), .B(new_n242), .C1(new_n1137), .C2(new_n782), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT54), .B(G143), .Z(new_n1139));
  AOI21_X1  g0939(.A(new_n1138), .B1(new_n795), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1134), .B(new_n1140), .C1(new_n275), .C2(new_n758), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n768), .A2(G128), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n847), .B2(new_n846), .C1(new_n800), .C2(new_n1008), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1132), .A2(new_n1133), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1128), .B1(new_n1144), .B2(new_n750), .ZN(new_n1145));
  XOR2_X1   g0945(.A(new_n1145), .B(KEYINPUT117), .Z(new_n1146));
  NAND2_X1  g0946(.A1(new_n1126), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1111), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1123), .B1(new_n1118), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n901), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1123), .A2(new_n1150), .B1(new_n1101), .B2(new_n1100), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1109), .A2(new_n1101), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1122), .A2(new_n916), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1152), .A2(new_n1114), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n460), .A2(G330), .A3(new_n897), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT116), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n460), .A2(KEYINPUT116), .A3(G330), .A4(new_n897), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1155), .A2(new_n1160), .A3(new_n937), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1116), .B1(new_n1106), .B2(new_n1115), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n1118), .A2(new_n1119), .A3(KEYINPUT115), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1149), .B(new_n1161), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1033), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1124), .A2(new_n1161), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1125), .B(new_n1147), .C1(new_n1165), .C2(new_n1166), .ZN(G378));
  OAI21_X1  g0967(.A(new_n935), .B1(new_n927), .B2(KEYINPUT102), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n921), .B(new_n923), .C1(new_n926), .C2(new_n917), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT122), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n904), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n902), .B1(new_n929), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n903), .B1(new_n925), .B2(new_n889), .ZN(new_n1173));
  OAI21_X1  g0973(.A(G330), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n286), .B1(new_n667), .B2(new_n668), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n871), .A2(new_n283), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(KEYINPUT55), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT55), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n871), .A2(new_n1178), .A3(new_n283), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1175), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1181));
  NAND2_X1  g0981(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n296), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1181), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1174), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT121), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1185), .A2(new_n1186), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1181), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT121), .B1(new_n1193), .B2(new_n1184), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1190), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g0995(.A(G330), .B(new_n1195), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1170), .A2(new_n1188), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1188), .A2(new_n1196), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1198), .A2(new_n936), .A3(KEYINPUT122), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1160), .A2(new_n937), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1164), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT57), .B1(new_n1200), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1201), .B1(new_n1124), .B2(new_n1161), .ZN(new_n1205));
  AOI21_X1  g1005(.A(KEYINPUT102), .B1(new_n918), .B2(new_n919), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1187), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n911), .B2(G330), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1196), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1208), .B(new_n928), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1188), .B(new_n1196), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(KEYINPUT57), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1033), .B1(new_n1205), .B2(new_n1214), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1204), .A2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n242), .A2(G41), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1038), .B(new_n1217), .C1(new_n344), .C2(new_n782), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n790), .A2(new_n464), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G68), .C2(new_n799), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n759), .A2(G58), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1220), .B(new_n1221), .C1(new_n1045), .C2(new_n763), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n784), .A2(G97), .B1(new_n593), .B2(new_n776), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT118), .Z(new_n1224));
  NOR2_X1   g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(KEYINPUT58), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(G33), .A2(G41), .ZN(new_n1227));
  OR3_X1    g1027(.A1(new_n1217), .A2(G50), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(KEYINPUT58), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1037), .A2(new_n1139), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n844), .A2(G128), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n846), .C2(new_n775), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G125), .B2(new_n768), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n1137), .B2(new_n847), .C1(new_n271), .C2(new_n800), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT59), .Z(new_n1235));
  NAND2_X1  g1035(.A1(new_n760), .A2(G124), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1227), .B(new_n1236), .C1(new_n758), .C2(new_n1008), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT119), .Z(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1226), .A2(new_n1228), .A3(new_n1229), .A4(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n750), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n748), .B1(new_n275), .B2(new_n858), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n1195), .C2(new_n806), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1200), .B2(new_n746), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1216), .A2(new_n1245), .ZN(G375));
  INV_X1    g1046(.A(new_n1161), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n975), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1155), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1201), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1247), .A2(new_n1248), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n916), .A2(new_n805), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n747), .B1(G68), .B2(new_n1127), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n764), .A2(G128), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n784), .A2(new_n1139), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n242), .B1(new_n782), .B2(new_n846), .C1(new_n1008), .C2(new_n780), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G132), .B2(new_n768), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1221), .A2(new_n1254), .A3(new_n1255), .A4(new_n1257), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n799), .A2(G50), .B1(G150), .B2(new_n776), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(KEYINPUT123), .Z(new_n1260));
  NAND2_X1  g1060(.A1(new_n795), .A2(G107), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n401), .B1(new_n782), .B2(new_n1045), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(G97), .B2(new_n1037), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G116), .A2(new_n784), .B1(new_n768), .B2(G294), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1261), .A2(new_n1035), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n322), .A2(new_n758), .B1(new_n763), .B2(new_n778), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1258), .A2(new_n1260), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1253), .B1(new_n1267), .B2(new_n750), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1155), .A2(new_n746), .B1(new_n1252), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1251), .A2(new_n1269), .ZN(G381));
  NOR2_X1   g1070(.A1(G393), .A2(G396), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1251), .A2(new_n861), .A3(new_n1269), .ZN(new_n1273));
  NOR4_X1   g1073(.A1(G387), .A2(new_n1272), .A3(G390), .A4(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(G375), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1149), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1147), .B1(new_n1276), .B2(new_n745), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1164), .A2(new_n1033), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1247), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1274), .A2(new_n1275), .A3(new_n1280), .ZN(G407));
  INV_X1    g1081(.A(G343), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(G213), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(KEYINPUT124), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1275), .A2(new_n1280), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(G407), .A2(new_n1285), .A3(G213), .ZN(G409));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G378), .B(new_n1245), .C1(new_n1204), .C2(new_n1215), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1200), .A2(new_n1203), .A3(new_n1248), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1212), .A2(new_n746), .A3(new_n1213), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1243), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1280), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1289), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT60), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1250), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1201), .A2(new_n1249), .A3(KEYINPUT60), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1296), .A2(new_n1033), .A3(new_n1247), .A4(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1269), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n861), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(G384), .A3(new_n1269), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  AND4_X1   g1102(.A1(new_n1288), .A2(new_n1294), .A3(new_n1283), .A4(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1283), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1289), .B2(new_n1293), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1288), .B1(new_n1305), .B2(new_n1302), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1287), .B1(new_n1303), .B2(new_n1306), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1305), .A2(KEYINPUT126), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1305), .A2(KEYINPUT126), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1300), .A2(new_n1301), .B1(G2897), .B2(new_n1284), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1304), .A2(G2897), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1302), .A2(new_n1311), .ZN(new_n1312));
  OAI22_X1  g1112(.A1(new_n1308), .A2(new_n1309), .B1(new_n1310), .B2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n823), .B1(new_n1034), .B2(new_n1070), .ZN(new_n1314));
  OR2_X1    g1114(.A1(new_n1271), .A2(new_n1314), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1004), .A2(G390), .A3(new_n1030), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G390), .B1(new_n1004), .B2(new_n1030), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1315), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(G390), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(G387), .A2(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1271), .A2(new_n1314), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1004), .A2(G390), .A3(new_n1030), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1318), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1284), .B1(new_n1289), .B2(new_n1293), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1326), .A2(KEYINPUT63), .A3(new_n1302), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1325), .B1(KEYINPUT127), .B2(new_n1327), .ZN(new_n1328));
  OR2_X1    g1128(.A1(new_n1327), .A2(KEYINPUT127), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1307), .A2(new_n1313), .A3(new_n1328), .A4(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1312), .A2(new_n1310), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1324), .B1(new_n1331), .B2(new_n1326), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1333), .B1(new_n1303), .B2(new_n1306), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1326), .A2(KEYINPUT62), .A3(new_n1302), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1332), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1318), .A2(new_n1323), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1330), .B1(new_n1336), .B2(new_n1338), .ZN(G405));
  NAND2_X1  g1139(.A1(G375), .A2(new_n1280), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1289), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1302), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1302), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1340), .A2(new_n1343), .A3(new_n1289), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1342), .A2(new_n1344), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1345), .B(new_n1337), .ZN(G402));
endmodule


