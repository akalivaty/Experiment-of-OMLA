//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  XNOR2_X1  g000(.A(G110), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n193), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  OAI21_X1  g010(.A(KEYINPUT3), .B1(new_n196), .B2(G107), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n198));
  INV_X1    g012(.A(G107), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(new_n199), .A3(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(G107), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(G101), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n195), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(G101), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n197), .A2(new_n200), .A3(new_n207), .A4(new_n201), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(KEYINPUT4), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT78), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT4), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n212), .B1(new_n202), .B2(G101), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT78), .A3(new_n208), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n205), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT83), .ZN(new_n216));
  AND3_X1   g030(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT5), .ZN(new_n217));
  OAI21_X1  g031(.A(G113), .B1(new_n190), .B2(KEYINPUT5), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G113), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n191), .A2(G119), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT5), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT5), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n223), .A2(KEYINPUT83), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n219), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n196), .A2(G107), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n199), .A2(G104), .ZN(new_n228));
  OAI21_X1  g042(.A(G101), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n208), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n193), .A2(new_n194), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n188), .B1(new_n215), .B2(new_n234), .ZN(new_n235));
  AND4_X1   g049(.A1(KEYINPUT78), .A2(new_n206), .A3(KEYINPUT4), .A4(new_n208), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT78), .B1(new_n213), .B2(new_n208), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n187), .B(new_n233), .C1(new_n238), .C2(new_n205), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(new_n239), .A3(KEYINPUT6), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT6), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n241), .B(new_n188), .C1(new_n215), .C2(new_n234), .ZN(new_n242));
  INV_X1    g056(.A(G146), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G143), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT67), .B(G128), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(G143), .B2(new_n243), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n247), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G125), .ZN(new_n252));
  XNOR2_X1  g066(.A(G143), .B(G146), .ZN(new_n253));
  INV_X1    g067(.A(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(KEYINPUT1), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n251), .A2(new_n252), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n244), .A2(new_n246), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT0), .B(G128), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n253), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G125), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G224), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G953), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n263), .B(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n240), .A2(new_n242), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT87), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n257), .A2(new_n262), .A3(KEYINPUT86), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT86), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n251), .A2(new_n256), .A3(new_n270), .A4(new_n252), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT7), .B1(new_n264), .B2(G953), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n268), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n263), .A2(new_n272), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n257), .A2(new_n262), .A3(KEYINPUT86), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n276), .A2(KEYINPUT87), .A3(new_n272), .A4(new_n271), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT85), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n224), .A2(KEYINPUT84), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT84), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n190), .A2(new_n192), .A3(new_n281), .A4(KEYINPUT5), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n282), .A3(new_n223), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n208), .A2(new_n229), .ZN(new_n284));
  INV_X1    g098(.A(new_n231), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n231), .B1(new_n219), .B2(new_n225), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(new_n284), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n187), .B(KEYINPUT8), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n279), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n279), .A3(new_n289), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n278), .A2(new_n239), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n267), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G210), .B1(G237), .B2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n267), .A2(new_n293), .A3(new_n294), .A4(new_n296), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  XOR2_X1   g115(.A(new_n301), .B(KEYINPUT81), .Z(new_n302));
  XOR2_X1   g116(.A(new_n302), .B(KEYINPUT82), .Z(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G122), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT90), .B1(new_n306), .B2(G116), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT90), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n191), .A3(G122), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n310), .B(new_n199), .C1(new_n191), .C2(G122), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT67), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G128), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n314), .A3(G143), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n245), .A2(G128), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G134), .ZN(new_n318));
  INV_X1    g132(.A(G134), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n315), .A2(new_n319), .A3(new_n316), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n310), .A2(KEYINPUT14), .B1(G116), .B2(new_n306), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT14), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n307), .A2(new_n309), .A3(new_n323), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n311), .B(new_n321), .C1(new_n325), .C2(new_n199), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n310), .B1(new_n191), .B2(G122), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G107), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n311), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT13), .B1(new_n245), .B2(G128), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT91), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT13), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n315), .B1(new_n332), .B2(new_n316), .ZN(new_n333));
  OAI21_X1  g147(.A(G134), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n329), .A2(new_n334), .A3(new_n320), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT9), .B(G234), .ZN(new_n336));
  INV_X1    g150(.A(G217), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n336), .A2(new_n337), .A3(G953), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n326), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT92), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT92), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n326), .A2(new_n335), .A3(new_n341), .A4(new_n338), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n326), .A2(new_n335), .ZN(new_n343));
  INV_X1    g157(.A(new_n338), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n340), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G478), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(KEYINPUT15), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n346), .A2(new_n294), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(new_n346), .B2(new_n294), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(G475), .A2(G902), .ZN(new_n353));
  INV_X1    g167(.A(G140), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G125), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n252), .A2(G140), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT72), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n354), .A2(KEYINPUT72), .A3(G125), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(KEYINPUT16), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT16), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n355), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G146), .ZN(new_n364));
  NOR2_X1   g178(.A1(G237), .A2(G953), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(G143), .A3(G214), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(G143), .B1(new_n365), .B2(G214), .ZN(new_n368));
  OAI21_X1  g182(.A(G131), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT17), .ZN(new_n370));
  INV_X1    g184(.A(G237), .ZN(new_n371));
  INV_X1    g185(.A(G953), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(G214), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n245), .ZN(new_n374));
  INV_X1    g188(.A(G131), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(new_n366), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n369), .A2(new_n370), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n360), .A2(new_n243), .A3(new_n362), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n375), .B1(new_n374), .B2(new_n366), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT17), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n364), .A2(new_n377), .A3(new_n378), .A4(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G113), .B(G122), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(new_n196), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n358), .A2(G146), .A3(new_n359), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n355), .A2(new_n356), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n243), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(KEYINPUT18), .A2(G131), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n374), .A2(new_n366), .A3(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(KEYINPUT18), .B(G131), .C1(new_n367), .C2(new_n368), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n381), .A2(new_n383), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT88), .ZN(new_n393));
  INV_X1    g207(.A(new_n376), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(new_n379), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT19), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(new_n358), .B2(new_n359), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n385), .A2(KEYINPUT19), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n243), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n369), .A2(KEYINPUT88), .A3(new_n376), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n395), .A2(new_n364), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n383), .B1(new_n401), .B2(new_n391), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n353), .B1(new_n392), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT20), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT89), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT89), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n406), .A3(KEYINPUT20), .ZN(new_n407));
  OR2_X1    g221(.A1(new_n392), .A2(new_n402), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n353), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n405), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G475), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n383), .B1(new_n381), .B2(new_n391), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n392), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n412), .B1(new_n414), .B2(new_n294), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(G234), .A2(G237), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(G952), .A3(new_n372), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(G902), .A3(G953), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(G898), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n352), .A2(new_n411), .A3(new_n416), .A4(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G221), .B1(new_n336), .B2(G902), .ZN(new_n426));
  XOR2_X1   g240(.A(new_n426), .B(KEYINPUT77), .Z(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G110), .B(G140), .ZN(new_n429));
  INV_X1    g243(.A(G227), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G953), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n429), .B(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n261), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n204), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n211), .B2(new_n214), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT1), .B1(new_n245), .B2(G146), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n436), .A2(G128), .B1(new_n244), .B2(new_n246), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n255), .A2(new_n244), .A3(new_n246), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n208), .B(new_n229), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT10), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n440), .B1(new_n251), .B2(new_n256), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(new_n284), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  AND2_X1   g258(.A1(KEYINPUT11), .A2(G134), .ZN(new_n445));
  OR2_X1    g259(.A1(KEYINPUT11), .A2(G134), .ZN(new_n446));
  INV_X1    g260(.A(G137), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AND2_X1   g263(.A1(KEYINPUT65), .A2(G137), .ZN(new_n450));
  NOR2_X1   g264(.A1(KEYINPUT65), .A2(G137), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT66), .B1(new_n452), .B2(new_n445), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n447), .ZN(new_n455));
  NAND2_X1  g269(.A1(KEYINPUT65), .A2(G137), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n445), .A3(KEYINPUT66), .A4(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n449), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G131), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(new_n456), .A3(new_n445), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n457), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n375), .A3(new_n449), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  NOR3_X1   g280(.A1(new_n435), .A2(new_n444), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n375), .B1(new_n464), .B2(new_n449), .ZN(new_n468));
  AOI211_X1 g282(.A(G131), .B(new_n448), .C1(new_n463), .C2(new_n457), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n433), .A2(new_n204), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n236), .B2(new_n237), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n440), .A2(new_n439), .B1(new_n442), .B2(new_n284), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n432), .B1(new_n467), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT12), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n476), .A2(KEYINPUT80), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(KEYINPUT80), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n230), .A2(new_n251), .A3(new_n256), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n479), .A2(new_n439), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n477), .B(new_n478), .C1(new_n470), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n472), .A2(new_n470), .A3(new_n473), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n439), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n466), .A2(KEYINPUT80), .A3(new_n476), .A4(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n432), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n481), .A2(new_n482), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n475), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G469), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(new_n294), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n294), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n432), .ZN(new_n494));
  INV_X1    g308(.A(new_n474), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n482), .A3(new_n485), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(new_n488), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n428), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n305), .A2(new_n425), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT22), .B(G137), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n372), .A2(G221), .A3(G234), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n501), .B(new_n502), .Z(new_n503));
  INV_X1    g317(.A(KEYINPUT75), .ZN(new_n504));
  INV_X1    g318(.A(G110), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT24), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G110), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT71), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n506), .B2(new_n508), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n254), .A2(G119), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(new_n248), .B2(G119), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT23), .B1(new_n254), .B2(G119), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(new_n513), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT23), .A4(G119), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n512), .A2(new_n514), .B1(new_n518), .B2(G110), .ZN(new_n519));
  INV_X1    g333(.A(new_n378), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n243), .B1(new_n360), .B2(new_n362), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT73), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT73), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n519), .B(new_n524), .C1(new_n520), .C2(new_n521), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT74), .B(G110), .Z(new_n527));
  NAND3_X1  g341(.A1(new_n516), .A2(new_n517), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n512), .B2(new_n514), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n364), .A2(new_n529), .A3(new_n386), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n504), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  AOI211_X1 g346(.A(KEYINPUT75), .B(new_n530), .C1(new_n523), .C2(new_n525), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n503), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n503), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n526), .A2(new_n531), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(KEYINPUT75), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n337), .B1(G234), .B2(new_n294), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(G902), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n534), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT76), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n534), .A2(KEYINPUT76), .A3(new_n537), .A4(new_n539), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n534), .A2(new_n545), .A3(new_n294), .A4(new_n537), .ZN(new_n546));
  INV_X1    g360(.A(new_n538), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n534), .A2(new_n294), .A3(new_n537), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n547), .B1(new_n548), .B2(KEYINPUT25), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n544), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n433), .B1(new_n468), .B2(new_n469), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT68), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(G131), .B1(new_n319), .B2(new_n447), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n452), .B2(new_n319), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n251), .B2(new_n256), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n465), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(KEYINPUT68), .B(new_n433), .C1(new_n468), .C2(new_n469), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n553), .A2(KEYINPUT30), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n261), .B(KEYINPUT64), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n557), .B1(new_n470), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n559), .A2(new_n195), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n195), .B1(new_n465), .B2(new_n556), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n553), .A2(new_n565), .A3(new_n558), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT69), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n365), .A2(G210), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT27), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT26), .B(G101), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n566), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n567), .B1(new_n566), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n564), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT31), .ZN(new_n575));
  INV_X1    g389(.A(new_n571), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT28), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n561), .A2(new_n195), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n577), .B1(new_n566), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT28), .B1(new_n551), .B2(new_n565), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n576), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT70), .B(KEYINPUT31), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n564), .B(new_n582), .C1(new_n572), .C2(new_n573), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n575), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT32), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n585), .A2(G472), .A3(G902), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n579), .A2(new_n580), .A3(new_n576), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n571), .B1(new_n564), .B2(new_n566), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT29), .ZN(new_n590));
  INV_X1    g404(.A(new_n580), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT29), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n576), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT68), .B1(new_n466), .B2(new_n433), .ZN(new_n594));
  INV_X1    g408(.A(new_n558), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n553), .A2(new_n557), .A3(new_n558), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n565), .A2(new_n596), .B1(new_n597), .B2(new_n195), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n591), .B(new_n593), .C1(new_n598), .C2(new_n577), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n294), .ZN(new_n600));
  OAI21_X1  g414(.A(G472), .B1(new_n590), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n587), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(G472), .A2(G902), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT32), .B1(new_n584), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n500), .B(new_n550), .C1(new_n602), .C2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  NAND2_X1  g420(.A1(new_n584), .A2(new_n294), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n607), .A2(G472), .B1(new_n603), .B2(new_n584), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n548), .A2(KEYINPUT25), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(new_n546), .A3(new_n538), .ZN(new_n610));
  AOI21_X1  g424(.A(G902), .B1(new_n475), .B2(new_n486), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n490), .B1(new_n611), .B2(new_n488), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n467), .A2(new_n432), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n613), .A2(new_n495), .B1(new_n493), .B2(new_n432), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G469), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n427), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  AND4_X1   g430(.A1(new_n610), .A2(new_n542), .A3(new_n543), .A4(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n608), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n346), .A2(new_n294), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n347), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n345), .A2(KEYINPUT33), .A3(new_n339), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n621), .A2(KEYINPUT93), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT33), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n346), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n621), .A2(KEYINPUT93), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n294), .A2(G478), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n620), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n411), .A2(new_n416), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n302), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n288), .A2(new_n279), .A3(new_n289), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n632), .A2(new_n633), .A3(new_n290), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n634), .B2(new_n239), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n296), .B1(new_n635), .B2(new_n267), .ZN(new_n636));
  INV_X1    g450(.A(new_n299), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n631), .B(new_n424), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n630), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n618), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  INV_X1    g456(.A(new_n410), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT94), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n403), .A2(new_n406), .A3(KEYINPUT20), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n406), .B1(new_n403), .B2(KEYINPUT20), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n405), .A2(KEYINPUT94), .A3(new_n407), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n643), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT95), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n416), .B1(new_n350), .B2(new_n351), .ZN(new_n651));
  NOR4_X1   g465(.A1(new_n638), .A2(new_n649), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n647), .A2(new_n648), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n651), .B1(new_n653), .B2(new_n410), .ZN(new_n654));
  AOI211_X1 g468(.A(new_n302), .B(new_n423), .C1(new_n298), .C2(new_n299), .ZN(new_n655));
  AOI21_X1  g469(.A(KEYINPUT95), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n618), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(KEYINPUT96), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT97), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT35), .B(G107), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  NOR2_X1   g477(.A1(new_n305), .A2(new_n425), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n535), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n536), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n539), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n499), .B1(new_n610), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n608), .A2(new_n664), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT37), .B(G110), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT98), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n669), .B(new_n671), .ZN(G12));
  AOI21_X1  g486(.A(new_n302), .B1(new_n298), .B2(new_n299), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n564), .A2(new_n566), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n576), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n566), .A2(new_n578), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n591), .B(new_n571), .C1(new_n677), .C2(new_n577), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n676), .A2(new_n678), .A3(new_n592), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n294), .A3(new_n599), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n680), .A2(G472), .B1(new_n584), .B2(new_n586), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n584), .A2(new_n603), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n585), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n674), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT99), .B(G900), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n421), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n418), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n649), .A2(new_n651), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n684), .A2(new_n668), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT100), .B(G128), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G30));
  NAND2_X1  g506(.A1(new_n597), .A2(new_n195), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n566), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n576), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n574), .A2(KEYINPUT101), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n294), .ZN(new_n697));
  AOI21_X1  g511(.A(KEYINPUT101), .B1(new_n574), .B2(new_n695), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n683), .A2(new_n587), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT102), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n300), .B(KEYINPUT38), .ZN(new_n702));
  OR2_X1    g516(.A1(new_n350), .A2(new_n351), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n629), .A2(new_n631), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n610), .A2(new_n667), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n687), .B(KEYINPUT39), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n616), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(KEYINPUT40), .Z(new_n709));
  NAND4_X1  g523(.A1(new_n701), .A2(new_n702), .A3(new_n706), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G143), .ZN(G45));
  NOR2_X1   g525(.A1(new_n630), .A2(new_n688), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n684), .A2(new_n668), .A3(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT103), .B(G146), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G48));
  AOI21_X1  g529(.A(new_n488), .B1(new_n487), .B2(new_n294), .ZN(new_n716));
  AOI211_X1 g530(.A(G469), .B(G902), .C1(new_n475), .C2(new_n486), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n426), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n550), .B(new_n721), .C1(new_n602), .C2(new_n604), .ZN(new_n722));
  INV_X1    g536(.A(new_n639), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT41), .B(G113), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G15));
  NOR2_X1   g540(.A1(new_n657), .A2(new_n722), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n191), .ZN(G18));
  AND3_X1   g542(.A1(new_n673), .A2(new_n426), .A3(new_n718), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n425), .B1(new_n610), .B2(new_n667), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n729), .B(new_n730), .C1(new_n602), .C2(new_n604), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  NAND4_X1  g546(.A1(new_n629), .A2(new_n718), .A3(new_n703), .A4(new_n426), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n638), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n607), .A2(G472), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n580), .B1(new_n694), .B2(KEYINPUT28), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n575), .B(new_n583), .C1(new_n571), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n603), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n734), .A2(new_n550), .A3(new_n735), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G122), .ZN(G24));
  AOI22_X1  g554(.A1(new_n607), .A2(G472), .B1(new_n603), .B2(new_n737), .ZN(new_n741));
  AND3_X1   g555(.A1(new_n741), .A2(new_n705), .A3(new_n712), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT104), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n729), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n741), .A2(new_n705), .A3(new_n712), .ZN(new_n745));
  INV_X1    g559(.A(new_n729), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT104), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G125), .ZN(G27));
  NAND2_X1  g563(.A1(new_n681), .A2(new_n683), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT105), .B1(new_n614), .B2(G469), .ZN(new_n751));
  AND4_X1   g565(.A1(KEYINPUT105), .A2(new_n494), .A3(G469), .A4(new_n496), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n720), .B1(new_n753), .B2(new_n612), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n298), .A2(new_n755), .A3(new_n299), .A4(new_n631), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n298), .A2(new_n299), .A3(new_n631), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT106), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n754), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n750), .A2(new_n759), .A3(new_n550), .A4(new_n712), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n610), .A2(new_n542), .A3(new_n543), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n681), .B2(new_n683), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(KEYINPUT42), .A3(new_n712), .A4(new_n759), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT107), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n762), .A2(new_n768), .A3(new_n765), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n375), .ZN(G33));
  NAND3_X1  g585(.A1(new_n764), .A2(new_n689), .A3(new_n759), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  NAND2_X1  g587(.A1(new_n758), .A2(new_n756), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n628), .A2(new_n411), .A3(new_n416), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT43), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n778), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n608), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n780), .A2(new_n781), .A3(new_n705), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n774), .B1(new_n782), .B2(KEYINPUT44), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n488), .B1(new_n497), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(new_n784), .B2(new_n497), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(KEYINPUT46), .A3(new_n491), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(KEYINPUT108), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT46), .B1(new_n786), .B2(new_n491), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n717), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n720), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(new_n707), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n783), .B(new_n792), .C1(KEYINPUT44), .C2(new_n782), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  NAND2_X1  g608(.A1(new_n712), .A2(new_n763), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n795), .A2(new_n750), .A3(new_n774), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n791), .A2(KEYINPUT47), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n791), .A2(KEYINPUT47), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  NOR3_X1   g614(.A1(new_n775), .A2(new_n303), .A3(new_n427), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n718), .B(KEYINPUT49), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n550), .A3(new_n802), .ZN(new_n803));
  OR3_X1    g617(.A1(new_n701), .A2(new_n702), .A3(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n780), .A2(new_n419), .ZN(new_n805));
  INV_X1    g619(.A(new_n774), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(new_n721), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n764), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(KEYINPUT48), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n805), .A2(new_n550), .A3(new_n741), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n746), .ZN(new_n812));
  INV_X1    g626(.A(G952), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n812), .A2(new_n813), .A3(G953), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n806), .A2(new_n550), .A3(new_n419), .A4(new_n721), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n701), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n810), .B(new_n814), .C1(new_n630), .C2(new_n816), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n817), .B(KEYINPUT116), .Z(new_n818));
  NOR3_X1   g632(.A1(new_n816), .A2(new_n629), .A3(new_n628), .ZN(new_n819));
  INV_X1    g633(.A(new_n721), .ZN(new_n820));
  OR4_X1    g634(.A1(new_n631), .A2(new_n811), .A3(new_n702), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(KEYINPUT115), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT50), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n819), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n821), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n808), .A2(new_n705), .A3(new_n741), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n797), .A2(new_n798), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n718), .A2(new_n427), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n774), .B(new_n811), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  OR3_X1    g645(.A1(new_n827), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n828), .B1(new_n827), .B2(new_n831), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n818), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n653), .A2(new_n410), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n415), .A2(new_n688), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(KEYINPUT110), .A3(new_n352), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT110), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n352), .A2(new_n836), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n838), .B1(new_n649), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n750), .A3(new_n668), .A4(new_n806), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n759), .A2(new_n705), .A3(new_n741), .A4(new_n712), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n772), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n605), .B(new_n669), .C1(new_n722), .C2(new_n723), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n304), .B(new_n424), .C1(new_n636), .C2(new_n637), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n703), .A2(new_n411), .A3(new_n416), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n846), .B1(new_n630), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n608), .A2(new_n617), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n731), .A3(new_n739), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n844), .A2(new_n845), .A3(new_n727), .A4(new_n850), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n684), .B(new_n668), .C1(new_n689), .C2(new_n712), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n673), .A2(new_n629), .A3(new_n703), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(new_n754), .ZN(new_n855));
  INV_X1    g669(.A(new_n705), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n856), .A2(KEYINPUT112), .A3(new_n687), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT112), .B1(new_n856), .B2(new_n687), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n700), .B(new_n855), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n747), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n745), .A2(KEYINPUT104), .A3(new_n746), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n852), .B(new_n859), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(KEYINPUT113), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n748), .A2(new_n852), .A3(new_n859), .A4(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n868), .B1(new_n762), .B2(new_n765), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n851), .A2(new_n865), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n845), .A2(new_n727), .A3(new_n850), .ZN(new_n871));
  INV_X1    g685(.A(new_n844), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n767), .A2(new_n871), .A3(new_n769), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT111), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT111), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n851), .A2(new_n875), .A3(new_n767), .A4(new_n769), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n862), .A2(new_n863), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n748), .A2(KEYINPUT52), .A3(new_n852), .A4(new_n859), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n874), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n870), .B1(new_n880), .B2(new_n868), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n880), .A2(KEYINPUT53), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n865), .A2(new_n867), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(new_n874), .A3(new_n868), .A4(new_n876), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(KEYINPUT54), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n883), .A2(KEYINPUT114), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT114), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n884), .A2(new_n889), .A3(KEYINPUT54), .A4(new_n886), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n834), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(G952), .A2(G953), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n804), .B1(new_n891), .B2(new_n892), .ZN(G75));
  NOR2_X1   g707(.A1(new_n372), .A2(G952), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n881), .A2(new_n294), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT56), .B1(new_n896), .B2(G210), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n240), .A2(new_n242), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(new_n266), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT55), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n895), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n897), .B2(new_n900), .ZN(G51));
  NAND2_X1  g716(.A1(new_n880), .A2(new_n868), .ZN(new_n903));
  INV_X1    g717(.A(new_n870), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT54), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT117), .B1(new_n881), .B2(new_n882), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n905), .A2(KEYINPUT117), .A3(KEYINPUT54), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n490), .B(KEYINPUT57), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n487), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n881), .A2(new_n294), .A3(new_n786), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n894), .B1(new_n912), .B2(new_n913), .ZN(G54));
  INV_X1    g728(.A(KEYINPUT58), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n915), .A2(new_n412), .A3(KEYINPUT118), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT118), .B1(new_n915), .B2(new_n412), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n896), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n408), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n920), .A2(new_n921), .A3(new_n894), .ZN(G60));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT59), .Z(new_n924));
  NOR2_X1   g738(.A1(new_n626), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n908), .A2(new_n909), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT119), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n926), .A2(new_n927), .A3(new_n895), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n927), .B1(new_n926), .B2(new_n895), .ZN(new_n929));
  INV_X1    g743(.A(new_n924), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n888), .A2(new_n890), .A3(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n931), .A2(new_n626), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n928), .A2(new_n929), .A3(new_n932), .ZN(G63));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n934), .A2(KEYINPUT121), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT120), .ZN(new_n936));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT60), .ZN(new_n938));
  INV_X1    g752(.A(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n905), .A2(new_n936), .A3(new_n666), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n534), .A2(new_n537), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n881), .B2(new_n938), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n895), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n881), .A2(new_n938), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n936), .B1(new_n944), .B2(new_n666), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n935), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n934), .A2(KEYINPUT121), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(G66));
  NOR2_X1   g762(.A1(new_n871), .A2(G953), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT122), .ZN(new_n950));
  OAI21_X1  g764(.A(G953), .B1(new_n422), .B2(new_n264), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n898), .B1(G898), .B2(new_n372), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G69));
  INV_X1    g768(.A(G900), .ZN(new_n955));
  OAI21_X1  g769(.A(G953), .B1(new_n430), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT125), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n559), .A2(new_n563), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n397), .A2(new_n398), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n748), .A2(new_n852), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n710), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(KEYINPUT123), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT123), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n969), .A3(KEYINPUT62), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n793), .A2(new_n799), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n708), .B1(new_n630), .B2(new_n847), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n764), .A2(new_n806), .A3(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n971), .A2(new_n972), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n964), .B1(new_n977), .B2(new_n372), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n792), .A2(new_n764), .A3(new_n854), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n965), .A2(new_n772), .A3(new_n980), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n981), .A2(new_n973), .A3(new_n770), .ZN(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n983), .A2(G953), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n964), .B1(new_n955), .B2(new_n372), .ZN(new_n985));
  OAI22_X1  g799(.A1(new_n978), .A2(new_n979), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n974), .B(new_n976), .C1(KEYINPUT62), .C2(new_n966), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n970), .B2(new_n968), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n963), .B1(new_n988), .B2(G953), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(KEYINPUT124), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n959), .B(new_n960), .C1(new_n986), .C2(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n984), .A2(new_n985), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n989), .B2(KEYINPUT124), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n978), .A2(new_n979), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n993), .A2(new_n994), .A3(KEYINPUT126), .A4(new_n958), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n991), .A2(new_n995), .ZN(G72));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  INV_X1    g812(.A(new_n871), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n998), .B1(new_n977), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n1000), .A2(new_n571), .A3(new_n675), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n574), .B1(new_n589), .B2(KEYINPUT127), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n589), .A2(KEYINPUT127), .ZN(new_n1003));
  OR2_X1    g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n884), .A2(new_n886), .A3(new_n998), .A4(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n998), .B1(new_n983), .B2(new_n999), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n675), .A2(new_n571), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n894), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1001), .A2(new_n1005), .A3(new_n1008), .ZN(G57));
endmodule


