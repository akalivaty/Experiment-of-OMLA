//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n569, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT67), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT66), .B1(new_n469), .B2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(new_n461), .B(new_n468), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n464), .B1(new_n465), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n475), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n461), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n473), .A2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n479), .B1(new_n474), .B2(KEYINPUT66), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(G2105), .A3(new_n468), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  INV_X1    g058(.A(new_n472), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(KEYINPUT68), .C1(G114), .C2(new_n461), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n461), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(new_n490), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n480), .A2(G126), .A3(G2105), .A4(new_n468), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n472), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n469), .A2(G2104), .ZN(new_n503));
  AND4_X1   g078(.A1(new_n461), .A2(new_n502), .A3(new_n479), .A4(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n498), .A2(new_n499), .A3(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n480), .A2(G138), .A3(new_n461), .A4(new_n468), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n504), .B1(new_n508), .B2(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n496), .A2(new_n497), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT69), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n511), .ZN(G164));
  AND2_X1   g087(.A1(KEYINPUT70), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT70), .A2(G651), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT6), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g092(.A(KEYINPUT71), .B(KEYINPUT6), .C1(new_n513), .C2(new_n514), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT72), .B1(new_n519), .B2(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n521), .A2(new_n522), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(KEYINPUT73), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(KEYINPUT5), .A3(G543), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n517), .A2(new_n518), .A3(new_n524), .A4(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G88), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n513), .A2(new_n514), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n530), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n531), .A2(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n517), .A2(G543), .A3(new_n518), .A4(new_n524), .ZN(new_n537));
  INV_X1    g112(.A(G50), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G166));
  NAND3_X1  g115(.A1(new_n530), .A2(G63), .A3(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT7), .ZN(new_n543));
  INV_X1    g118(.A(G51), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n541), .B(new_n543), .C1(new_n537), .C2(new_n544), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT74), .B(G89), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n531), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G168));
  INV_X1    g124(.A(G64), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n527), .B2(new_n529), .ZN(new_n551));
  AND2_X1   g126(.A1(G77), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n533), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(G90), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n531), .B2(new_n554), .ZN(new_n555));
  XOR2_X1   g130(.A(KEYINPUT75), .B(G52), .Z(new_n556));
  NOR2_X1   g131(.A1(new_n537), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(G171));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(new_n527), .B2(new_n529), .ZN(new_n560));
  AND2_X1   g135(.A1(G68), .A2(G543), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n533), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G43), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n537), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G81), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n531), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  AND3_X1   g143(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G36), .ZN(G176));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT8), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(G188));
  AND2_X1   g148(.A1(new_n530), .A2(G65), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT77), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n531), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G91), .ZN(new_n579));
  NOR2_X1   g154(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n580));
  INV_X1    g155(.A(new_n537), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(G53), .ZN(new_n582));
  INV_X1    g157(.A(G53), .ZN(new_n583));
  XOR2_X1   g158(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n584));
  NOR3_X1   g159(.A1(new_n537), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n577), .B(new_n579), .C1(new_n582), .C2(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  OR2_X1    g162(.A1(new_n545), .A2(new_n548), .ZN(G286));
  OR2_X1    g163(.A1(new_n536), .A2(new_n539), .ZN(G303));
  OAI21_X1  g164(.A(G651), .B1(new_n530), .B2(G74), .ZN(new_n590));
  INV_X1    g165(.A(G87), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n531), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G49), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n537), .A2(new_n593), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n592), .A2(new_n594), .ZN(G288));
  AOI22_X1  g170(.A1(new_n530), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n534), .ZN(new_n597));
  INV_X1    g172(.A(G86), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n531), .ZN(new_n599));
  INV_X1    g174(.A(G48), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n537), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G305));
  AND2_X1   g178(.A1(new_n578), .A2(G85), .ZN(new_n604));
  INV_X1    g179(.A(G47), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n530), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n537), .A2(new_n605), .B1(new_n534), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  AND3_X1   g185(.A1(new_n517), .A2(new_n518), .A3(new_n524), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n612));
  NAND4_X1  g187(.A1(new_n611), .A2(new_n612), .A3(G92), .A4(new_n530), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT78), .B1(new_n531), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT10), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT79), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n530), .A2(G66), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n519), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(new_n581), .B2(G54), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n615), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n618), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n610), .B1(new_n626), .B2(G868), .ZN(G284));
  OAI21_X1  g202(.A(new_n610), .B1(new_n626), .B2(G868), .ZN(G321));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  INV_X1    g204(.A(G299), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G868), .ZN(G280));
  XOR2_X1   g206(.A(G280), .B(KEYINPUT80), .Z(G297));
  INV_X1    g207(.A(G559), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n626), .B1(new_n633), .B2(G860), .ZN(G148));
  NAND2_X1  g209(.A1(new_n626), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G868), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(KEYINPUT81), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(KEYINPUT81), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n637), .B(new_n638), .C1(G868), .C2(new_n567), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT82), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n463), .A2(new_n475), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT12), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2100), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n482), .A2(G123), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n484), .A2(G135), .ZN(new_n647));
  OR2_X1    g222(.A1(G99), .A2(G2105), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n648), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(G2096), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n645), .A2(new_n651), .ZN(G156));
  XOR2_X1   g227(.A(KEYINPUT15), .B(G2435), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2438), .ZN(new_n654));
  XOR2_X1   g229(.A(G2427), .B(G2430), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT83), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT14), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2446), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n658), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT84), .B(KEYINPUT85), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT16), .B(G2443), .Z(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(G14), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(G401));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT86), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  NOR2_X1   g248(.A1(G2072), .A2(G2078), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n672), .B(new_n673), .C1(new_n443), .C2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n672), .A2(new_n673), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n443), .A2(new_n674), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT17), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n681), .B(KEYINPUT88), .Z(new_n684));
  OAI211_X1 g259(.A(new_n677), .B(new_n683), .C1(new_n679), .C2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2096), .B(G2100), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT19), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n689), .A2(new_n690), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n692), .A2(new_n694), .A3(new_n696), .ZN(new_n700));
  OAI211_X1 g275(.A(new_n699), .B(new_n700), .C1(new_n698), .C2(new_n697), .ZN(new_n701));
  XOR2_X1   g276(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1991), .B(G1996), .ZN(new_n704));
  INV_X1    g279(.A(G1981), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n703), .B(new_n707), .ZN(G229));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G23), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n592), .A2(new_n594), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT33), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1976), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n709), .A2(G6), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n602), .B2(new_n709), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT32), .B(G1981), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G16), .A2(G22), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G166), .B2(G16), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1971), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  AND3_X1   g298(.A1(new_n714), .A2(new_n715), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n715), .B1(new_n714), .B2(new_n723), .ZN(new_n726));
  NOR3_X1   g301(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G25), .ZN(new_n729));
  OR2_X1    g304(.A1(G95), .A2(G2105), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n730), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n731));
  INV_X1    g306(.A(G131), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n472), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G119), .B2(new_n482), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n729), .B1(new_n734), .B2(new_n728), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(G16), .A2(G24), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n608), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT89), .ZN(new_n740));
  INV_X1    g315(.A(G1986), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n727), .A2(new_n737), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT31), .B(G11), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n743), .A2(new_n744), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n709), .A2(KEYINPUT23), .A3(G20), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT23), .ZN(new_n749));
  INV_X1    g324(.A(G20), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n750), .B2(G16), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n748), .B(new_n751), .C1(new_n630), .C2(new_n709), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G1956), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT91), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G29), .B2(G33), .ZN(new_n755));
  OR3_X1    g330(.A1(new_n754), .A2(G29), .A3(G33), .ZN(new_n756));
  AOI22_X1  g331(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n757), .A2(new_n461), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G139), .B2(new_n484), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT25), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g338(.A(new_n755), .B(new_n756), .C1(new_n763), .C2(new_n728), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G2072), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n728), .A2(G27), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G164), .B2(new_n728), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n765), .B1(new_n767), .B2(G2078), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n753), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n626), .A2(G16), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G4), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G1348), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n771), .A2(new_n772), .B1(G2078), .B2(new_n767), .ZN(new_n773));
  NOR2_X1   g348(.A1(G29), .A2(G35), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G162), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT29), .B(G2090), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G16), .A2(G19), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n567), .B2(G16), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n777), .B1(G1341), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n728), .A2(G26), .ZN(new_n781));
  OR2_X1    g356(.A1(G104), .A2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n782), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n783));
  INV_X1    g358(.A(G140), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n472), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G128), .B2(new_n482), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n781), .B1(new_n786), .B2(new_n728), .ZN(new_n787));
  MUX2_X1   g362(.A(new_n781), .B(new_n787), .S(KEYINPUT28), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2067), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n779), .A2(G1341), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n650), .A2(new_n728), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT95), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n769), .A2(new_n773), .A3(new_n780), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G5), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G171), .B2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT97), .B(G1961), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT94), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G16), .B2(G21), .ZN(new_n800));
  NAND2_X1  g375(.A1(G168), .A2(G16), .ZN(new_n801));
  MUX2_X1   g376(.A(new_n799), .B(new_n800), .S(new_n801), .Z(new_n802));
  INV_X1    g377(.A(G1966), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n798), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT96), .B(KEYINPUT30), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G28), .ZN(new_n807));
  OAI22_X1  g382(.A1(new_n771), .A2(new_n772), .B1(G29), .B2(new_n807), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n794), .A2(new_n804), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n482), .A2(G129), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n463), .A2(G105), .ZN(new_n812));
  NAND3_X1  g387(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT26), .Z(new_n814));
  NAND2_X1  g389(.A1(new_n484), .A2(G141), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n811), .A2(new_n812), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT92), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT93), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(G29), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G29), .B2(G32), .ZN(new_n823));
  XOR2_X1   g398(.A(KEYINPUT27), .B(G1996), .Z(new_n824));
  XOR2_X1   g399(.A(new_n823), .B(new_n824), .Z(new_n825));
  OR2_X1    g400(.A1(KEYINPUT24), .A2(G34), .ZN(new_n826));
  NAND2_X1  g401(.A1(KEYINPUT24), .A2(G34), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n826), .A2(new_n728), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G160), .B2(new_n728), .ZN(new_n829));
  INV_X1    g404(.A(G2084), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n810), .A2(new_n825), .A3(new_n832), .ZN(G311));
  AND3_X1   g408(.A1(new_n745), .A2(new_n747), .A3(new_n809), .ZN(new_n834));
  INV_X1    g409(.A(new_n825), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n834), .A2(new_n835), .A3(new_n831), .A4(new_n746), .ZN(G150));
  INV_X1    g411(.A(G67), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n527), .B2(new_n529), .ZN(new_n838));
  AND2_X1   g413(.A1(G80), .A2(G543), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n533), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G55), .ZN(new_n841));
  INV_X1    g416(.A(G93), .ZN(new_n842));
  OAI221_X1 g417(.A(new_n840), .B1(new_n537), .B2(new_n841), .C1(new_n842), .C2(new_n531), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT98), .B(G860), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NOR2_X1   g421(.A1(new_n625), .A2(new_n633), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n843), .A2(new_n567), .ZN(new_n849));
  OAI221_X1 g424(.A(new_n562), .B1(new_n537), .B2(new_n563), .C1(new_n565), .C2(new_n531), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n840), .B1(new_n537), .B2(new_n841), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n531), .A2(new_n842), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT39), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n848), .B(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n846), .B1(new_n857), .B2(new_n844), .ZN(G145));
  NOR2_X1   g433(.A1(new_n509), .A2(new_n510), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n734), .ZN(new_n860));
  XNOR2_X1  g435(.A(G160), .B(KEYINPUT99), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n488), .ZN(new_n862));
  INV_X1    g437(.A(new_n650), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n862), .A2(new_n863), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n860), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n862), .A2(new_n863), .ZN(new_n868));
  INV_X1    g443(.A(new_n860), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n864), .A3(new_n869), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n643), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n763), .B1(new_n819), .B2(new_n820), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n817), .A2(new_n763), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n872), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n873), .A2(new_n872), .A3(new_n875), .ZN(new_n878));
  INV_X1    g453(.A(new_n786), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n484), .A2(G142), .ZN(new_n880));
  INV_X1    g455(.A(G130), .ZN(new_n881));
  OAI21_X1  g456(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n461), .A2(G118), .ZN(new_n883));
  OAI221_X1 g458(.A(new_n880), .B1(new_n881), .B2(new_n481), .C1(new_n882), .C2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n879), .B(new_n884), .ZN(new_n885));
  NOR3_X1   g460(.A1(new_n877), .A2(new_n878), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  INV_X1    g462(.A(new_n873), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(new_n643), .A3(new_n874), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n889), .B2(new_n876), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n871), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n885), .B1(new_n877), .B2(new_n878), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n867), .A2(new_n870), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n876), .A3(new_n887), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT100), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n891), .A2(new_n895), .A3(new_n899), .A4(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g477(.A1(G303), .A2(G288), .ZN(new_n903));
  NAND2_X1  g478(.A1(G166), .A2(new_n711), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n903), .A2(G305), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(G305), .B1(new_n903), .B2(new_n904), .ZN(new_n906));
  OR3_X1    g481(.A1(new_n905), .A2(new_n906), .A3(G290), .ZN(new_n907));
  OAI21_X1  g482(.A(G290), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n635), .B(new_n855), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n613), .A2(KEYINPUT10), .A3(new_n615), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT10), .B1(new_n613), .B2(new_n615), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(G299), .A3(new_n623), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n625), .A2(new_n630), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(G299), .B1(new_n915), .B2(new_n623), .ZN(new_n922));
  AND4_X1   g497(.A1(G299), .A2(new_n618), .A3(new_n623), .A4(new_n624), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT101), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT101), .B1(new_n625), .B2(new_n630), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n921), .B1(new_n927), .B2(new_n920), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n919), .B1(new_n928), .B2(new_n912), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n911), .B(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(G868), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(G868), .B2(new_n853), .ZN(G295));
  OAI21_X1  g507(.A(new_n931), .B1(G868), .B2(new_n853), .ZN(G331));
  NOR2_X1   g508(.A1(new_n922), .A2(new_n923), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n925), .B1(new_n918), .B2(KEYINPUT101), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n578), .A2(G90), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n537), .A2(new_n556), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .A4(new_n553), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT103), .B1(new_n555), .B2(new_n557), .ZN(new_n941));
  NAND3_X1  g516(.A1(G286), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(G168), .A2(new_n939), .A3(G171), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n855), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n849), .A2(new_n854), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n946), .A2(new_n942), .A3(new_n943), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n936), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n947), .A2(new_n936), .ZN(new_n949));
  OAI22_X1  g524(.A1(new_n935), .A2(new_n920), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n946), .A2(new_n942), .A3(new_n943), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n946), .B1(new_n943), .B2(new_n942), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n934), .B1(new_n950), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n935), .B(KEYINPUT41), .C1(new_n948), .C2(new_n949), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n909), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n948), .A2(new_n949), .A3(new_n934), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n934), .A2(KEYINPUT41), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n935), .B2(KEYINPUT41), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n961), .B2(new_n954), .ZN(new_n962));
  INV_X1    g537(.A(new_n909), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n958), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT104), .B1(new_n951), .B2(new_n952), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n947), .A2(new_n936), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n918), .A3(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n928), .B2(new_n953), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n909), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n964), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n966), .B1(new_n972), .B2(new_n965), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n976));
  AOI22_X1  g551(.A1(new_n927), .A2(KEYINPUT41), .B1(new_n967), .B2(new_n968), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n918), .B1(new_n977), .B2(new_n953), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n963), .B1(new_n978), .B2(new_n956), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n963), .B(new_n969), .C1(new_n928), .C2(new_n953), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n896), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n976), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n958), .A2(new_n964), .A3(KEYINPUT105), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(KEYINPUT43), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n964), .A2(new_n965), .A3(new_n971), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n985), .A2(KEYINPUT44), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n984), .A2(KEYINPUT106), .A3(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT106), .B1(new_n984), .B2(new_n986), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n975), .B1(new_n987), .B2(new_n988), .ZN(G397));
  NAND2_X1  g564(.A1(new_n498), .A2(new_n506), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT107), .B(G1384), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n477), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n484), .A2(G137), .B1(new_n463), .B2(G101), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(G40), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1996), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n821), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n786), .B(G2067), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n817), .A2(G1996), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n734), .A2(new_n736), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n734), .A2(new_n736), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n608), .A2(new_n741), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT110), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n608), .A2(new_n741), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT109), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n999), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1384), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n507), .A2(new_n511), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT50), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n990), .A2(new_n1018), .A3(new_n1015), .ZN(new_n1019));
  INV_X1    g594(.A(new_n998), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT118), .ZN(new_n1022));
  INV_X1    g597(.A(G1961), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1017), .A2(new_n1019), .A3(new_n1024), .A4(new_n1020), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n990), .A2(new_n1015), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n998), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(G2078), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1029), .B(new_n1031), .C1(new_n1016), .C2(new_n994), .ZN(new_n1032));
  INV_X1    g607(.A(G160), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n1016), .B2(new_n994), .ZN(new_n1034));
  INV_X1    g609(.A(G40), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1035), .B1(new_n992), .B2(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1030), .B1(new_n1037), .B2(G2078), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1026), .A2(new_n1032), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(G171), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1036), .A2(new_n1031), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n997), .B(KEYINPUT125), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1041), .A2(new_n996), .A3(new_n995), .A4(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1026), .A2(new_n1043), .A3(G301), .A4(new_n1038), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT54), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1045), .A2(KEYINPUT126), .ZN(new_n1046));
  OAI21_X1  g621(.A(G1981), .B1(new_n599), .B2(new_n601), .ZN(new_n1047));
  INV_X1    g622(.A(new_n601), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n578), .A2(G86), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(new_n705), .A4(new_n597), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1027), .A2(new_n998), .ZN(new_n1054));
  INV_X1    g629(.A(G8), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1047), .A2(KEYINPUT49), .A3(new_n1050), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1053), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT111), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT111), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1053), .A2(new_n1056), .A3(new_n1060), .A4(new_n1057), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1056), .B1(new_n1062), .B2(G288), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1059), .A2(new_n1061), .B1(KEYINPUT52), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n998), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(KEYINPUT50), .B2(new_n1016), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(G2090), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1971), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G303), .A2(G8), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1070), .B(KEYINPUT55), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1071), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1021), .A2(G2090), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1073), .B(G8), .C1(new_n1074), .C2(new_n1068), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n711), .A2(G1976), .ZN(new_n1076));
  OR3_X1    g651(.A1(new_n1063), .A2(KEYINPUT52), .A3(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1064), .A2(new_n1072), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1029), .B1(new_n1016), .B2(new_n994), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n803), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1017), .A2(new_n1019), .A3(new_n830), .A4(new_n1020), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(G168), .A3(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(G8), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1083), .B1(new_n1082), .B2(G8), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1055), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(G286), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1078), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1045), .A2(KEYINPUT126), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1026), .A2(new_n1043), .A3(new_n1038), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1094), .B(KEYINPUT54), .C1(G171), .C2(new_n1039), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1046), .A2(new_n1091), .A3(new_n1092), .A4(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1034), .A2(new_n1036), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT116), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  OAI22_X1  g675(.A1(new_n537), .A2(new_n583), .B1(KEYINPUT76), .B2(KEYINPUT9), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n581), .A2(G53), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(new_n584), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT57), .B1(new_n1103), .B2(KEYINPUT115), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(G299), .ZN(new_n1105));
  INV_X1    g680(.A(G1956), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1066), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1034), .A2(new_n1036), .A3(KEYINPUT116), .A4(new_n1097), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1100), .A2(new_n1105), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT117), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1100), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1105), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT121), .B(KEYINPUT61), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1109), .A2(KEYINPUT122), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1116), .A2(new_n1113), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1109), .A2(KEYINPUT122), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1114), .A2(new_n1115), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1022), .A2(new_n772), .A3(new_n1025), .ZN(new_n1122));
  INV_X1    g697(.A(G2067), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1054), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n625), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1122), .A2(KEYINPUT123), .A3(KEYINPUT60), .A4(new_n1124), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1130), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1127), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT120), .B(G1996), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT58), .B(G1341), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1037), .A2(new_n1136), .B1(new_n1054), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n567), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT59), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1121), .A2(new_n1135), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1125), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1113), .B1(new_n1142), .B2(new_n625), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1110), .A2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT119), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1096), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT114), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT113), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1089), .A2(new_n1148), .A3(G168), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1148), .B1(new_n1089), .B2(G168), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1147), .B1(new_n1152), .B2(new_n1078), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1064), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1089), .A2(G168), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT113), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1149), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1154), .A2(new_n1157), .A3(KEYINPUT114), .A4(new_n1072), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1153), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(G8), .B1(new_n1074), .B2(new_n1068), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1159), .B1(new_n1161), .B2(new_n1071), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1154), .A2(new_n1157), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1087), .A2(new_n1086), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1165), .A2(new_n1090), .A3(new_n1084), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1078), .B1(new_n1166), .B2(KEYINPUT62), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1040), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1167), .B(new_n1168), .C1(KEYINPUT62), .C2(new_n1166), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1170), .A2(new_n1062), .A3(new_n711), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(new_n1050), .ZN(new_n1172));
  XOR2_X1   g747(.A(new_n1056), .B(KEYINPUT112), .Z(new_n1173));
  AND2_X1   g748(.A1(new_n1064), .A2(new_n1077), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1075), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1172), .A2(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1164), .A2(new_n1169), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1014), .B1(new_n1146), .B2(new_n1177), .ZN(new_n1178));
  OAI22_X1  g753(.A1(new_n1004), .A2(new_n1006), .B1(G2067), .B2(new_n879), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1179), .A2(new_n999), .ZN(new_n1180));
  NOR3_X1   g755(.A1(new_n995), .A2(G1996), .A3(new_n998), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n1181), .A2(KEYINPUT46), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1002), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n999), .B1(new_n1183), .B2(new_n817), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1181), .A2(KEYINPUT46), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1182), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT47), .Z(new_n1187));
  NAND2_X1  g762(.A1(new_n1008), .A2(new_n999), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1012), .A2(new_n999), .ZN(new_n1189));
  XOR2_X1   g764(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1190));
  XNOR2_X1  g765(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  AOI211_X1 g766(.A(new_n1180), .B(new_n1187), .C1(new_n1188), .C2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1178), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g768(.A(new_n687), .B1(new_n667), .B2(new_n668), .ZN(new_n1195));
  AOI21_X1  g769(.A(new_n1195), .B1(new_n898), .B2(new_n900), .ZN(new_n1196));
  INV_X1    g770(.A(G229), .ZN(new_n1197));
  NAND4_X1  g771(.A1(new_n1196), .A2(new_n973), .A3(G319), .A4(new_n1197), .ZN(G225));
  INV_X1    g772(.A(G225), .ZN(G308));
endmodule


