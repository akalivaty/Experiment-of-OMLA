
module locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, 
        G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450;

  NOR2_X2 U258 ( .A1(n391), .A2(n390), .ZN(n392) );
  XOR2_X1 U259 ( .A(KEYINPUT41), .B(n442), .Z(n406) );
  NOR2_X1 U260 ( .A1(n419), .A2(n418), .ZN(n437) );
  XOR2_X1 U261 ( .A(n264), .B(n263), .Z(n412) );
  XOR2_X1 U262 ( .A(n293), .B(n292), .Z(n423) );
  XOR2_X1 U263 ( .A(G218GAT), .B(G106GAT), .Z(n226) );
  NOR2_X1 U264 ( .A1(n448), .A2(n445), .ZN(n387) );
  XNOR2_X1 U265 ( .A(n318), .B(n226), .ZN(n260) );
  XNOR2_X1 U266 ( .A(n261), .B(n260), .ZN(n262) );
  XOR2_X1 U267 ( .A(n420), .B(KEYINPUT28), .Z(n395) );
  XOR2_X1 U268 ( .A(G50GAT), .B(G36GAT), .Z(n228) );
  NAND2_X1 U269 ( .A1(G229GAT), .A2(G233GAT), .ZN(n227) );
  XNOR2_X1 U270 ( .A(n228), .B(n227), .ZN(n240) );
  XOR2_X1 U271 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n230) );
  XNOR2_X1 U272 ( .A(G169GAT), .B(G8GAT), .ZN(n229) );
  XNOR2_X1 U273 ( .A(n230), .B(n229), .ZN(n234) );
  XOR2_X1 U274 ( .A(G113GAT), .B(G197GAT), .Z(n232) );
  XNOR2_X1 U275 ( .A(G29GAT), .B(G141GAT), .ZN(n231) );
  XNOR2_X1 U276 ( .A(n232), .B(n231), .ZN(n233) );
  XOR2_X1 U277 ( .A(n234), .B(n233), .Z(n238) );
  XNOR2_X1 U278 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n235) );
  XNOR2_X1 U279 ( .A(n235), .B(KEYINPUT7), .ZN(n257) );
  XNOR2_X1 U280 ( .A(G22GAT), .B(G15GAT), .ZN(n236) );
  XNOR2_X1 U281 ( .A(n236), .B(G1GAT), .ZN(n272) );
  XNOR2_X1 U282 ( .A(n257), .B(n272), .ZN(n237) );
  XNOR2_X1 U283 ( .A(n238), .B(n237), .ZN(n239) );
  XNOR2_X1 U284 ( .A(n240), .B(n239), .ZN(n438) );
  INV_X1 U285 ( .A(n438), .ZN(n424) );
  XNOR2_X1 U286 ( .A(G71GAT), .B(G57GAT), .ZN(n241) );
  XNOR2_X1 U287 ( .A(n241), .B(KEYINPUT13), .ZN(n271) );
  XOR2_X1 U288 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n243) );
  NAND2_X1 U289 ( .A1(G230GAT), .A2(G233GAT), .ZN(n242) );
  XNOR2_X1 U290 ( .A(n243), .B(n242), .ZN(n244) );
  XOR2_X1 U291 ( .A(n244), .B(KEYINPUT32), .Z(n248) );
  XNOR2_X1 U292 ( .A(G106GAT), .B(G78GAT), .ZN(n245) );
  XNOR2_X1 U293 ( .A(n245), .B(G148GAT), .ZN(n296) );
  XNOR2_X1 U294 ( .A(G99GAT), .B(G85GAT), .ZN(n246) );
  XNOR2_X1 U295 ( .A(n246), .B(G92GAT), .ZN(n256) );
  XNOR2_X1 U296 ( .A(n296), .B(n256), .ZN(n247) );
  XNOR2_X1 U297 ( .A(n248), .B(n247), .ZN(n249) );
  XOR2_X1 U298 ( .A(G176GAT), .B(G64GAT), .Z(n324) );
  XOR2_X1 U299 ( .A(n249), .B(n324), .Z(n251) );
  XNOR2_X1 U300 ( .A(G120GAT), .B(G204GAT), .ZN(n250) );
  XNOR2_X1 U301 ( .A(n251), .B(n250), .ZN(n252) );
  XOR2_X1 U302 ( .A(n271), .B(n252), .Z(n442) );
  NAND2_X1 U303 ( .A1(n424), .A2(n442), .ZN(n358) );
  XOR2_X1 U304 ( .A(G50GAT), .B(G162GAT), .Z(n306) );
  XOR2_X1 U305 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n254) );
  NAND2_X1 U306 ( .A1(G232GAT), .A2(G233GAT), .ZN(n253) );
  XNOR2_X1 U307 ( .A(n254), .B(n253), .ZN(n255) );
  XOR2_X1 U308 ( .A(n255), .B(KEYINPUT9), .Z(n259) );
  XNOR2_X1 U309 ( .A(n257), .B(n256), .ZN(n258) );
  XNOR2_X1 U310 ( .A(n259), .B(n258), .ZN(n261) );
  XOR2_X1 U311 ( .A(G29GAT), .B(G134GAT), .Z(n318) );
  XNOR2_X1 U312 ( .A(n306), .B(n262), .ZN(n264) );
  XNOR2_X1 U313 ( .A(G36GAT), .B(G190GAT), .ZN(n329) );
  INV_X1 U314 ( .A(n329), .ZN(n263) );
  INV_X1 U315 ( .A(n412), .ZN(n433) );
  XOR2_X1 U316 ( .A(G8GAT), .B(G183GAT), .Z(n327) );
  XOR2_X1 U317 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n266) );
  XNOR2_X1 U318 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n265) );
  XNOR2_X1 U319 ( .A(n266), .B(n265), .ZN(n270) );
  XOR2_X1 U320 ( .A(G78GAT), .B(G155GAT), .Z(n268) );
  XNOR2_X1 U321 ( .A(G127GAT), .B(G211GAT), .ZN(n267) );
  XNOR2_X1 U322 ( .A(n268), .B(n267), .ZN(n269) );
  XOR2_X1 U323 ( .A(n270), .B(n269), .Z(n274) );
  XNOR2_X1 U324 ( .A(n272), .B(n271), .ZN(n273) );
  XNOR2_X1 U325 ( .A(n274), .B(n273), .ZN(n275) );
  XOR2_X1 U326 ( .A(n327), .B(n275), .Z(n277) );
  NAND2_X1 U327 ( .A1(G231GAT), .A2(G233GAT), .ZN(n276) );
  XOR2_X1 U328 ( .A(n277), .B(n276), .Z(n445) );
  NOR2_X1 U329 ( .A1(n433), .A2(n445), .ZN(n278) );
  XNOR2_X1 U330 ( .A(n278), .B(KEYINPUT16), .ZN(n347) );
  XOR2_X1 U331 ( .A(G120GAT), .B(G127GAT), .Z(n280) );
  XNOR2_X1 U332 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n279) );
  XNOR2_X1 U333 ( .A(n280), .B(n279), .ZN(n315) );
  XOR2_X1 U334 ( .A(n315), .B(G15GAT), .Z(n282) );
  NAND2_X1 U335 ( .A1(G227GAT), .A2(G233GAT), .ZN(n281) );
  XNOR2_X1 U336 ( .A(n282), .B(n281), .ZN(n286) );
  XOR2_X1 U337 ( .A(G176GAT), .B(G183GAT), .Z(n284) );
  XNOR2_X1 U338 ( .A(G71GAT), .B(KEYINPUT20), .ZN(n283) );
  XNOR2_X1 U339 ( .A(n284), .B(n283), .ZN(n285) );
  XOR2_X1 U340 ( .A(n286), .B(n285), .Z(n293) );
  XOR2_X1 U341 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n288) );
  XNOR2_X1 U342 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n287) );
  XNOR2_X1 U343 ( .A(n288), .B(n287), .ZN(n334) );
  XOR2_X1 U344 ( .A(G134GAT), .B(G190GAT), .Z(n290) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(G99GAT), .ZN(n289) );
  XNOR2_X1 U346 ( .A(n290), .B(n289), .ZN(n291) );
  XNOR2_X1 U347 ( .A(n334), .B(n291), .ZN(n292) );
  INV_X1 U348 ( .A(n423), .ZN(n336) );
  XOR2_X1 U349 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n295) );
  XNOR2_X1 U350 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n297) );
  XOR2_X1 U352 ( .A(n297), .B(n296), .Z(n304) );
  XOR2_X1 U353 ( .A(G211GAT), .B(G218GAT), .Z(n299) );
  XNOR2_X1 U354 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U356 ( .A(G197GAT), .B(n300), .Z(n330) );
  XOR2_X1 U357 ( .A(G155GAT), .B(KEYINPUT3), .Z(n302) );
  XNOR2_X1 U358 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n301) );
  XNOR2_X1 U359 ( .A(n302), .B(n301), .ZN(n313) );
  XNOR2_X1 U360 ( .A(n330), .B(n313), .ZN(n303) );
  XNOR2_X1 U361 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U362 ( .A(n306), .B(n305), .Z(n308) );
  NAND2_X1 U363 ( .A1(G228GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n420) );
  XOR2_X1 U365 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n310) );
  XNOR2_X1 U366 ( .A(G148GAT), .B(KEYINPUT6), .ZN(n309) );
  XNOR2_X1 U367 ( .A(n310), .B(n309), .ZN(n323) );
  XOR2_X1 U368 ( .A(KEYINPUT1), .B(G57GAT), .Z(n312) );
  NAND2_X1 U369 ( .A1(G225GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U370 ( .A(n312), .B(n311), .ZN(n314) );
  XOR2_X1 U371 ( .A(n314), .B(n313), .Z(n317) );
  XNOR2_X1 U372 ( .A(G1GAT), .B(n315), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n319) );
  XOR2_X1 U374 ( .A(n319), .B(n318), .Z(n321) );
  XNOR2_X1 U375 ( .A(G162GAT), .B(G85GAT), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U377 ( .A(n323), .B(n322), .ZN(n343) );
  INV_X1 U378 ( .A(n343), .ZN(n419) );
  XOR2_X1 U379 ( .A(n324), .B(G92GAT), .Z(n326) );
  NAND2_X1 U380 ( .A1(G226GAT), .A2(G233GAT), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n328) );
  XOR2_X1 U382 ( .A(n328), .B(n327), .Z(n332) );
  XOR2_X1 U383 ( .A(n330), .B(n329), .Z(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U385 ( .A(n334), .B(n333), .ZN(n414) );
  XNOR2_X1 U386 ( .A(n414), .B(KEYINPUT27), .ZN(n338) );
  NAND2_X1 U387 ( .A1(n419), .A2(n338), .ZN(n393) );
  NOR2_X1 U388 ( .A1(n395), .A2(n393), .ZN(n335) );
  NAND2_X1 U389 ( .A1(n336), .A2(n335), .ZN(n346) );
  NOR2_X1 U390 ( .A1(n423), .A2(n420), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n337), .B(KEYINPUT26), .ZN(n436) );
  NAND2_X1 U392 ( .A1(n436), .A2(n338), .ZN(n342) );
  NAND2_X1 U393 ( .A1(n423), .A2(n414), .ZN(n339) );
  NAND2_X1 U394 ( .A1(n420), .A2(n339), .ZN(n340) );
  XOR2_X1 U395 ( .A(KEYINPUT25), .B(n340), .Z(n341) );
  NAND2_X1 U396 ( .A1(n342), .A2(n341), .ZN(n344) );
  NAND2_X1 U397 ( .A1(n344), .A2(n343), .ZN(n345) );
  NAND2_X1 U398 ( .A1(n346), .A2(n345), .ZN(n355) );
  NAND2_X1 U399 ( .A1(n347), .A2(n355), .ZN(n367) );
  NOR2_X1 U400 ( .A1(n358), .A2(n367), .ZN(n353) );
  NAND2_X1 U401 ( .A1(n353), .A2(n419), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n348), .B(KEYINPUT34), .ZN(n349) );
  XNOR2_X1 U403 ( .A(G1GAT), .B(n349), .ZN(G1324GAT) );
  NAND2_X1 U404 ( .A1(n414), .A2(n353), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n350), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U406 ( .A(G15GAT), .B(KEYINPUT35), .Z(n352) );
  NAND2_X1 U407 ( .A1(n353), .A2(n423), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(G1326GAT) );
  NAND2_X1 U409 ( .A1(n353), .A2(n395), .ZN(n354) );
  XNOR2_X1 U410 ( .A(n354), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U411 ( .A(G29GAT), .B(KEYINPUT39), .Z(n361) );
  XOR2_X1 U412 ( .A(KEYINPUT36), .B(n433), .Z(n448) );
  NAND2_X1 U413 ( .A1(n445), .A2(n355), .ZN(n356) );
  NOR2_X1 U414 ( .A1(n448), .A2(n356), .ZN(n357) );
  XNOR2_X1 U415 ( .A(KEYINPUT37), .B(n357), .ZN(n376) );
  NOR2_X1 U416 ( .A1(n376), .A2(n358), .ZN(n359) );
  XNOR2_X1 U417 ( .A(KEYINPUT38), .B(n359), .ZN(n365) );
  NAND2_X1 U418 ( .A1(n419), .A2(n365), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n361), .B(n360), .ZN(G1328GAT) );
  NAND2_X1 U420 ( .A1(n365), .A2(n414), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n362), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U422 ( .A1(n365), .A2(n423), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n363), .B(KEYINPUT40), .ZN(n364) );
  XNOR2_X1 U424 ( .A(G43GAT), .B(n364), .ZN(G1330GAT) );
  NAND2_X1 U425 ( .A1(n365), .A2(n395), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n366), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U427 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n369) );
  INV_X1 U428 ( .A(n406), .ZN(n426) );
  NAND2_X1 U429 ( .A1(n438), .A2(n426), .ZN(n375) );
  NOR2_X1 U430 ( .A1(n375), .A2(n367), .ZN(n372) );
  NAND2_X1 U431 ( .A1(n419), .A2(n372), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n369), .B(n368), .ZN(G1332GAT) );
  NAND2_X1 U433 ( .A1(n414), .A2(n372), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n370), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U435 ( .A1(n423), .A2(n372), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n371), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U437 ( .A(G78GAT), .B(KEYINPUT43), .Z(n374) );
  NAND2_X1 U438 ( .A1(n372), .A2(n395), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(G1335GAT) );
  NOR2_X1 U440 ( .A1(n376), .A2(n375), .ZN(n380) );
  NAND2_X1 U441 ( .A1(n419), .A2(n380), .ZN(n377) );
  XNOR2_X1 U442 ( .A(G85GAT), .B(n377), .ZN(G1336GAT) );
  NAND2_X1 U443 ( .A1(n414), .A2(n380), .ZN(n378) );
  XNOR2_X1 U444 ( .A(n378), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U445 ( .A1(n423), .A2(n380), .ZN(n379) );
  XNOR2_X1 U446 ( .A(n379), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U447 ( .A1(n380), .A2(n395), .ZN(n381) );
  XNOR2_X1 U448 ( .A(n381), .B(KEYINPUT44), .ZN(n382) );
  XNOR2_X1 U449 ( .A(G106GAT), .B(n382), .ZN(G1339GAT) );
  INV_X1 U450 ( .A(n445), .ZN(n430) );
  NOR2_X1 U451 ( .A1(n406), .A2(n438), .ZN(n383) );
  XNOR2_X1 U452 ( .A(n383), .B(KEYINPUT46), .ZN(n384) );
  NOR2_X1 U453 ( .A1(n430), .A2(n384), .ZN(n385) );
  NAND2_X1 U454 ( .A1(n385), .A2(n412), .ZN(n386) );
  XNOR2_X1 U455 ( .A(KEYINPUT47), .B(n386), .ZN(n391) );
  XNOR2_X1 U456 ( .A(KEYINPUT45), .B(n387), .ZN(n388) );
  NAND2_X1 U457 ( .A1(n388), .A2(n442), .ZN(n389) );
  NOR2_X1 U458 ( .A1(n424), .A2(n389), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n392), .B(KEYINPUT48), .ZN(n416) );
  NOR2_X1 U460 ( .A1(n416), .A2(n393), .ZN(n404) );
  NAND2_X1 U461 ( .A1(n404), .A2(n423), .ZN(n394) );
  NOR2_X1 U462 ( .A1(n395), .A2(n394), .ZN(n401) );
  NAND2_X1 U463 ( .A1(n424), .A2(n401), .ZN(n396) );
  XNOR2_X1 U464 ( .A(G113GAT), .B(n396), .ZN(G1340GAT) );
  XOR2_X1 U465 ( .A(G120GAT), .B(KEYINPUT49), .Z(n398) );
  NAND2_X1 U466 ( .A1(n401), .A2(n426), .ZN(n397) );
  XNOR2_X1 U467 ( .A(n398), .B(n397), .ZN(G1341GAT) );
  NAND2_X1 U468 ( .A1(n401), .A2(n430), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n399), .B(KEYINPUT50), .ZN(n400) );
  XNOR2_X1 U470 ( .A(G127GAT), .B(n400), .ZN(G1342GAT) );
  XOR2_X1 U471 ( .A(G134GAT), .B(KEYINPUT51), .Z(n403) );
  NAND2_X1 U472 ( .A1(n401), .A2(n433), .ZN(n402) );
  XNOR2_X1 U473 ( .A(n403), .B(n402), .ZN(G1343GAT) );
  NAND2_X1 U474 ( .A1(n404), .A2(n436), .ZN(n411) );
  NOR2_X1 U475 ( .A1(n438), .A2(n411), .ZN(n405) );
  XOR2_X1 U476 ( .A(G141GAT), .B(n405), .Z(G1344GAT) );
  NOR2_X1 U477 ( .A1(n406), .A2(n411), .ZN(n408) );
  XNOR2_X1 U478 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n407) );
  XNOR2_X1 U479 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U480 ( .A(G148GAT), .B(n409), .ZN(G1345GAT) );
  NOR2_X1 U481 ( .A1(n445), .A2(n411), .ZN(n410) );
  XOR2_X1 U482 ( .A(G155GAT), .B(n410), .Z(G1346GAT) );
  NOR2_X1 U483 ( .A1(n412), .A2(n411), .ZN(n413) );
  XOR2_X1 U484 ( .A(G162GAT), .B(n413), .Z(G1347GAT) );
  INV_X1 U485 ( .A(n414), .ZN(n415) );
  NOR2_X1 U486 ( .A1(n416), .A2(n415), .ZN(n417) );
  XOR2_X1 U487 ( .A(KEYINPUT54), .B(n417), .Z(n418) );
  NAND2_X1 U488 ( .A1(n420), .A2(n437), .ZN(n421) );
  XNOR2_X1 U489 ( .A(KEYINPUT55), .B(n421), .ZN(n422) );
  AND2_X2 U490 ( .A1(n423), .A2(n422), .ZN(n432) );
  NAND2_X1 U491 ( .A1(n432), .A2(n424), .ZN(n425) );
  XNOR2_X1 U492 ( .A(n425), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U493 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n428) );
  NAND2_X1 U494 ( .A1(n432), .A2(n426), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U496 ( .A(G176GAT), .B(n429), .ZN(G1349GAT) );
  NAND2_X1 U497 ( .A1(n432), .A2(n430), .ZN(n431) );
  XNOR2_X1 U498 ( .A(n431), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U499 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n435) );
  NAND2_X1 U500 ( .A1(n433), .A2(n432), .ZN(n434) );
  XNOR2_X1 U501 ( .A(n435), .B(n434), .ZN(G1351GAT) );
  NAND2_X1 U502 ( .A1(n437), .A2(n436), .ZN(n447) );
  NOR2_X1 U503 ( .A1(n438), .A2(n447), .ZN(n440) );
  XNOR2_X1 U504 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n439) );
  XNOR2_X1 U505 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U506 ( .A(G197GAT), .B(n441), .ZN(G1352GAT) );
  NOR2_X1 U507 ( .A1(n442), .A2(n447), .ZN(n444) );
  XNOR2_X1 U508 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n443) );
  XNOR2_X1 U509 ( .A(n444), .B(n443), .ZN(G1353GAT) );
  NOR2_X1 U510 ( .A1(n445), .A2(n447), .ZN(n446) );
  XOR2_X1 U511 ( .A(G211GAT), .B(n446), .Z(G1354GAT) );
  NOR2_X1 U512 ( .A1(n448), .A2(n447), .ZN(n449) );
  XOR2_X1 U513 ( .A(KEYINPUT62), .B(n449), .Z(n450) );
  XNOR2_X1 U514 ( .A(G218GAT), .B(n450), .ZN(G1355GAT) );
endmodule

