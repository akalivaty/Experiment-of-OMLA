

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580;

  INV_X1 U319 ( .A(n293), .ZN(n290) );
  AND2_X1 U320 ( .A1(G232GAT), .A2(G233GAT), .ZN(n287) );
  OR2_X1 U321 ( .A1(n377), .A2(n376), .ZN(n378) );
  XNOR2_X1 U322 ( .A(KEYINPUT70), .B(G92GAT), .ZN(n293) );
  XNOR2_X1 U323 ( .A(n289), .B(n409), .ZN(n297) );
  XNOR2_X1 U324 ( .A(n297), .B(n356), .ZN(n298) );
  XNOR2_X1 U325 ( .A(n349), .B(n287), .ZN(n350) );
  XNOR2_X1 U326 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U327 ( .A(n351), .B(n350), .ZN(n353) );
  XNOR2_X1 U328 ( .A(n305), .B(n304), .ZN(n383) );
  NOR2_X1 U329 ( .A1(n526), .A2(n449), .ZN(n557) );
  XNOR2_X1 U330 ( .A(n530), .B(KEYINPUT117), .ZN(n539) );
  XOR2_X1 U331 ( .A(KEYINPUT28), .B(n468), .Z(n528) );
  XNOR2_X1 U332 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U333 ( .A(n453), .B(n452), .ZN(G1349GAT) );
  INV_X1 U334 ( .A(KEYINPUT41), .ZN(n306) );
  XNOR2_X1 U335 ( .A(G176GAT), .B(G64GAT), .ZN(n288) );
  XNOR2_X1 U336 ( .A(n288), .B(G204GAT), .ZN(n396) );
  XOR2_X1 U337 ( .A(G71GAT), .B(KEYINPUT13), .Z(n336) );
  XOR2_X1 U338 ( .A(n396), .B(n336), .Z(n289) );
  XOR2_X1 U339 ( .A(G120GAT), .B(G57GAT), .Z(n409) );
  XNOR2_X1 U340 ( .A(G99GAT), .B(G106GAT), .ZN(n291) );
  NAND2_X1 U341 ( .A1(n290), .A2(n291), .ZN(n295) );
  INV_X1 U342 ( .A(n291), .ZN(n292) );
  NAND2_X1 U343 ( .A1(n293), .A2(n292), .ZN(n294) );
  NAND2_X1 U344 ( .A1(n295), .A2(n294), .ZN(n296) );
  XOR2_X1 U345 ( .A(G85GAT), .B(n296), .Z(n356) );
  XOR2_X1 U346 ( .A(G148GAT), .B(G78GAT), .Z(n431) );
  XOR2_X1 U347 ( .A(n298), .B(n431), .Z(n305) );
  XOR2_X1 U348 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n300) );
  NAND2_X1 U349 ( .A1(G230GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U351 ( .A(KEYINPUT33), .B(n301), .ZN(n303) );
  XNOR2_X1 U352 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n302) );
  XNOR2_X1 U353 ( .A(n306), .B(n383), .ZN(n374) );
  XOR2_X1 U354 ( .A(n374), .B(KEYINPUT106), .Z(n532) );
  XOR2_X1 U355 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n308) );
  XNOR2_X1 U356 ( .A(G176GAT), .B(KEYINPUT79), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n326) );
  XOR2_X1 U358 ( .A(G99GAT), .B(G190GAT), .Z(n310) );
  XNOR2_X1 U359 ( .A(G43GAT), .B(G134GAT), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U361 ( .A(G71GAT), .B(G120GAT), .Z(n312) );
  XNOR2_X1 U362 ( .A(G169GAT), .B(G15GAT), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U364 ( .A(n314), .B(n313), .Z(n324) );
  XOR2_X1 U365 ( .A(KEYINPUT17), .B(G183GAT), .Z(n316) );
  XNOR2_X1 U366 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U368 ( .A(KEYINPUT80), .B(n317), .Z(n394) );
  XOR2_X1 U369 ( .A(G127GAT), .B(KEYINPUT78), .Z(n319) );
  XNOR2_X1 U370 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n412) );
  XOR2_X1 U372 ( .A(n412), .B(KEYINPUT20), .Z(n321) );
  NAND2_X1 U373 ( .A1(G227GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n394), .B(n322), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U377 ( .A(n326), .B(n325), .ZN(n526) );
  XOR2_X1 U378 ( .A(KEYINPUT114), .B(KEYINPUT48), .Z(n390) );
  XOR2_X1 U379 ( .A(KEYINPUT47), .B(KEYINPUT112), .Z(n379) );
  XOR2_X1 U380 ( .A(G211GAT), .B(KEYINPUT75), .Z(n328) );
  XNOR2_X1 U381 ( .A(G78GAT), .B(G64GAT), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U383 ( .A(KEYINPUT76), .B(KEYINPUT12), .Z(n330) );
  XNOR2_X1 U384 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U386 ( .A(n332), .B(n331), .ZN(n344) );
  XOR2_X1 U387 ( .A(G57GAT), .B(G155GAT), .Z(n334) );
  XNOR2_X1 U388 ( .A(G8GAT), .B(G127GAT), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U390 ( .A(n336), .B(n335), .Z(n338) );
  NAND2_X1 U391 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U393 ( .A(n339), .B(KEYINPUT77), .Z(n342) );
  XNOR2_X1 U394 ( .A(G1GAT), .B(G22GAT), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n340), .B(G15GAT), .ZN(n365) );
  XNOR2_X1 U396 ( .A(n365), .B(G183GAT), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n535) );
  XOR2_X1 U399 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n346) );
  XOR2_X1 U400 ( .A(G29GAT), .B(G134GAT), .Z(n413) );
  XOR2_X1 U401 ( .A(G50GAT), .B(G162GAT), .Z(n440) );
  XNOR2_X1 U402 ( .A(n413), .B(n440), .ZN(n345) );
  XNOR2_X1 U403 ( .A(n346), .B(n345), .ZN(n351) );
  XOR2_X1 U404 ( .A(KEYINPUT73), .B(KEYINPUT9), .Z(n348) );
  XNOR2_X1 U405 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U407 ( .A(G36GAT), .B(G190GAT), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n352), .B(G218GAT), .ZN(n400) );
  XOR2_X1 U409 ( .A(n353), .B(n400), .Z(n358) );
  XOR2_X1 U410 ( .A(G43GAT), .B(KEYINPUT7), .Z(n355) );
  XNOR2_X1 U411 ( .A(KEYINPUT66), .B(KEYINPUT8), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n369) );
  XNOR2_X1 U413 ( .A(n369), .B(n356), .ZN(n357) );
  XNOR2_X1 U414 ( .A(n358), .B(n357), .ZN(n553) );
  NAND2_X1 U415 ( .A1(n535), .A2(n553), .ZN(n377) );
  XOR2_X1 U416 ( .A(G141GAT), .B(G36GAT), .Z(n360) );
  XNOR2_X1 U417 ( .A(G50GAT), .B(G29GAT), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U419 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n362) );
  XNOR2_X1 U420 ( .A(G113GAT), .B(G197GAT), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n373) );
  XOR2_X1 U423 ( .A(G169GAT), .B(G8GAT), .Z(n395) );
  XOR2_X1 U424 ( .A(n365), .B(n395), .Z(n367) );
  NAND2_X1 U425 ( .A1(G229GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U427 ( .A(n368), .B(KEYINPUT65), .Z(n371) );
  XNOR2_X1 U428 ( .A(n369), .B(KEYINPUT67), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n373), .B(n372), .ZN(n522) );
  NOR2_X1 U431 ( .A1(n522), .A2(n374), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n375), .B(KEYINPUT46), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n388) );
  INV_X1 U434 ( .A(KEYINPUT74), .ZN(n380) );
  XNOR2_X1 U435 ( .A(n380), .B(n553), .ZN(n472) );
  XOR2_X1 U436 ( .A(KEYINPUT36), .B(KEYINPUT102), .Z(n381) );
  XNOR2_X1 U437 ( .A(n472), .B(n381), .ZN(n578) );
  NOR2_X1 U438 ( .A1(n535), .A2(n578), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n382), .B(KEYINPUT45), .ZN(n384) );
  INV_X1 U440 ( .A(n383), .ZN(n568) );
  NAND2_X1 U441 ( .A1(n384), .A2(n383), .ZN(n385) );
  XNOR2_X1 U442 ( .A(KEYINPUT113), .B(n385), .ZN(n386) );
  NAND2_X1 U443 ( .A1(n386), .A2(n522), .ZN(n387) );
  NAND2_X1 U444 ( .A1(n388), .A2(n387), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n523) );
  XOR2_X1 U446 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n392) );
  XNOR2_X1 U447 ( .A(G197GAT), .B(G211GAT), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U449 ( .A(KEYINPUT86), .B(n393), .ZN(n446) );
  XOR2_X1 U450 ( .A(n394), .B(n446), .Z(n404) );
  XOR2_X1 U451 ( .A(n396), .B(n395), .Z(n398) );
  NAND2_X1 U452 ( .A1(G226GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U453 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U454 ( .A(n399), .B(KEYINPUT75), .Z(n402) );
  XNOR2_X1 U455 ( .A(G92GAT), .B(n400), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U457 ( .A(n404), .B(n403), .ZN(n516) );
  NOR2_X1 U458 ( .A1(n523), .A2(n516), .ZN(n405) );
  XNOR2_X1 U459 ( .A(KEYINPUT54), .B(n405), .ZN(n426) );
  XOR2_X1 U460 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n407) );
  XNOR2_X1 U461 ( .A(G162GAT), .B(G85GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U463 ( .A(n408), .B(KEYINPUT91), .Z(n411) );
  XNOR2_X1 U464 ( .A(G1GAT), .B(n409), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n417) );
  XOR2_X1 U466 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U467 ( .A1(G225GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U469 ( .A(n417), .B(n416), .Z(n425) );
  XOR2_X1 U470 ( .A(KEYINPUT87), .B(KEYINPUT2), .Z(n419) );
  XNOR2_X1 U471 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n418) );
  XNOR2_X1 U472 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U473 ( .A(G141GAT), .B(n420), .Z(n441) );
  XOR2_X1 U474 ( .A(G148GAT), .B(KEYINPUT6), .Z(n422) );
  XNOR2_X1 U475 ( .A(KEYINPUT5), .B(KEYINPUT92), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n441), .B(n423), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n464) );
  XNOR2_X1 U479 ( .A(KEYINPUT93), .B(n464), .ZN(n513) );
  NAND2_X1 U480 ( .A1(n426), .A2(n513), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n427), .B(KEYINPUT64), .ZN(n561) );
  XOR2_X1 U482 ( .A(KEYINPUT24), .B(KEYINPUT90), .Z(n429) );
  XNOR2_X1 U483 ( .A(G106GAT), .B(G218GAT), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U485 ( .A(n430), .B(G204GAT), .Z(n433) );
  XNOR2_X1 U486 ( .A(G22GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n445) );
  XOR2_X1 U488 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n435) );
  XNOR2_X1 U489 ( .A(KEYINPUT83), .B(KEYINPUT89), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U491 ( .A(KEYINPUT84), .B(KEYINPUT23), .Z(n437) );
  NAND2_X1 U492 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U494 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n447), .B(n446), .ZN(n468) );
  NOR2_X1 U499 ( .A1(n561), .A2(n468), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n448), .B(KEYINPUT55), .ZN(n449) );
  NAND2_X1 U501 ( .A1(n532), .A2(n557), .ZN(n453) );
  XOR2_X1 U502 ( .A(G176GAT), .B(KEYINPUT56), .Z(n451) );
  XNOR2_X1 U503 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n450) );
  NOR2_X1 U504 ( .A1(n522), .A2(n568), .ZN(n488) );
  XNOR2_X1 U505 ( .A(KEYINPUT25), .B(KEYINPUT98), .ZN(n454) );
  XNOR2_X1 U506 ( .A(n454), .B(KEYINPUT97), .ZN(n457) );
  NOR2_X1 U507 ( .A1(n516), .A2(n526), .ZN(n455) );
  NOR2_X1 U508 ( .A1(n468), .A2(n455), .ZN(n456) );
  XNOR2_X1 U509 ( .A(n457), .B(n456), .ZN(n462) );
  NAND2_X1 U510 ( .A1(n468), .A2(n526), .ZN(n458) );
  XNOR2_X1 U511 ( .A(n458), .B(KEYINPUT96), .ZN(n459) );
  XNOR2_X1 U512 ( .A(KEYINPUT26), .B(n459), .ZN(n560) );
  XNOR2_X1 U513 ( .A(n516), .B(KEYINPUT94), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n460), .B(KEYINPUT27), .ZN(n466) );
  NOR2_X1 U515 ( .A1(n560), .A2(n466), .ZN(n461) );
  NOR2_X1 U516 ( .A1(n462), .A2(n461), .ZN(n463) );
  NOR2_X1 U517 ( .A1(n464), .A2(n463), .ZN(n465) );
  XOR2_X1 U518 ( .A(KEYINPUT99), .B(n465), .Z(n471) );
  NOR2_X1 U519 ( .A1(n513), .A2(n466), .ZN(n467) );
  XNOR2_X1 U520 ( .A(n467), .B(KEYINPUT95), .ZN(n524) );
  NAND2_X1 U521 ( .A1(n526), .A2(n528), .ZN(n469) );
  NOR2_X1 U522 ( .A1(n524), .A2(n469), .ZN(n470) );
  NOR2_X1 U523 ( .A1(n471), .A2(n470), .ZN(n484) );
  NOR2_X1 U524 ( .A1(n472), .A2(n535), .ZN(n473) );
  XOR2_X1 U525 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  NOR2_X1 U526 ( .A1(n484), .A2(n474), .ZN(n499) );
  NAND2_X1 U527 ( .A1(n488), .A2(n499), .ZN(n481) );
  NOR2_X1 U528 ( .A1(n513), .A2(n481), .ZN(n475) );
  XOR2_X1 U529 ( .A(KEYINPUT34), .B(n475), .Z(n476) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(n476), .ZN(G1324GAT) );
  NOR2_X1 U531 ( .A1(n516), .A2(n481), .ZN(n477) );
  XOR2_X1 U532 ( .A(G8GAT), .B(n477), .Z(G1325GAT) );
  NOR2_X1 U533 ( .A1(n526), .A2(n481), .ZN(n479) );
  XNOR2_X1 U534 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U535 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U536 ( .A(G15GAT), .B(n480), .ZN(G1326GAT) );
  NOR2_X1 U537 ( .A1(n528), .A2(n481), .ZN(n483) );
  XNOR2_X1 U538 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n483), .B(n482), .ZN(G1327GAT) );
  NOR2_X1 U540 ( .A1(n484), .A2(n578), .ZN(n485) );
  NAND2_X1 U541 ( .A1(n535), .A2(n485), .ZN(n487) );
  XOR2_X1 U542 ( .A(KEYINPUT103), .B(KEYINPUT37), .Z(n486) );
  XNOR2_X1 U543 ( .A(n487), .B(n486), .ZN(n512) );
  NAND2_X1 U544 ( .A1(n488), .A2(n512), .ZN(n489) );
  XNOR2_X1 U545 ( .A(n489), .B(KEYINPUT38), .ZN(n496) );
  NOR2_X1 U546 ( .A1(n496), .A2(n513), .ZN(n491) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  NOR2_X1 U549 ( .A1(n516), .A2(n496), .ZN(n492) );
  XOR2_X1 U550 ( .A(KEYINPUT104), .B(n492), .Z(n493) );
  XNOR2_X1 U551 ( .A(G36GAT), .B(n493), .ZN(G1329GAT) );
  NOR2_X1 U552 ( .A1(n496), .A2(n526), .ZN(n494) );
  XOR2_X1 U553 ( .A(KEYINPUT40), .B(n494), .Z(n495) );
  XNOR2_X1 U554 ( .A(G43GAT), .B(n495), .ZN(G1330GAT) );
  NOR2_X1 U555 ( .A1(n496), .A2(n528), .ZN(n498) );
  XNOR2_X1 U556 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1331GAT) );
  AND2_X1 U558 ( .A1(n522), .A2(n532), .ZN(n511) );
  NAND2_X1 U559 ( .A1(n511), .A2(n499), .ZN(n506) );
  NOR2_X1 U560 ( .A1(n513), .A2(n506), .ZN(n500) );
  XOR2_X1 U561 ( .A(G57GAT), .B(n500), .Z(n501) );
  XNOR2_X1 U562 ( .A(KEYINPUT42), .B(n501), .ZN(G1332GAT) );
  NOR2_X1 U563 ( .A1(n516), .A2(n506), .ZN(n503) );
  XNOR2_X1 U564 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U566 ( .A(G64GAT), .B(n504), .ZN(G1333GAT) );
  NOR2_X1 U567 ( .A1(n526), .A2(n506), .ZN(n505) );
  XOR2_X1 U568 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  NOR2_X1 U569 ( .A1(n506), .A2(n528), .ZN(n510) );
  XOR2_X1 U570 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n508) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT110), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U574 ( .A1(n512), .A2(n511), .ZN(n519) );
  NOR2_X1 U575 ( .A1(n513), .A2(n519), .ZN(n515) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n515), .B(n514), .ZN(G1336GAT) );
  NOR2_X1 U578 ( .A1(n516), .A2(n519), .ZN(n517) );
  XOR2_X1 U579 ( .A(G92GAT), .B(n517), .Z(G1337GAT) );
  NOR2_X1 U580 ( .A1(n526), .A2(n519), .ZN(n518) );
  XOR2_X1 U581 ( .A(G99GAT), .B(n518), .Z(G1338GAT) );
  NOR2_X1 U582 ( .A1(n528), .A2(n519), .ZN(n520) );
  XOR2_X1 U583 ( .A(KEYINPUT44), .B(n520), .Z(n521) );
  XNOR2_X1 U584 ( .A(G106GAT), .B(n521), .ZN(G1339GAT) );
  INV_X1 U585 ( .A(n522), .ZN(n563) );
  NOR2_X1 U586 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n525), .B(KEYINPUT115), .ZN(n543) );
  NOR2_X1 U588 ( .A1(n526), .A2(n543), .ZN(n527) );
  XNOR2_X1 U589 ( .A(n527), .B(KEYINPUT116), .ZN(n529) );
  NAND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U591 ( .A1(n563), .A2(n539), .ZN(n531) );
  XNOR2_X1 U592 ( .A(n531), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U594 ( .A1(n539), .A2(n532), .ZN(n533) );
  XNOR2_X1 U595 ( .A(n534), .B(n533), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n537) );
  INV_X1 U597 ( .A(n535), .ZN(n571) );
  NAND2_X1 U598 ( .A1(n539), .A2(n571), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U600 ( .A(n538), .B(G127GAT), .Z(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U602 ( .A1(n539), .A2(n472), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U604 ( .A(G134GAT), .B(n542), .Z(G1343GAT) );
  NOR2_X1 U605 ( .A1(n543), .A2(n560), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n549), .A2(n563), .ZN(n544) );
  XNOR2_X1 U607 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n548) );
  INV_X1 U611 ( .A(n549), .ZN(n552) );
  NOR2_X1 U612 ( .A1(n374), .A2(n552), .ZN(n547) );
  XOR2_X1 U613 ( .A(n548), .B(n547), .Z(G1345GAT) );
  XOR2_X1 U614 ( .A(G155GAT), .B(KEYINPUT121), .Z(n551) );
  NAND2_X1 U615 ( .A1(n549), .A2(n571), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n551), .B(n550), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n554), .Z(G1347GAT) );
  NAND2_X1 U619 ( .A1(n563), .A2(n557), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U621 ( .A1(n571), .A2(n557), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n472), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT58), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G190GAT), .B(n559), .ZN(G1351GAT) );
  NOR2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(KEYINPUT123), .B(n562), .Z(n576) );
  NAND2_X1 U628 ( .A1(n563), .A2(n576), .ZN(n567) );
  XOR2_X1 U629 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n565) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(G204GAT), .B(KEYINPUT61), .Z(n570) );
  NAND2_X1 U634 ( .A1(n576), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1353GAT) );
  XOR2_X1 U636 ( .A(G211GAT), .B(KEYINPUT125), .Z(n573) );
  NAND2_X1 U637 ( .A1(n576), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1354GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n575) );
  XNOR2_X1 U640 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n580) );
  INV_X1 U642 ( .A(n576), .ZN(n577) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(n580), .B(n579), .Z(G1355GAT) );
endmodule

