//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT88), .Z(new_n204));
  XNOR2_X1  g003(.A(G211gat), .B(G218gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT74), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  AND2_X1   g007(.A1(G211gat), .A2(G218gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(KEYINPUT22), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n207), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT83), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G162gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n221));
  INV_X1    g020(.A(G148gat), .ZN(new_n222));
  NOR3_X1   g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G141gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(G148gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n219), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  AND2_X1   g025(.A1(KEYINPUT82), .A2(G155gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(KEYINPUT82), .A2(G155gat), .ZN(new_n228));
  OAI21_X1  g027(.A(G162gat), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n229), .A2(KEYINPUT2), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n213), .B1(new_n226), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT81), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n224), .ZN(new_n233));
  NAND2_X1  g032(.A1(KEYINPUT81), .A2(G141gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(G148gat), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n225), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n218), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n229), .A2(KEYINPUT2), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(KEYINPUT83), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n231), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G141gat), .B(G148gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n218), .B1(new_n241), .B2(KEYINPUT2), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT29), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n212), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT29), .B1(new_n210), .B2(new_n205), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n205), .B2(new_n210), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT89), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n244), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(new_n250), .B2(new_n249), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n252), .A2(new_n243), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n204), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G22gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n242), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n211), .B1(new_n257), .B2(KEYINPUT29), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n244), .B1(new_n211), .B2(KEYINPUT29), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n203), .B1(new_n259), .B2(new_n256), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n254), .A2(new_n255), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT90), .ZN(new_n263));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT31), .B(G50gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n254), .A2(new_n261), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G22gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(new_n262), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n263), .A2(new_n269), .A3(new_n262), .A4(new_n266), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT65), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT27), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G183gat), .ZN(new_n276));
  INV_X1    g075(.A(G183gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT27), .ZN(new_n278));
  INV_X1    g077(.A(G190gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n274), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n274), .A3(new_n281), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n276), .A2(new_n278), .A3(KEYINPUT28), .A4(new_n279), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT27), .B(G183gat), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n288), .A2(KEYINPUT66), .A3(KEYINPUT28), .A4(new_n279), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n283), .A2(new_n284), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G169gat), .ZN(new_n291));
  INV_X1    g090(.A(G176gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n293), .A2(KEYINPUT26), .A3(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n277), .A2(new_n279), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n294), .A2(KEYINPUT26), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n299), .B1(new_n301), .B2(new_n296), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT64), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT25), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT23), .B1(new_n291), .B2(new_n292), .ZN(new_n305));
  INV_X1    g104(.A(new_n294), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT23), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n302), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n308), .B1(new_n306), .B2(new_n305), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n312), .B(new_n302), .C1(new_n303), .C2(KEYINPUT25), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n290), .A2(new_n298), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(G127gat), .A2(G134gat), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT67), .B(G127gat), .Z(new_n316));
  AOI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(G134gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(G113gat), .B2(G120gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G113gat), .ZN(new_n321));
  INV_X1    g120(.A(G120gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT68), .B(G120gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G113gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(G127gat), .A2(G134gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n315), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n319), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n317), .A2(new_n323), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n313), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n284), .A2(new_n287), .A3(new_n289), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n298), .B1(new_n333), .B2(new_n282), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n329), .ZN(new_n336));
  NAND2_X1  g135(.A1(G227gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n331), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT32), .ZN(new_n340));
  XNOR2_X1  g139(.A(G15gat), .B(G43gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(G71gat), .B(G99gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT33), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n343), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT69), .B1(new_n339), .B2(new_n344), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n339), .A2(KEYINPUT69), .A3(new_n344), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n346), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n314), .A2(new_n330), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n335), .A2(new_n329), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n355), .A2(KEYINPUT34), .A3(new_n338), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT72), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT71), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n359), .B1(new_n353), .B2(new_n354), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n331), .A2(new_n336), .A3(KEYINPUT71), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n337), .A3(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n363));
  AOI21_X1  g162(.A(new_n358), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AND3_X1   g163(.A1(new_n362), .A2(new_n358), .A3(new_n363), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n352), .B(new_n357), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n367));
  INV_X1    g166(.A(new_n346), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n357), .B1(new_n365), .B2(new_n364), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n273), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT0), .ZN(new_n375));
  XNOR2_X1  g174(.A(G57gat), .B(G85gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  NAND2_X1  g176(.A1(new_n235), .A2(new_n236), .ZN(new_n378));
  AND4_X1   g177(.A1(KEYINPUT83), .A2(new_n238), .A3(new_n378), .A4(new_n219), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT83), .B1(new_n237), .B2(new_n238), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n242), .B(new_n329), .C1(new_n379), .C2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT85), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n240), .A2(KEYINPUT85), .A3(new_n242), .A4(new_n329), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT86), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT86), .A4(KEYINPUT4), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT84), .B(KEYINPUT4), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n243), .A2(new_n329), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n329), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n245), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(KEYINPUT5), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n391), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n389), .B1(new_n243), .B2(new_n329), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT4), .B1(new_n383), .B2(new_n384), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n393), .B(new_n394), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT5), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n383), .B(new_n384), .C1(new_n243), .C2(new_n329), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n401), .B1(new_n402), .B2(new_n395), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n377), .B1(new_n397), .B2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(KEYINPUT87), .B(KEYINPUT6), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n397), .A2(new_n377), .A3(new_n404), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n405), .A2(new_n407), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G226gat), .A2(G233gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(KEYINPUT75), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT76), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n332), .A2(new_n334), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n414), .B1(new_n332), .B2(new_n334), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n413), .B1(new_n417), .B2(new_n246), .ZN(new_n418));
  INV_X1    g217(.A(new_n413), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n314), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n211), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n335), .A2(KEYINPUT76), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n332), .A2(new_n334), .A3(new_n414), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n413), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT78), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT77), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT29), .B1(new_n332), .B2(new_n334), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n413), .ZN(new_n429));
  OAI211_X1 g228(.A(KEYINPUT77), .B(new_n419), .C1(new_n314), .C2(KEYINPUT29), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n422), .A2(KEYINPUT78), .A3(new_n413), .A4(new_n423), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n426), .A2(new_n431), .A3(new_n212), .A4(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(G8gat), .B(G36gat), .Z(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT79), .ZN(new_n435));
  XNOR2_X1  g234(.A(G64gat), .B(G92gat), .ZN(new_n436));
  XOR2_X1   g235(.A(new_n435), .B(new_n436), .Z(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT80), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT30), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n438), .B1(new_n421), .B2(new_n433), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n411), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n202), .B1(new_n373), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n445), .B1(new_n441), .B2(KEYINPUT30), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n451), .A2(KEYINPUT92), .A3(new_n444), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT92), .B1(new_n451), .B2(new_n444), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n366), .A2(new_n371), .A3(KEYINPUT73), .ZN(new_n455));
  OR3_X1    g254(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT73), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n271), .A2(new_n272), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n410), .A2(new_n409), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n405), .A2(new_n407), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT96), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT96), .B1(new_n405), .B2(new_n407), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n457), .A2(new_n202), .A3(new_n458), .A4(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n450), .B1(new_n454), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT36), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n366), .A2(new_n371), .A3(KEYINPUT73), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT73), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n273), .B1(new_n411), .B2(new_n447), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n467), .B1(new_n366), .B2(new_n371), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n472), .B1(new_n457), .B2(new_n467), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n477), .A2(KEYINPUT91), .A3(new_n471), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT37), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n421), .B2(new_n433), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n421), .A2(new_n480), .A3(new_n433), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n437), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT38), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n484), .A2(new_n439), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT38), .ZN(new_n486));
  AND4_X1   g285(.A1(new_n211), .A2(new_n426), .A3(new_n432), .A4(new_n431), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n422), .A2(new_n246), .A3(new_n423), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n420), .B1(new_n488), .B2(new_n419), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT37), .B1(new_n489), .B2(new_n211), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n486), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT95), .ZN(new_n492));
  OR3_X1    g291(.A1(new_n483), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n483), .B2(new_n491), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n485), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n458), .B1(new_n496), .B2(new_n464), .ZN(new_n497));
  NOR3_X1   g296(.A1(new_n452), .A2(new_n453), .A3(new_n405), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT39), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT93), .ZN(new_n500));
  AOI211_X1 g299(.A(new_n500), .B(new_n394), .C1(new_n391), .C2(new_n393), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n385), .A2(new_n386), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n388), .A2(new_n390), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n393), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT93), .B1(new_n504), .B2(new_n395), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n499), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n393), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n388), .A2(new_n390), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(new_n387), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n500), .B1(new_n509), .B2(new_n394), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n504), .A2(KEYINPUT93), .A3(new_n395), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n402), .A2(new_n395), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(new_n499), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n506), .A2(new_n377), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT40), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n506), .A2(new_n514), .A3(KEYINPUT40), .A4(new_n377), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n519), .A3(KEYINPUT94), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT94), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT92), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n447), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n405), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n451), .A2(KEYINPUT92), .A3(new_n444), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n517), .A2(new_n518), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n521), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n497), .B1(new_n520), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n466), .B1(new_n479), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n531), .A2(G1gat), .ZN(new_n532));
  INV_X1    g331(.A(G8gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT16), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n531), .B1(new_n534), .B2(G1gat), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n533), .B1(new_n532), .B2(new_n535), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT14), .ZN(new_n540));
  INV_X1    g339(.A(G29gat), .ZN(new_n541));
  INV_X1    g340(.A(G36gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n543), .A2(new_n544), .B1(G29gat), .B2(G36gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(G43gat), .B(G50gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT15), .ZN(new_n547));
  OR2_X1    g346(.A1(G43gat), .A2(G50gat), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549));
  NAND2_X1  g348(.A1(G43gat), .A2(G50gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n545), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT99), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n545), .A2(new_n547), .A3(KEYINPUT99), .A4(new_n551), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n544), .A2(KEYINPUT98), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n544), .A2(KEYINPUT98), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n543), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G29gat), .A2(G36gat), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n547), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n556), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n539), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n561), .B1(new_n554), .B2(new_n555), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n538), .B1(new_n566), .B2(KEYINPUT17), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT17), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n564), .B(new_n565), .C1(new_n567), .C2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT100), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n571), .A2(KEYINPUT18), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n563), .A2(new_n568), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n566), .A2(KEYINPUT17), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n576), .A3(new_n538), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n577), .A2(new_n564), .A3(new_n565), .A4(new_n572), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n565), .B(KEYINPUT13), .Z(new_n579));
  NOR2_X1   g378(.A1(new_n539), .A2(new_n563), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n566), .A2(new_n538), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT101), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(KEYINPUT101), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n574), .A2(new_n578), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G113gat), .B(G141gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(G197gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(KEYINPUT11), .B(G169gat), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT12), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n592), .B(KEYINPUT97), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n574), .A2(new_n578), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n584), .A2(new_n585), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n595), .A2(new_n596), .A3(new_n592), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(KEYINPUT102), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT102), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n599), .B1(new_n586), .B2(new_n592), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n594), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G134gat), .B(G162gat), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT106), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT7), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT7), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(G85gat), .A3(G92gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n607), .A2(new_n609), .B1(new_n605), .B2(new_n606), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT8), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(new_n612), .B2(KEYINPUT107), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(KEYINPUT107), .B2(new_n612), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(G99gat), .B(G106gat), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n610), .A2(new_n618), .A3(new_n614), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n575), .A2(new_n576), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  AND2_X1   g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n563), .A2(new_n622), .B1(KEYINPUT41), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(G190gat), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n621), .A2(new_n279), .A3(new_n624), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G218gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n623), .A2(KEYINPUT41), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n626), .A2(new_n627), .A3(G218gat), .ZN(new_n633));
  AND4_X1   g432(.A1(new_n604), .A2(new_n630), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT106), .B1(new_n628), .B2(new_n629), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n632), .B1(new_n635), .B2(new_n633), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n603), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n630), .A2(new_n604), .A3(new_n633), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n631), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n635), .A2(new_n632), .A3(new_n633), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n639), .A2(new_n602), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G71gat), .B(G78gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT103), .ZN(new_n645));
  XOR2_X1   g444(.A(G57gat), .B(G64gat), .Z(new_n646));
  INV_X1    g445(.A(KEYINPUT9), .ZN(new_n647));
  INV_X1    g446(.A(G71gat), .ZN(new_n648));
  INV_X1    g447(.A(G78gat), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n643), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n645), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n644), .A2(new_n646), .A3(KEYINPUT103), .A4(new_n650), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(KEYINPUT21), .ZN(new_n657));
  NAND2_X1  g456(.A1(G231gat), .A2(G233gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G127gat), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n654), .A2(KEYINPUT105), .A3(new_n655), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT105), .B1(new_n654), .B2(new_n655), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n539), .B1(new_n664), .B2(KEYINPUT21), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n660), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT104), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G155gat), .ZN(new_n669));
  XOR2_X1   g468(.A(G183gat), .B(G211gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n666), .B(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n642), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n620), .A2(new_n656), .ZN(new_n674));
  NAND2_X1  g473(.A1(G230gat), .A2(G233gat), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n617), .A2(new_n619), .B1(new_n654), .B2(new_n655), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n617), .A2(KEYINPUT10), .A3(new_n619), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n663), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT10), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(new_n674), .B2(new_n676), .ZN(new_n682));
  INV_X1    g481(.A(new_n679), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n683), .B(KEYINPUT108), .C1(new_n661), .C2(new_n662), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n680), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n677), .B1(new_n685), .B2(new_n675), .ZN(new_n686));
  XOR2_X1   g485(.A(G120gat), .B(G148gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT109), .ZN(new_n688));
  XNOR2_X1  g487(.A(G176gat), .B(G204gat), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n688), .B(new_n689), .Z(new_n690));
  OR2_X1    g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n686), .A2(KEYINPUT110), .A3(new_n690), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT110), .B1(new_n686), .B2(new_n690), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n673), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n530), .A2(new_n601), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT111), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT111), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n530), .A2(new_n700), .A3(new_n601), .A4(new_n697), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n411), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT112), .B(G1gat), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(G1324gat));
  INV_X1    g504(.A(new_n454), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT16), .B(G8gat), .ZN(new_n707));
  AOI211_X1 g506(.A(new_n706), .B(new_n707), .C1(new_n699), .C2(new_n701), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n708), .A2(KEYINPUT42), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n533), .B1(new_n702), .B2(new_n454), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT42), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(G1325gat));
  INV_X1    g511(.A(new_n457), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(G15gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n702), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(G15gat), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n477), .B1(new_n699), .B2(new_n701), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT113), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n715), .B(new_n720), .C1(new_n716), .C2(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(G1326gat));
  NAND2_X1  g521(.A1(new_n702), .A2(new_n273), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT43), .B(G22gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1327gat));
  AND2_X1   g524(.A1(new_n530), .A2(new_n601), .ZN(new_n726));
  INV_X1    g525(.A(new_n642), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n672), .A2(new_n695), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n726), .A2(new_n541), .A3(new_n411), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT45), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n466), .B1(new_n529), .B2(new_n474), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n642), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  AOI22_X1  g534(.A1(new_n733), .A2(new_n734), .B1(new_n530), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n597), .A2(KEYINPUT102), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n586), .A2(new_n599), .A3(new_n592), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n737), .A2(new_n738), .B1(new_n587), .B2(new_n593), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n728), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n411), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT114), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G29gat), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n741), .A2(KEYINPUT114), .A3(new_n742), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n731), .B1(new_n744), .B2(new_n745), .ZN(G1328gat));
  NAND4_X1  g545(.A1(new_n726), .A2(new_n542), .A3(new_n454), .A4(new_n729), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT46), .Z(new_n748));
  OAI21_X1  g547(.A(G36gat), .B1(new_n741), .B2(new_n706), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1329gat));
  INV_X1    g549(.A(new_n465), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n449), .B1(new_n751), .B2(new_n706), .ZN(new_n752));
  INV_X1    g551(.A(new_n497), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT94), .B1(new_n498), .B2(new_n519), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n526), .A2(new_n527), .A3(new_n521), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n474), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n752), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n734), .B1(new_n758), .B2(new_n727), .ZN(new_n759));
  INV_X1    g558(.A(new_n477), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n530), .A2(new_n735), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n759), .A2(new_n760), .A3(new_n761), .A4(new_n740), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G43gat), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n713), .A2(G43gat), .ZN(new_n764));
  AND4_X1   g563(.A1(new_n530), .A2(new_n601), .A3(new_n729), .A4(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT47), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n765), .B1(new_n762), .B2(G43gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n770), .A2(KEYINPUT115), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n769), .A2(new_n772), .ZN(G1330gat));
  NAND3_X1  g572(.A1(new_n726), .A2(new_n273), .A3(new_n729), .ZN(new_n774));
  INV_X1    g573(.A(G50gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n273), .A2(G50gat), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n741), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(KEYINPUT48), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n776), .B(new_n780), .C1(new_n741), .C2(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(G1331gat));
  NOR4_X1   g581(.A1(new_n642), .A2(new_n672), .A3(new_n601), .A4(new_n695), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n732), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n411), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g586(.A1(new_n784), .A2(new_n706), .ZN(new_n788));
  NOR2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  AND2_X1   g588(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n788), .B2(new_n789), .ZN(G1333gat));
  OAI21_X1  g591(.A(G71gat), .B1(new_n784), .B2(new_n477), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n457), .A2(new_n648), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n784), .B2(new_n794), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n795), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g595(.A1(new_n784), .A2(new_n458), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(new_n649), .ZN(G1335gat));
  NAND2_X1  g597(.A1(new_n672), .A2(new_n739), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n695), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT116), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n736), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G85gat), .B1(new_n802), .B2(new_n742), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n758), .A2(new_n727), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT117), .ZN(new_n805));
  INV_X1    g604(.A(new_n799), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n804), .A2(new_n805), .A3(KEYINPUT51), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n732), .A2(new_n642), .A3(new_n806), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT117), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n411), .A2(new_n605), .A3(new_n694), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n803), .B1(new_n813), .B2(new_n814), .ZN(G1336gat));
  NAND3_X1  g614(.A1(new_n736), .A2(new_n454), .A3(new_n801), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(new_n816), .B2(G92gat), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n706), .A2(G92gat), .A3(new_n695), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT52), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n808), .A2(new_n822), .A3(KEYINPUT51), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT51), .B1(new_n808), .B2(new_n822), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI22_X1  g624(.A1(new_n825), .A2(new_n818), .B1(new_n816), .B2(G92gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n820), .B1(new_n821), .B2(new_n826), .ZN(G1337gat));
  XOR2_X1   g626(.A(KEYINPUT119), .B(G99gat), .Z(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n802), .B2(new_n477), .ZN(new_n829));
  OR3_X1    g628(.A1(new_n713), .A2(new_n695), .A3(new_n828), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n829), .B1(new_n813), .B2(new_n830), .ZN(G1338gat));
  NOR3_X1   g630(.A1(new_n458), .A2(G106gat), .A3(new_n695), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT53), .B1(new_n812), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n736), .A2(new_n834), .A3(new_n273), .A4(new_n801), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n759), .A2(new_n273), .A3(new_n761), .A4(new_n801), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT121), .ZN(new_n837));
  XNOR2_X1  g636(.A(KEYINPUT120), .B(G106gat), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n833), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n832), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n823), .A2(new_n824), .A3(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n836), .A2(new_n839), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT53), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n845), .ZN(G1339gat));
  NOR2_X1   g645(.A1(new_n696), .A2(new_n601), .ZN(new_n847));
  INV_X1    g646(.A(new_n672), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n565), .B1(new_n577), .B2(new_n564), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n580), .A2(new_n581), .A3(new_n579), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n591), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n694), .B(new_n852), .C1(new_n598), .C2(new_n600), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n685), .A2(new_n675), .ZN(new_n855));
  INV_X1    g654(.A(new_n675), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n680), .A2(new_n684), .A3(new_n856), .A4(new_n682), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n855), .A2(KEYINPUT54), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n685), .A2(new_n859), .A3(new_n675), .ZN(new_n860));
  INV_X1    g659(.A(new_n690), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n854), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n677), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n855), .A2(new_n864), .A3(new_n690), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT110), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n686), .A2(KEYINPUT110), .A3(new_n690), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n855), .A2(KEYINPUT54), .A3(new_n857), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n870), .A2(KEYINPUT55), .A3(new_n861), .A4(new_n860), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n863), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n853), .B1(new_n739), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(new_n641), .A3(new_n637), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n863), .A2(new_n869), .A3(new_n871), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n737), .A2(new_n738), .B1(new_n591), .B2(new_n851), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n642), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n848), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n847), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(new_n742), .A3(new_n454), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n713), .A2(new_n273), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(new_n321), .A3(new_n739), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n880), .A2(new_n373), .A3(new_n601), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n321), .B2(new_n884), .ZN(G1340gat));
  OAI21_X1  g684(.A(G120gat), .B1(new_n882), .B2(new_n695), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n880), .A2(new_n373), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n695), .A2(new_n324), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n889), .B(KEYINPUT122), .Z(G1341gat));
  OAI21_X1  g689(.A(new_n316), .B1(new_n882), .B2(new_n672), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n672), .A2(new_n316), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n887), .B2(new_n892), .ZN(G1342gat));
  NOR2_X1   g692(.A1(new_n879), .A2(new_n742), .ZN(new_n894));
  INV_X1    g693(.A(G134gat), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n454), .A2(new_n727), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n894), .A2(new_n895), .A3(new_n373), .A4(new_n896), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n897), .B(KEYINPUT56), .Z(new_n898));
  OAI21_X1  g697(.A(G134gat), .B1(new_n882), .B2(new_n727), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1343gat));
  OAI21_X1  g699(.A(new_n273), .B1(new_n847), .B2(new_n878), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT57), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n454), .A2(new_n742), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n477), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n902), .A2(new_n739), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n220), .A2(new_n221), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n894), .A2(KEYINPUT123), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n894), .A2(KEYINPUT123), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n760), .A2(new_n458), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n908), .A2(new_n706), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n601), .A2(new_n224), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT58), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n915));
  OAI221_X1 g714(.A(new_n915), .B1(new_n911), .B2(new_n912), .C1(new_n905), .C2(new_n906), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1344gat));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n875), .A2(new_n601), .B1(new_n876), .B2(new_n694), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n642), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n870), .A2(new_n861), .A3(new_n860), .ZN(new_n921));
  AOI22_X1  g720(.A1(new_n921), .A2(new_n854), .B1(new_n867), .B2(new_n868), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n876), .A2(new_n871), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n923), .B1(new_n641), .B2(new_n637), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT124), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n874), .A2(new_n877), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n925), .A2(new_n927), .A3(new_n672), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n697), .A2(new_n739), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT57), .B1(new_n930), .B2(new_n273), .ZN(new_n931));
  OAI211_X1 g730(.A(KEYINPUT57), .B(new_n273), .C1(new_n847), .C2(new_n878), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n934), .A2(new_n477), .A3(new_n694), .A4(new_n903), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n918), .B1(new_n935), .B2(G148gat), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n902), .A2(new_n695), .A3(new_n904), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(KEYINPUT59), .A3(new_n222), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n694), .A2(new_n222), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n936), .A2(new_n938), .B1(new_n911), .B2(new_n939), .ZN(G1345gat));
  NOR3_X1   g739(.A1(new_n902), .A2(new_n672), .A3(new_n904), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n227), .A2(new_n228), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n848), .A2(new_n943), .ZN(new_n944));
  OAI22_X1  g743(.A1(new_n941), .A2(new_n943), .B1(new_n911), .B2(new_n944), .ZN(G1346gat));
  NOR3_X1   g744(.A1(new_n902), .A2(new_n727), .A3(new_n904), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n896), .A2(new_n214), .ZN(new_n948));
  OAI22_X1  g747(.A1(new_n946), .A2(new_n214), .B1(new_n947), .B2(new_n948), .ZN(G1347gat));
  NOR2_X1   g748(.A1(new_n879), .A2(new_n411), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n454), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n951), .A2(new_n273), .A3(new_n372), .ZN(new_n952));
  AOI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n601), .ZN(new_n953));
  INV_X1    g752(.A(new_n881), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n739), .A2(new_n291), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1348gat));
  NAND3_X1  g756(.A1(new_n952), .A2(new_n292), .A3(new_n694), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n951), .A2(new_n954), .A3(new_n695), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n292), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT125), .ZN(G1349gat));
  NAND3_X1  g760(.A1(new_n952), .A2(new_n288), .A3(new_n848), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n951), .A2(new_n954), .A3(new_n672), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n277), .B2(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g764(.A1(new_n952), .A2(new_n279), .A3(new_n642), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n955), .A2(new_n642), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(G190gat), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(G1351gat));
  NAND2_X1  g770(.A1(new_n910), .A2(new_n454), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n972), .A2(KEYINPUT126), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(KEYINPUT126), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n973), .A2(new_n950), .A3(new_n974), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(G197gat), .B1(new_n976), .B2(new_n601), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n760), .A2(new_n411), .A3(new_n706), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n934), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n601), .A2(G197gat), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(G1352gat));
  NOR3_X1   g780(.A1(new_n975), .A2(G204gat), .A3(new_n695), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT62), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n934), .A2(new_n694), .A3(new_n978), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G204gat), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(new_n985), .ZN(G1353gat));
  INV_X1    g785(.A(G211gat), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n976), .A2(new_n987), .A3(new_n848), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n848), .B(new_n978), .C1(new_n931), .C2(new_n933), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n989), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n990));
  AOI21_X1  g789(.A(KEYINPUT63), .B1(new_n989), .B2(G211gat), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI211_X1 g793(.A(KEYINPUT127), .B(new_n988), .C1(new_n990), .C2(new_n991), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(G1354gat));
  NAND3_X1  g795(.A1(new_n976), .A2(new_n629), .A3(new_n642), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n979), .A2(new_n642), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n997), .B1(new_n998), .B2(new_n629), .ZN(G1355gat));
endmodule


