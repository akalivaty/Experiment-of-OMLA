//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(G120gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G113gat), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G120gat), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT1), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G134gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G127gat), .ZN(new_n210));
  INV_X1    g009(.A(G127gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G134gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n208), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT69), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(new_n212), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n210), .A2(new_n215), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n205), .A2(new_n207), .ZN(new_n219));
  OAI22_X1  g018(.A1(new_n217), .A2(new_n218), .B1(new_n219), .B2(KEYINPUT1), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT69), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n208), .A2(new_n221), .A3(new_n210), .A4(new_n212), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n214), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(G155gat), .ZN(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G141gat), .B(G148gat), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n224), .B(new_n227), .C1(new_n228), .C2(KEYINPUT75), .ZN(new_n229));
  INV_X1    g028(.A(G148gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G141gat), .ZN(new_n231));
  INV_X1    g030(.A(G141gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G148gat), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n231), .A2(new_n233), .B1(KEYINPUT2), .B2(new_n224), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n229), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(new_n233), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n224), .A2(KEYINPUT2), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT75), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n232), .A2(G148gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n230), .A2(G141gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n238), .A2(new_n242), .A3(new_n224), .A4(new_n227), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n235), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n223), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT4), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n235), .A2(new_n243), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n235), .B2(new_n243), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n248), .B1(new_n252), .B2(new_n223), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n203), .B(new_n246), .C1(new_n253), .C2(new_n245), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n214), .A2(new_n220), .A3(new_n222), .ZN(new_n255));
  INV_X1    g054(.A(new_n244), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n223), .A2(new_n244), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n203), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n254), .A2(KEYINPUT5), .A3(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n236), .A2(new_n239), .B1(G155gat), .B2(G162gat), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n238), .B1(new_n263), .B2(new_n227), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n229), .A2(new_n234), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT3), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n235), .A2(new_n243), .A3(new_n249), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n223), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(KEYINPUT4), .A3(new_n257), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n245), .A2(new_n248), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n203), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G1gat), .B(G29gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT0), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(G57gat), .ZN(new_n277));
  INV_X1    g076(.A(G85gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n262), .A2(new_n279), .A3(new_n273), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n281), .A2(KEYINPUT77), .A3(new_n282), .A4(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT77), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n274), .B(new_n280), .C1(new_n285), .C2(KEYINPUT6), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OR2_X1    g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(KEYINPUT66), .B2(KEYINPUT24), .ZN(new_n291));
  AND2_X1   g090(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n288), .B(new_n289), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n294), .A2(G169gat), .A3(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(G169gat), .ZN(new_n296));
  INV_X1    g095(.A(G176gat), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT65), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT23), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT23), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n296), .A2(new_n297), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n293), .A2(new_n299), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT64), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n306), .A2(new_n288), .A3(new_n307), .A4(new_n289), .ZN(new_n308));
  NOR2_X1   g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT25), .B1(new_n309), .B2(KEYINPUT23), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(new_n288), .A3(new_n289), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n312), .A2(KEYINPUT64), .B1(new_n302), .B2(new_n301), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n304), .A2(KEYINPUT25), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT67), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(new_n309), .ZN(new_n317));
  INV_X1    g116(.A(new_n316), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n318), .A2(KEYINPUT67), .A3(new_n302), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n295), .A2(new_n298), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n317), .B(new_n319), .C1(new_n320), .C2(KEYINPUT26), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT27), .B(G183gat), .ZN(new_n322));
  INV_X1    g121(.A(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT28), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT28), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n322), .A2(new_n326), .A3(new_n323), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n321), .A2(new_n290), .A3(new_n325), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n314), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT73), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n330), .A2(G226gat), .A3(G233gat), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G226gat), .A2(G233gat), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n334), .B(KEYINPUT72), .Z(new_n335));
  INV_X1    g134(.A(new_n329), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(KEYINPUT29), .ZN(new_n337));
  XNOR2_X1  g136(.A(G197gat), .B(G204gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT22), .ZN(new_n339));
  INV_X1    g138(.A(G211gat), .ZN(new_n340));
  INV_X1    g139(.A(G218gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G211gat), .B(G218gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n338), .A3(new_n342), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n337), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n336), .A2(new_n335), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT29), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n330), .A2(new_n352), .A3(new_n332), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n353), .B2(new_n334), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n350), .B1(new_n354), .B2(new_n349), .ZN(new_n355));
  XOR2_X1   g154(.A(G8gat), .B(G36gat), .Z(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(G64gat), .ZN(new_n357));
  INV_X1    g156(.A(G92gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT30), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT30), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n355), .A2(new_n363), .A3(new_n360), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n350), .B(new_n359), .C1(new_n354), .C2(new_n349), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT74), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n366), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n362), .A2(new_n364), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT31), .B(G50gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G78gat), .B(G106gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n267), .A2(new_n376), .A3(new_n352), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n376), .B1(new_n267), .B2(new_n352), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n377), .A2(new_n378), .A3(new_n348), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT3), .B1(new_n348), .B2(new_n352), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n256), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n375), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n380), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n244), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT79), .B1(new_n256), .B2(new_n380), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n267), .A2(new_n352), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n349), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n385), .A2(new_n386), .A3(new_n388), .A4(new_n374), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT78), .B1(new_n390), .B2(G22gat), .ZN(new_n391));
  INV_X1    g190(.A(G22gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n382), .A2(new_n392), .A3(new_n389), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n373), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT78), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n387), .A2(KEYINPUT80), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n267), .A2(new_n376), .A3(new_n352), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n349), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n381), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n374), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AND4_X1   g199(.A1(new_n374), .A2(new_n385), .A3(new_n386), .A4(new_n388), .ZN(new_n401));
  OAI21_X1  g200(.A(G22gat), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND4_X1   g201(.A1(new_n395), .A2(new_n402), .A3(new_n373), .A4(new_n393), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n371), .B1(new_n394), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n391), .A2(new_n373), .A3(new_n393), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n393), .A3(new_n395), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n372), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n407), .A3(new_n370), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n287), .A2(new_n369), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT36), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n329), .A2(new_n255), .ZN(new_n411));
  INV_X1    g210(.A(G227gat), .ZN(new_n412));
  INV_X1    g211(.A(G233gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n314), .A2(new_n328), .A3(new_n223), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT32), .ZN(new_n417));
  XOR2_X1   g216(.A(KEYINPUT70), .B(KEYINPUT33), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G15gat), .B(G43gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(G71gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(G99gat), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n417), .A2(new_n420), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n411), .A2(new_n415), .ZN(new_n426));
  INV_X1    g225(.A(new_n414), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(KEYINPUT71), .A3(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n416), .B(KEYINPUT32), .C1(new_n419), .C2(new_n423), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n425), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n428), .B1(new_n425), .B2(new_n429), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT71), .B1(new_n426), .B2(new_n427), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n433), .A2(KEYINPUT34), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n431), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n425), .A2(new_n429), .ZN(new_n437));
  INV_X1    g236(.A(new_n428), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n439), .B2(new_n430), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n410), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n435), .B1(new_n431), .B2(new_n432), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(new_n434), .A3(new_n430), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT36), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n409), .A2(new_n445), .ZN(new_n446));
  AOI211_X1 g245(.A(KEYINPUT5), .B(new_n260), .C1(new_n269), .C2(new_n270), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n268), .A2(new_n247), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n260), .B1(new_n448), .B2(new_n257), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n272), .B1(new_n449), .B2(new_n246), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n447), .B1(new_n450), .B2(new_n261), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT83), .ZN(new_n452));
  NOR4_X1   g251(.A1(new_n451), .A2(new_n452), .A3(new_n282), .A4(new_n279), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n279), .B1(new_n262), .B2(new_n273), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT83), .B1(new_n454), .B2(KEYINPUT6), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n283), .A2(new_n282), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n454), .A2(KEYINPUT81), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n460));
  AOI211_X1 g259(.A(new_n460), .B(new_n279), .C1(new_n262), .C2(new_n273), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n458), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n354), .A2(new_n349), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n333), .A2(new_n337), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n463), .B(KEYINPUT37), .C1(new_n349), .C2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(KEYINPUT82), .B(KEYINPUT37), .Z(new_n466));
  NAND2_X1  g265(.A1(new_n355), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n465), .A2(new_n467), .A3(new_n468), .A4(new_n359), .ZN(new_n469));
  INV_X1    g268(.A(new_n361), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT37), .B(new_n350), .C1(new_n354), .C2(new_n349), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n359), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n472), .B2(KEYINPUT38), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n456), .A2(new_n462), .A3(new_n469), .A4(new_n473), .ZN(new_n474));
  AND2_X1   g273(.A1(new_n404), .A2(new_n408), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n362), .A2(new_n364), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n367), .A2(new_n368), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n460), .B1(new_n451), .B2(new_n279), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n454), .A2(KEYINPUT81), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n269), .A2(new_n260), .A3(new_n270), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n482), .B(KEYINPUT39), .C1(new_n260), .C2(new_n259), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n483), .B(new_n279), .C1(KEYINPUT39), .C2(new_n482), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT40), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n478), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n474), .A2(new_n475), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n274), .A2(KEYINPUT6), .A3(new_n280), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n452), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n454), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n457), .B1(new_n479), .B2(new_n480), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n369), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT35), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n442), .A2(new_n443), .ZN(new_n497));
  AND4_X1   g296(.A1(new_n496), .A2(new_n497), .A3(new_n404), .A4(new_n408), .ZN(new_n498));
  OAI211_X1 g297(.A(KEYINPUT84), .B(new_n369), .C1(new_n491), .C2(new_n492), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n497), .A2(new_n404), .A3(new_n408), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n287), .A2(new_n369), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT35), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI221_X4 g302(.A(new_n202), .B1(new_n446), .B2(new_n487), .C1(new_n500), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n500), .A2(new_n503), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n446), .A2(new_n487), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT85), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508));
  OR3_X1    g307(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(KEYINPUT86), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n511), .B1(KEYINPUT86), .B2(new_n510), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT87), .B(G29gat), .ZN(new_n513));
  INV_X1    g312(.A(G36gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(KEYINPUT15), .B(new_n508), .C1(new_n512), .C2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n509), .B1(new_n515), .B2(new_n510), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n508), .A2(KEYINPUT15), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT88), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT88), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n516), .A2(new_n523), .A3(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(G15gat), .B(G22gat), .Z(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  OR3_X1    g327(.A1(new_n527), .A2(KEYINPUT89), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n527), .B2(KEYINPUT89), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n529), .B(new_n530), .C1(KEYINPUT16), .C2(new_n527), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G8gat), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n522), .A2(new_n535), .A3(new_n524), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT17), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n532), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G229gat), .A2(G233gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT18), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(KEYINPUT90), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n540), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n534), .A2(new_n538), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT90), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT18), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n525), .B(new_n532), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n540), .B(KEYINPUT91), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT13), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n543), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(G197gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT11), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(new_n296), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT12), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n543), .A2(new_n547), .A3(new_n557), .A4(new_n551), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT99), .ZN(new_n563));
  XOR2_X1   g362(.A(G57gat), .B(G64gat), .Z(new_n564));
  NAND2_X1  g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(KEYINPUT9), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G71gat), .B(G78gat), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n568), .A2(KEYINPUT92), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(KEYINPUT92), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT93), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n564), .B(new_n568), .C1(KEYINPUT9), .C2(new_n566), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n567), .B(KEYINPUT93), .C1(new_n569), .C2(new_n570), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G99gat), .B(G106gat), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT97), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(KEYINPUT8), .A2(new_n580), .B1(new_n278), .B2(new_n358), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT7), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n577), .B(KEYINPUT97), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n581), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n563), .B(KEYINPUT10), .C1(new_n576), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(KEYINPUT98), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n588), .B1(new_n576), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n594));
  NOR3_X1   g393(.A1(new_n576), .A2(new_n591), .A3(new_n588), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n594), .B1(new_n595), .B2(KEYINPUT99), .ZN(new_n596));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n593), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n595), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n599), .A2(new_n592), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G120gat), .B(G148gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n297), .ZN(new_n603));
  INV_X1    g402(.A(G204gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT100), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n601), .A2(new_n605), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n601), .A2(KEYINPUT100), .A3(new_n605), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n562), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(G162gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n536), .A2(new_n537), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n588), .ZN(new_n620));
  NAND3_X1  g419(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n620), .B(new_n621), .C1(new_n526), .C2(new_n588), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G134gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n622), .B(new_n209), .ZN(new_n626));
  INV_X1    g425(.A(new_n624), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n618), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n623), .A2(new_n624), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n617), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT21), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n533), .B1(new_n634), .B2(new_n576), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n576), .A2(new_n634), .ZN(new_n638));
  XOR2_X1   g437(.A(G183gat), .B(G211gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G127gat), .B(G155gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT20), .ZN(new_n643));
  NAND2_X1  g442(.A1(G231gat), .A2(G233gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n641), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n648), .ZN(new_n649));
  NOR4_X1   g448(.A1(new_n504), .A2(new_n507), .A3(new_n615), .A4(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n287), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT101), .B(G1gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(G1324gat));
  NAND2_X1  g453(.A1(new_n650), .A2(new_n478), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n655), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(G8gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  MUX2_X1   g460(.A(new_n659), .B(new_n661), .S(KEYINPUT42), .Z(G1325gat));
  AOI21_X1  g461(.A(G15gat), .B1(new_n650), .B2(new_n497), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n445), .A2(G15gat), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n663), .B1(new_n650), .B2(new_n664), .ZN(G1326gat));
  INV_X1    g464(.A(new_n475), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n504), .A2(new_n507), .ZN(new_n670));
  INV_X1    g469(.A(new_n648), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n629), .A2(new_n632), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n670), .A2(new_n614), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n651), .A3(new_n513), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n648), .B(KEYINPUT103), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n614), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n505), .A2(new_n506), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n202), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n505), .A2(KEYINPUT85), .A3(new_n506), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n682), .A2(new_n683), .A3(new_n672), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT44), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n506), .A2(KEYINPUT104), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n446), .A2(new_n487), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n633), .B1(new_n689), .B2(new_n505), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n680), .B1(new_n685), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n287), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n677), .B1(new_n513), .B2(new_n695), .ZN(G1328gat));
  NAND2_X1  g495(.A1(new_n674), .A2(new_n514), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT46), .B1(new_n697), .B2(new_n369), .ZN(new_n698));
  OAI21_X1  g497(.A(G36gat), .B1(new_n694), .B2(new_n369), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n697), .A2(KEYINPUT46), .A3(new_n369), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n700), .A2(KEYINPUT106), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(KEYINPUT106), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n698), .B(new_n699), .C1(new_n701), .C2(new_n702), .ZN(G1329gat));
  INV_X1    g502(.A(new_n445), .ZN(new_n704));
  OAI21_X1  g503(.A(G43gat), .B1(new_n694), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n673), .A2(G43gat), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(new_n497), .ZN(new_n708));
  INV_X1    g507(.A(new_n497), .ZN(new_n709));
  NOR4_X1   g508(.A1(new_n673), .A2(KEYINPUT107), .A3(G43gat), .A4(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n705), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g512(.A(new_n705), .B(KEYINPUT47), .C1(new_n708), .C2(new_n710), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1330gat));
  NOR2_X1   g514(.A1(new_n475), .A2(G50gat), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  AOI211_X1 g516(.A(new_n475), .B(new_n680), .C1(new_n685), .C2(new_n692), .ZN(new_n718));
  INV_X1    g517(.A(G50gat), .ZN(new_n719));
  OAI221_X1 g518(.A(KEYINPUT48), .B1(new_n673), .B2(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT108), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n673), .B2(new_n717), .ZN(new_n723));
  NOR4_X1   g522(.A1(new_n504), .A2(new_n507), .A3(new_n615), .A4(new_n633), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n724), .A2(KEYINPUT108), .A3(new_n671), .A4(new_n716), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n723), .B(new_n725), .C1(new_n718), .C2(new_n719), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT48), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n721), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n719), .B1(new_n693), .B2(new_n666), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n723), .A2(new_n725), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n721), .B(new_n727), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n720), .B1(new_n728), .B2(new_n732), .ZN(G1331gat));
  NAND2_X1  g532(.A1(new_n689), .A2(new_n505), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n649), .A2(new_n561), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(new_n613), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n287), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g537(.A(new_n736), .B(KEYINPUT110), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n478), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT49), .B(G64gat), .Z(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(G1333gat));
  INV_X1    g542(.A(G71gat), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n739), .B2(new_n445), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746));
  OR3_X1    g545(.A1(new_n736), .A2(new_n746), .A3(new_n709), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n736), .B2(new_n709), .ZN(new_n748));
  AOI21_X1  g547(.A(G71gat), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g550(.A1(new_n739), .A2(new_n666), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g552(.A1(new_n685), .A2(new_n692), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n671), .A2(new_n562), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT112), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(new_n613), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(G85gat), .B1(new_n757), .B2(new_n287), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n690), .A2(KEYINPUT51), .A3(new_n756), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n759), .A2(KEYINPUT113), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n690), .A2(new_n756), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n763), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n613), .A2(new_n278), .A3(new_n651), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT114), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n758), .B1(new_n766), .B2(new_n768), .ZN(G1336gat));
  NAND4_X1  g568(.A1(new_n754), .A2(new_n613), .A3(new_n478), .A4(new_n756), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT52), .B1(new_n770), .B2(G92gat), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n612), .A2(new_n369), .A3(G92gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n764), .A2(new_n765), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(new_n763), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n777), .A2(new_n772), .B1(G92gat), .B2(new_n770), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n774), .B1(new_n778), .B2(new_n779), .ZN(G1337gat));
  OAI21_X1  g579(.A(G99gat), .B1(new_n757), .B2(new_n704), .ZN(new_n781));
  OR3_X1    g580(.A1(new_n612), .A2(new_n709), .A3(G99gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n766), .B2(new_n782), .ZN(G1338gat));
  NOR3_X1   g582(.A1(new_n475), .A2(new_n612), .A3(G106gat), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n764), .A2(new_n765), .A3(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n754), .A2(new_n613), .A3(new_n666), .A4(new_n756), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  XOR2_X1   g586(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n788));
  NAND3_X1  g587(.A1(new_n785), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n777), .A2(new_n784), .B1(G106gat), .B2(new_n786), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(G1339gat));
  NAND2_X1  g591(.A1(new_n593), .A2(new_n596), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(G230gat), .A3(G233gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(KEYINPUT54), .A3(new_n598), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n593), .A2(new_n596), .A3(new_n796), .A4(new_n597), .ZN(new_n797));
  AND3_X1   g596(.A1(new_n797), .A2(KEYINPUT117), .A3(new_n605), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT117), .B1(new_n797), .B2(new_n605), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n607), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(KEYINPUT118), .B(new_n607), .C1(new_n800), .C2(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n800), .A2(new_n801), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n804), .A2(new_n561), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  OAI22_X1  g606(.A1(new_n539), .A2(new_n540), .B1(new_n548), .B2(new_n550), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n556), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n560), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n613), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n633), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n804), .A2(new_n805), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n814), .A2(new_n672), .A3(new_n810), .A4(new_n806), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n678), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n649), .A2(new_n561), .A3(new_n613), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n287), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n501), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT119), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n561), .A2(new_n206), .ZN(new_n824));
  XOR2_X1   g623(.A(new_n824), .B(KEYINPUT120), .Z(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n369), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n822), .A2(new_n478), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(G113gat), .B1(new_n828), .B2(new_n562), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n826), .A2(new_n829), .ZN(G1340gat));
  NAND4_X1  g629(.A1(new_n823), .A2(new_n204), .A3(new_n613), .A4(new_n369), .ZN(new_n831));
  OAI21_X1  g630(.A(G120gat), .B1(new_n828), .B2(new_n612), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1341gat));
  NAND3_X1  g632(.A1(new_n823), .A2(new_n369), .A3(new_n648), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n679), .A2(new_n211), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n834), .A2(new_n211), .B1(new_n827), .B2(new_n835), .ZN(G1342gat));
  NOR2_X1   g635(.A1(new_n633), .A2(new_n478), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n823), .A2(new_n209), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT56), .ZN(new_n839));
  INV_X1    g638(.A(new_n837), .ZN(new_n840));
  OAI21_X1  g639(.A(G134gat), .B1(new_n822), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT56), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n823), .A2(new_n842), .A3(new_n209), .A4(new_n837), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n839), .A2(new_n841), .A3(new_n843), .ZN(G1343gat));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n845), .B(new_n666), .C1(new_n816), .C2(new_n818), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n704), .A2(new_n651), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n478), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n800), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n795), .B(KEYINPUT121), .C1(new_n798), .C2(new_n799), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n801), .A3(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n802), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n851), .A2(KEYINPUT122), .A3(new_n801), .A4(new_n852), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n855), .A2(new_n856), .A3(new_n561), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n811), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n858), .A2(KEYINPUT123), .A3(new_n811), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n633), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n648), .B1(new_n863), .B2(new_n815), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n666), .B1(new_n864), .B2(new_n818), .ZN(new_n865));
  AOI211_X1 g664(.A(new_n562), .B(new_n849), .C1(new_n865), .C2(KEYINPUT57), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT124), .B1(new_n866), .B2(new_n232), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n817), .A2(new_n819), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n666), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n869), .A2(new_n478), .A3(new_n847), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n232), .A3(new_n561), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n866), .B2(new_n232), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n867), .A2(new_n872), .A3(KEYINPUT58), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  OAI221_X1 g673(.A(new_n871), .B1(KEYINPUT124), .B2(new_n874), .C1(new_n866), .C2(new_n232), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1344gat));
  NAND3_X1  g675(.A1(new_n870), .A2(new_n230), .A3(new_n613), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n849), .B1(new_n865), .B2(KEYINPUT57), .ZN(new_n878));
  AOI211_X1 g677(.A(KEYINPUT59), .B(new_n230), .C1(new_n878), .C2(new_n613), .ZN(new_n879));
  XNOR2_X1  g678(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n869), .A2(KEYINPUT57), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n845), .B(new_n666), .C1(new_n864), .C2(new_n818), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n881), .A2(new_n882), .A3(new_n613), .A4(new_n848), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n883), .B2(G148gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n877), .B1(new_n879), .B2(new_n884), .ZN(G1345gat));
  INV_X1    g684(.A(new_n878), .ZN(new_n886));
  OAI21_X1  g685(.A(G155gat), .B1(new_n886), .B2(new_n679), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n225), .A3(new_n648), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1346gat));
  OAI21_X1  g688(.A(G162gat), .B1(new_n886), .B2(new_n633), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n837), .A2(new_n226), .A3(new_n651), .A4(new_n704), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n869), .B2(new_n891), .ZN(G1347gat));
  NOR2_X1   g691(.A1(new_n651), .A2(new_n369), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n868), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n821), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n562), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(new_n296), .ZN(G1348gat));
  NOR2_X1   g696(.A1(new_n895), .A2(new_n612), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(new_n297), .ZN(G1349gat));
  OAI21_X1  g698(.A(G183gat), .B1(new_n895), .B2(new_n679), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n648), .A2(new_n322), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n895), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT60), .ZN(G1350gat));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G190gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n895), .A2(new_n633), .ZN(new_n906));
  MUX2_X1   g705(.A(new_n904), .B(new_n905), .S(new_n906), .Z(G1351gat));
  AND2_X1   g706(.A1(new_n881), .A2(new_n882), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n704), .A2(new_n893), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n561), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(KEYINPUT126), .B(G197gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n869), .A2(new_n909), .ZN(new_n914));
  INV_X1    g713(.A(new_n912), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n561), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n913), .A2(new_n916), .ZN(G1352gat));
  NOR3_X1   g716(.A1(new_n475), .A2(new_n612), .A3(G204gat), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n868), .A2(new_n910), .A3(new_n918), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n919), .B(KEYINPUT62), .Z(new_n920));
  AND3_X1   g719(.A1(new_n908), .A2(new_n613), .A3(new_n910), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n604), .ZN(G1353gat));
  NAND4_X1  g721(.A1(new_n881), .A2(new_n882), .A3(new_n648), .A4(new_n910), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G211gat), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(KEYINPUT63), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(KEYINPUT63), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n914), .A2(new_n340), .A3(new_n648), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT127), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(G1354gat));
  AOI21_X1  g728(.A(G218gat), .B1(new_n914), .B2(new_n672), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n908), .A2(new_n910), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n633), .A2(new_n341), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(G1355gat));
endmodule


