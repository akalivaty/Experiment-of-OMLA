//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1320, new_n1321,
    new_n1322, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n201), .B(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  AND2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NOR2_X1   g0009(.A1(G58), .A2(G68), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(G13), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT0), .Z(new_n221));
  INV_X1    g0021(.A(KEYINPUT65), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n217), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(new_n222), .B2(new_n221), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT66), .Z(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT67), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n218), .B1(new_n227), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n225), .A2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(KEYINPUT71), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n215), .A2(G1), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  AND3_X1   g0055(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n214), .ZN(new_n256));
  AOI21_X1  g0056(.A(KEYINPUT70), .B1(new_n255), .B2(new_n214), .ZN(new_n257));
  OR2_X1    g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n254), .A2(new_n261), .B1(new_n251), .B2(new_n260), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(KEYINPUT7), .B1(new_n265), .B2(new_n215), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT7), .ZN(new_n267));
  NOR4_X1   g0067(.A1(new_n263), .A2(new_n264), .A3(new_n267), .A4(G20), .ZN(new_n268));
  OAI21_X1  g0068(.A(G68), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G58), .ZN(new_n270));
  INV_X1    g0070(.A(G68), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(G20), .B1(new_n272), .B2(new_n210), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G159), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n269), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT16), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n258), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n269), .A2(KEYINPUT16), .A3(new_n277), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n262), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G169), .ZN(new_n283));
  OR2_X1    g0083(.A1(G223), .A2(G1698), .ZN(new_n284));
  INV_X1    g0084(.A(G226), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G1698), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n284), .B(new_n286), .C1(new_n263), .C2(new_n264), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G87), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G41), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G1), .A3(G13), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  INV_X1    g0094(.A(G45), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(G1), .A2(G13), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n259), .A2(new_n296), .B1(new_n297), .B2(new_n290), .ZN(new_n298));
  INV_X1    g0098(.A(G274), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n297), .B2(new_n290), .ZN(new_n300));
  AOI21_X1  g0100(.A(G1), .B1(new_n294), .B2(new_n295), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n298), .A2(G232), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT75), .B1(new_n293), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n291), .B1(new_n287), .B2(new_n288), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n301), .A2(new_n291), .A3(G274), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n291), .A2(G232), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT75), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n304), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n283), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n304), .A2(new_n308), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT18), .B1(new_n282), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G200), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n303), .B2(new_n310), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n304), .A2(new_n308), .A3(G190), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n282), .A2(KEYINPUT17), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT17), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT3), .B(G33), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n267), .B1(new_n324), .B2(G20), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n215), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n271), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n279), .B1(new_n327), .B2(new_n276), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n256), .A2(new_n257), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n281), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT71), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n250), .B(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n332), .A2(new_n252), .ZN(new_n333));
  INV_X1    g0133(.A(new_n260), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n333), .A2(new_n335), .B1(new_n332), .B2(new_n334), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n293), .A2(KEYINPUT75), .A3(new_n302), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n309), .B1(new_n304), .B2(new_n308), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n319), .B1(new_n340), .B2(new_n317), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n323), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n340), .A2(new_n283), .B1(new_n313), .B2(new_n312), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT18), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n337), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n316), .A2(new_n322), .A3(new_n342), .A4(new_n345), .ZN(new_n346));
  OR2_X1    g0146(.A1(new_n346), .A2(KEYINPUT76), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(KEYINPUT76), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n274), .A2(G50), .B1(G20), .B2(new_n271), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n215), .A2(G33), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n204), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n329), .A2(new_n351), .A3(KEYINPUT74), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT74), .B1(new_n329), .B2(new_n351), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT11), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n329), .A2(new_n351), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT74), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT11), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n358), .A2(new_n352), .A3(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n252), .A2(new_n271), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT12), .B1(new_n260), .B2(G68), .ZN(new_n362));
  OR3_X1    g0162(.A1(new_n260), .A2(KEYINPUT12), .A3(G68), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n335), .A2(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n355), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  INV_X1    g0166(.A(new_n305), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n291), .A2(new_n306), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT68), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT68), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n291), .A2(new_n370), .A3(new_n306), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n367), .B1(new_n372), .B2(G238), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT13), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n324), .A2(G232), .A3(G1698), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G33), .A2(G97), .ZN(new_n376));
  INV_X1    g0176(.A(G1698), .ZN(new_n377));
  OAI211_X1 g0177(.A(G226), .B(new_n377), .C1(new_n263), .C2(new_n264), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n292), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n373), .A2(new_n374), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n374), .B1(new_n373), .B2(new_n380), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n366), .B(G169), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n371), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n370), .B1(new_n291), .B2(new_n306), .ZN(new_n385));
  OAI21_X1  g0185(.A(G238), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n380), .A2(new_n386), .A3(new_n305), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT13), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n373), .A2(new_n374), .A3(new_n380), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(G179), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n383), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n388), .A2(new_n389), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n366), .B1(new_n392), .B2(G169), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n365), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n355), .A2(new_n360), .A3(new_n364), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n388), .A2(G190), .A3(new_n389), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n381), .A2(new_n382), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n395), .B(new_n396), .C1(new_n397), .C2(new_n317), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n347), .A2(new_n348), .A3(new_n394), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n274), .A2(G150), .ZN(new_n400));
  OAI221_X1 g0200(.A(new_n400), .B1(new_n203), .B2(new_n215), .C1(new_n332), .C2(new_n350), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n329), .ZN(new_n402));
  INV_X1    g0202(.A(G50), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n252), .A2(new_n403), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n335), .A2(new_n404), .B1(new_n403), .B2(new_n334), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT9), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n402), .A2(KEYINPUT9), .A3(new_n405), .ZN(new_n409));
  AND2_X1   g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT10), .ZN(new_n411));
  OR2_X1    g0211(.A1(KEYINPUT3), .A2(G33), .ZN(new_n412));
  NAND2_X1  g0212(.A1(KEYINPUT3), .A2(G33), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n377), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n414), .A2(G223), .B1(new_n265), .B2(G77), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n324), .A2(G222), .A3(new_n377), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT69), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n291), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n418), .B2(new_n417), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n367), .B1(new_n372), .B2(G226), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(G190), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n421), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(G200), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n410), .A2(new_n411), .A3(new_n422), .A4(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n424), .A2(new_n408), .A3(new_n422), .A4(new_n409), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT10), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n423), .A2(G179), .ZN(new_n429));
  INV_X1    g0229(.A(new_n406), .ZN(new_n430));
  AOI21_X1  g0230(.A(G169), .B1(new_n420), .B2(new_n421), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n414), .A2(G238), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n324), .A2(G232), .A3(new_n377), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n434), .B(new_n435), .C1(new_n207), .C2(new_n324), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n292), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n372), .A2(G244), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n437), .A2(new_n305), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n313), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(new_n305), .A3(new_n438), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n283), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n252), .A2(new_n204), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n335), .A2(new_n443), .B1(new_n204), .B2(new_n334), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G20), .A2(G77), .ZN(new_n445));
  INV_X1    g0245(.A(new_n274), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT15), .B(G87), .ZN(new_n447));
  OAI221_X1 g0247(.A(new_n445), .B1(new_n250), .B2(new_n446), .C1(new_n350), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n329), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT72), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT72), .B1(new_n448), .B2(new_n329), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n444), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n440), .A2(new_n442), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n437), .A2(G190), .A3(new_n305), .A4(new_n438), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n456), .B(new_n444), .C1(new_n452), .C2(new_n451), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n439), .A2(new_n317), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n428), .A2(new_n433), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT73), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n461), .A2(new_n462), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n399), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n260), .A2(G116), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n467), .B(KEYINPUT84), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n259), .A2(G33), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n260), .B(new_n469), .C1(new_n256), .C2(new_n257), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n468), .B1(G116), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT85), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n206), .A2(KEYINPUT77), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT77), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G97), .ZN(new_n476));
  AOI21_X1  g0276(.A(G33), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G283), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n215), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n473), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n479), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT77), .B(G97), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n481), .B(KEYINPUT85), .C1(new_n482), .C2(G33), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n255), .A2(new_n214), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n215), .B2(G116), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT20), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n489), .B(new_n486), .C1(new_n480), .C2(new_n483), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n472), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n324), .A2(KEYINPUT82), .A3(G264), .A4(G1698), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(G1698), .B1(new_n412), .B2(new_n413), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(G257), .B1(new_n265), .B2(G303), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n496), .A2(KEYINPUT83), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT83), .B1(new_n496), .B2(new_n498), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n292), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n295), .A2(G1), .ZN(new_n502));
  XNOR2_X1  g0302(.A(KEYINPUT5), .B(G41), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n292), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G270), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n300), .A2(new_n502), .A3(new_n503), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n313), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n491), .A2(new_n501), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT21), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n283), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n491), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n496), .A2(new_n498), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT83), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n496), .A2(KEYINPUT83), .A3(new_n498), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n507), .B1(new_n517), .B2(new_n292), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n509), .B1(new_n512), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT86), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT86), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n509), .B(new_n521), .C1(new_n512), .C2(new_n518), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n491), .A2(G169), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n510), .B1(new_n523), .B2(new_n518), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n291), .B1(new_n515), .B2(new_n516), .ZN(new_n525));
  OAI21_X1  g0325(.A(G200), .B1(new_n525), .B2(new_n507), .ZN(new_n526));
  INV_X1    g0326(.A(new_n491), .ZN(new_n527));
  INV_X1    g0327(.A(G190), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n501), .A2(new_n505), .A3(new_n506), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n520), .A2(new_n522), .A3(new_n524), .A4(new_n530), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n291), .A2(G274), .A3(new_n502), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G116), .ZN(new_n533));
  INV_X1    g0333(.A(G244), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G1698), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(G238), .B2(G1698), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n533), .B1(new_n536), .B2(new_n265), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n532), .B1(new_n537), .B2(new_n292), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT78), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n295), .B2(G1), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n259), .A2(KEYINPUT78), .A3(G45), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n291), .A2(new_n540), .A3(G250), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT79), .ZN(new_n543));
  INV_X1    g0343(.A(G250), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n297), .B2(new_n290), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT79), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n541), .A4(new_n540), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n538), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G190), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT81), .ZN(new_n552));
  OR2_X1    g0352(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n553));
  NAND2_X1  g0353(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n376), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n552), .B1(new_n555), .B2(G20), .ZN(new_n556));
  INV_X1    g0356(.A(new_n376), .ZN(new_n557));
  AND2_X1   g0357(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n558));
  NOR2_X1   g0358(.A1(KEYINPUT80), .A2(KEYINPUT19), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(KEYINPUT81), .A3(new_n215), .ZN(new_n561));
  NOR2_X1   g0361(.A1(G87), .A2(G107), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n482), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n556), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n265), .A2(G20), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n474), .A2(new_n476), .ZN(new_n566));
  INV_X1    g0366(.A(new_n350), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n558), .A2(new_n559), .ZN(new_n569));
  AOI22_X1  g0369(.A1(G68), .A2(new_n565), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n329), .B1(new_n334), .B2(new_n447), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n549), .A2(G200), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n471), .A2(G87), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n551), .A2(new_n572), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n447), .A2(new_n334), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n470), .A2(new_n447), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n324), .A2(new_n215), .A3(G68), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n482), .A2(new_n350), .ZN(new_n579));
  INV_X1    g0379(.A(new_n569), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n560), .A2(new_n215), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n582), .A2(new_n552), .B1(new_n482), .B2(new_n562), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n581), .B1(new_n583), .B2(new_n561), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n576), .B(new_n577), .C1(new_n584), .C2(new_n258), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n549), .A2(new_n283), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n550), .A2(new_n313), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n575), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(G250), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n591));
  OAI211_X1 g0391(.A(G244), .B(new_n377), .C1(new_n263), .C2(new_n264), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT4), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n478), .B(new_n591), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(KEYINPUT4), .B1(new_n497), .B2(G244), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n292), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n503), .A2(new_n502), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n504), .A2(G257), .B1(new_n597), .B2(new_n300), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G200), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n260), .A2(G97), .ZN(new_n601));
  OAI21_X1  g0401(.A(G107), .B1(new_n266), .B2(new_n268), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n274), .A2(G77), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n207), .A2(KEYINPUT6), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n474), .B2(new_n476), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G97), .A2(G107), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT6), .B1(new_n208), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(G20), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n602), .A2(new_n603), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n601), .B1(new_n609), .B2(new_n329), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n471), .A2(G97), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n596), .A2(new_n598), .A3(G190), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n600), .A2(new_n610), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n215), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT22), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT22), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n324), .A2(new_n616), .A3(new_n215), .A4(G87), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT24), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n533), .A2(G20), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT23), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n215), .B2(G107), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g0424(.A1(new_n618), .A2(new_n619), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n619), .B1(new_n618), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n329), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n503), .A2(new_n502), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(G264), .A3(new_n291), .ZN(new_n629));
  NOR2_X1   g0429(.A1(G250), .A2(G1698), .ZN(new_n630));
  INV_X1    g0430(.A(G257), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n630), .B1(new_n631), .B2(G1698), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n632), .A2(new_n324), .B1(G33), .B2(G294), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n629), .B(new_n506), .C1(new_n633), .C2(new_n291), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n317), .ZN(new_n635));
  NAND2_X1  g0435(.A1(G33), .A2(G294), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n631), .A2(G1698), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(G250), .B2(G1698), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n638), .B2(new_n265), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n292), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n640), .A2(new_n528), .A3(new_n506), .A4(new_n629), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n334), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT87), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT25), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n260), .B2(G107), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n646), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n647), .A2(new_n648), .B1(G107), .B2(new_n471), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n627), .A2(new_n642), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n608), .A2(new_n603), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n207), .B1(new_n325), .B2(new_n326), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n329), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n601), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(new_n611), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n599), .A2(new_n283), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n596), .A2(new_n598), .A3(new_n313), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n613), .A2(new_n650), .A3(new_n658), .ZN(new_n659));
  OR3_X1    g0459(.A1(new_n634), .A2(KEYINPUT88), .A3(new_n313), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n634), .A2(new_n313), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT88), .B1(new_n634), .B2(G169), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n627), .A2(new_n649), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n590), .A2(new_n659), .A3(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n466), .A2(new_n531), .A3(new_n666), .ZN(G372));
  AND3_X1   g0467(.A1(new_n337), .A2(new_n343), .A3(new_n344), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n344), .B1(new_n337), .B2(new_n343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n394), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n455), .B2(new_n398), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n322), .A2(new_n342), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT90), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n674), .A2(new_n675), .B1(new_n427), .B2(new_n425), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n432), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n588), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n576), .B(new_n574), .C1(new_n584), .C2(new_n258), .ZN(new_n680));
  INV_X1    g0480(.A(new_n573), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT89), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT89), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n572), .A2(new_n683), .A3(new_n573), .A4(new_n574), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n682), .A2(new_n551), .A3(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n659), .A2(new_n588), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n529), .A2(new_n491), .A3(new_n511), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n524), .A2(new_n687), .A3(new_n509), .A4(new_n665), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n679), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n658), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n685), .A2(new_n588), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n590), .A2(KEYINPUT26), .A3(new_n690), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n678), .B1(new_n466), .B2(new_n697), .ZN(G369));
  NAND3_X1  g0498(.A1(new_n259), .A2(new_n215), .A3(G13), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G213), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G343), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n527), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n531), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT91), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n491), .A2(G169), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT21), .B1(new_n709), .B2(new_n529), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n706), .B1(new_n710), .B2(new_n519), .ZN(new_n711));
  AND3_X1   g0511(.A1(new_n707), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n708), .B1(new_n707), .B2(new_n711), .ZN(new_n713));
  OAI21_X1  g0513(.A(G330), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n665), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n704), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n664), .A2(new_n704), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n665), .A2(new_n650), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n714), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n710), .B1(KEYINPUT86), .B2(new_n519), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n704), .B1(new_n723), .B2(new_n522), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n650), .A3(new_n665), .A4(new_n717), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT92), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n665), .A2(new_n704), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n726), .B1(new_n725), .B2(new_n728), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n722), .B1(new_n729), .B2(new_n730), .ZN(G399));
  INV_X1    g0531(.A(new_n219), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G41), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G1), .ZN(new_n735));
  INV_X1    g0535(.A(G116), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n482), .A2(new_n736), .A3(new_n562), .ZN(new_n737));
  OAI22_X1  g0537(.A1(new_n735), .A2(new_n737), .B1(new_n212), .B2(new_n734), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT96), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n685), .A2(KEYINPUT26), .A3(new_n588), .A4(new_n690), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n692), .B1(new_n589), .B2(new_n658), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n520), .A2(new_n522), .A3(new_n524), .A4(new_n665), .ZN(new_n743));
  AOI221_X4 g0543(.A(new_n679), .B1(new_n741), .B2(new_n742), .C1(new_n743), .C2(new_n686), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n740), .B1(new_n744), .B2(new_n704), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n743), .A2(new_n686), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n741), .A2(new_n742), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n746), .A2(new_n588), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(KEYINPUT96), .A3(new_n705), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT29), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT29), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n696), .A2(KEYINPUT95), .A3(new_n705), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT95), .B1(new_n696), .B2(new_n705), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n599), .ZN(new_n758));
  AND4_X1   g0558(.A1(new_n548), .A2(new_n538), .A3(new_n629), .A4(new_n640), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n501), .A2(new_n508), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT30), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND3_X1   g0562(.A1(new_n596), .A2(new_n598), .A3(KEYINPUT30), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n501), .A2(new_n763), .A3(new_n508), .A4(new_n759), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n599), .A2(new_n313), .A3(new_n549), .A4(new_n634), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n762), .B(new_n764), .C1(new_n518), .C2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(KEYINPUT31), .B1(new_n766), .B2(new_n704), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT93), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n590), .A2(new_n659), .A3(new_n665), .A4(new_n705), .ZN(new_n769));
  OAI22_X1  g0569(.A1(new_n767), .A2(new_n768), .B1(new_n531), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n760), .A2(new_n761), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n764), .B1(new_n518), .B2(new_n765), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n704), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT31), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n766), .A2(KEYINPUT31), .A3(new_n704), .ZN(new_n776));
  AOI21_X1  g0576(.A(KEYINPUT93), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(G330), .B1(new_n770), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(KEYINPUT94), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT94), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n781), .B(G330), .C1(new_n770), .C2(new_n777), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n757), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n739), .B1(new_n786), .B2(G1), .ZN(G364));
  OR3_X1    g0587(.A1(new_n712), .A2(new_n713), .A3(G330), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n215), .A2(G13), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n259), .B1(new_n789), .B2(G45), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n733), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n788), .A2(new_n714), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n732), .A2(new_n265), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G355), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(G116), .B2(new_n219), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n245), .A2(new_n295), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n732), .A2(new_n324), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n295), .B2(new_n213), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n797), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G13), .A2(G33), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(G20), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT97), .Z(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n214), .B1(G20), .B2(new_n283), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n792), .B1(new_n802), .B2(new_n810), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT99), .B(G159), .Z(new_n812));
  NOR2_X1   g0612(.A1(new_n215), .A2(G179), .ZN(new_n813));
  NOR2_X1   g0613(.A1(G190), .A2(G200), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT32), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n528), .A2(G179), .A3(G200), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n215), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n816), .A2(new_n817), .B1(new_n206), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n816), .A2(new_n817), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n215), .A2(new_n313), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n822), .A2(G190), .A3(new_n317), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n814), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n821), .B1(new_n270), .B2(new_n823), .C1(new_n204), .C2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT98), .ZN(new_n826));
  INV_X1    g0626(.A(new_n822), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n827), .B2(new_n317), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n822), .A2(KEYINPUT98), .A3(G200), .ZN(new_n829));
  AND3_X1   g0629(.A1(new_n828), .A2(G190), .A3(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(new_n820), .B(new_n825), .C1(G50), .C2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n813), .A2(new_n528), .A3(G200), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G107), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n813), .A2(G190), .A3(G200), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G87), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n834), .A2(new_n837), .A3(new_n324), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT100), .Z(new_n839));
  NAND3_X1  g0639(.A1(new_n828), .A2(new_n528), .A3(new_n829), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n831), .B(new_n839), .C1(new_n271), .C2(new_n840), .ZN(new_n841));
  OR2_X1    g0641(.A1(new_n841), .A2(KEYINPUT101), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(KEYINPUT101), .ZN(new_n843));
  INV_X1    g0643(.A(G322), .ZN(new_n844));
  INV_X1    g0644(.A(G329), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n823), .A2(new_n844), .B1(new_n815), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n824), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n324), .B(new_n846), .C1(G311), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G283), .ZN(new_n849));
  INV_X1    g0649(.A(G303), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n849), .A2(new_n832), .B1(new_n835), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n819), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n851), .B1(G294), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n848), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n830), .ZN(new_n855));
  INV_X1    g0655(.A(G326), .ZN(new_n856));
  XNOR2_X1  g0656(.A(KEYINPUT102), .B(KEYINPUT33), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(G317), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n855), .A2(new_n856), .B1(new_n840), .B2(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n842), .B(new_n843), .C1(new_n854), .C2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n811), .B1(new_n860), .B2(new_n808), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n707), .A2(new_n711), .A3(new_n807), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n794), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G396));
  NAND2_X1  g0665(.A1(new_n460), .A2(new_n705), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n688), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n659), .A2(new_n588), .A3(new_n685), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n588), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR3_X1   g0670(.A1(new_n589), .A2(new_n692), .A3(new_n658), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n871), .B1(new_n692), .B2(new_n691), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n867), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OR2_X1    g0673(.A1(new_n754), .A2(new_n755), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n453), .A2(new_n704), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n454), .B1(new_n459), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n455), .A2(new_n705), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n874), .A2(KEYINPUT107), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT107), .B1(new_n874), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n873), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n792), .B1(new_n881), .B2(new_n784), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n784), .B2(new_n881), .ZN(new_n883));
  INV_X1    g0683(.A(new_n808), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n804), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n792), .B1(G77), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n833), .A2(G87), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n887), .B1(new_n207), .B2(new_n835), .C1(new_n206), .C2(new_n819), .ZN(new_n888));
  INV_X1    g0688(.A(new_n823), .ZN(new_n889));
  INV_X1    g0689(.A(new_n815), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n889), .A2(G294), .B1(new_n890), .B2(G311), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(new_n265), .C1(new_n736), .C2(new_n824), .ZN(new_n892));
  AOI211_X1 g0692(.A(new_n888), .B(new_n892), .C1(G303), .C2(new_n830), .ZN(new_n893));
  INV_X1    g0693(.A(new_n840), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n894), .A2(KEYINPUT103), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(KEYINPUT103), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n893), .B1(new_n849), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT104), .ZN(new_n900));
  INV_X1    g0700(.A(new_n812), .ZN(new_n901));
  AOI22_X1  g0701(.A1(G143), .A2(new_n889), .B1(new_n901), .B2(new_n847), .ZN(new_n902));
  INV_X1    g0702(.A(G150), .ZN(new_n903));
  INV_X1    g0703(.A(G137), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n902), .B1(new_n903), .B2(new_n840), .C1(new_n855), .C2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT34), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n906), .ZN(new_n908));
  INV_X1    g0708(.A(G132), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n324), .B1(new_n815), .B2(new_n909), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n403), .A2(new_n835), .B1(new_n832), .B2(new_n271), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n910), .B(new_n911), .C1(G58), .C2(new_n852), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n907), .A2(new_n908), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n900), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n886), .B1(new_n914), .B2(new_n808), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT105), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n803), .B2(new_n878), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT106), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n883), .A2(new_n919), .ZN(G384));
  OR2_X1    g0720(.A1(new_n605), .A2(new_n607), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n921), .A2(KEYINPUT35), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(KEYINPUT35), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n922), .A2(G116), .A3(new_n216), .A4(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT36), .Z(new_n925));
  OR3_X1    g0725(.A1(new_n212), .A2(new_n204), .A3(new_n272), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n403), .A2(G68), .ZN(new_n927));
  AOI211_X1 g0727(.A(new_n259), .B(G13), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n751), .A2(new_n756), .A3(new_n465), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n678), .ZN(new_n931));
  INV_X1    g0731(.A(new_n702), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n670), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT37), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n337), .A2(new_n932), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT110), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n337), .A2(new_n343), .ZN(new_n938));
  AOI21_X1  g0738(.A(G200), .B1(new_n338), .B2(new_n339), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n330), .B(new_n336), .C1(new_n939), .C2(new_n319), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n938), .A2(new_n935), .A3(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n937), .B(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n282), .A2(new_n702), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n346), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT38), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(KEYINPUT37), .B1(new_n943), .B2(KEYINPUT110), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n941), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n937), .A2(new_n938), .A3(new_n940), .A4(new_n935), .ZN(new_n948));
  AND4_X1   g0748(.A1(KEYINPUT38), .A2(new_n944), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT39), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n942), .A2(KEYINPUT38), .A3(new_n944), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n941), .A2(new_n934), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n938), .A2(new_n935), .A3(KEYINPUT37), .A4(new_n940), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT111), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n673), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n322), .A2(new_n342), .A3(KEYINPUT111), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n956), .A2(new_n670), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n954), .B1(new_n958), .B2(new_n943), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n951), .B1(new_n959), .B2(KEYINPUT38), .ZN(new_n960));
  XNOR2_X1  g0760(.A(KEYINPUT112), .B(KEYINPUT39), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n950), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n671), .A2(new_n705), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n933), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n945), .A2(new_n949), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n395), .A2(KEYINPUT109), .A3(new_n705), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT109), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n365), .B2(new_n704), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n394), .A2(new_n971), .A3(new_n398), .ZN(new_n972));
  OAI21_X1  g0772(.A(KEYINPUT14), .B1(new_n397), .B2(new_n283), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n398), .A2(new_n973), .A3(new_n390), .A4(new_n383), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n395), .A2(new_n705), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n866), .B1(new_n689), .B2(new_n695), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT108), .ZN(new_n979));
  INV_X1    g0779(.A(new_n877), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT108), .B1(new_n873), .B2(new_n877), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n967), .B(new_n977), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n966), .A2(new_n983), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n931), .B(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT38), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n670), .A2(new_n957), .ZN(new_n987));
  AOI21_X1  g0787(.A(KEYINPUT111), .B1(new_n322), .B2(new_n342), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n943), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n954), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n949), .B1(new_n986), .B2(new_n991), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n775), .B(new_n776), .C1(new_n531), .C2(new_n769), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n878), .B1(new_n972), .B2(new_n976), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n993), .A2(new_n994), .A3(KEYINPUT40), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT113), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n993), .A2(KEYINPUT40), .A3(new_n994), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT113), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n998), .A3(new_n960), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n993), .B(new_n994), .C1(new_n945), .C2(new_n949), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT40), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n465), .A2(new_n993), .ZN(new_n1005));
  OAI21_X1  g0805(.A(G330), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n985), .A2(new_n1007), .B1(new_n259), .B2(new_n789), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n985), .A2(new_n1007), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n929), .B1(new_n1008), .B2(new_n1009), .ZN(G367));
  NAND2_X1  g0810(.A1(new_n690), .A2(new_n704), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n655), .A2(new_n704), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n613), .A2(new_n658), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT114), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n722), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n680), .A2(new_n704), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n685), .A2(new_n588), .A3(new_n1018), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n588), .A2(new_n1018), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT43), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1021), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT43), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1014), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n725), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT42), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1015), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n690), .B1(new_n1029), .B2(new_n715), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT115), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n704), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1031), .B2(new_n1030), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1022), .B(new_n1025), .C1(new_n1028), .C2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1028), .A2(new_n1033), .A3(new_n1024), .A4(new_n1023), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  OR3_X1    g0836(.A1(new_n1017), .A2(new_n1034), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1017), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n733), .B(KEYINPUT41), .Z(new_n1040));
  OAI21_X1  g0840(.A(new_n1014), .B1(new_n729), .B2(new_n730), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT45), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g0843(.A(KEYINPUT45), .B(new_n1014), .C1(new_n729), .C2(new_n730), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n723), .A2(new_n522), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n705), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(new_n718), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT92), .B1(new_n1048), .B2(new_n727), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n725), .A2(new_n726), .A3(new_n728), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1049), .A2(new_n1050), .A3(new_n1026), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT44), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1049), .A2(KEYINPUT44), .A3(new_n1050), .A4(new_n1026), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n722), .B1(new_n1045), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n725), .B1(new_n724), .B2(new_n719), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n714), .A2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(G330), .C1(new_n712), .C2(new_n713), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n757), .A2(new_n1062), .A3(new_n784), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1045), .A2(new_n722), .A3(new_n1055), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1057), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1040), .B1(new_n1066), .B2(new_n786), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1039), .B1(new_n1067), .B2(new_n791), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n809), .B1(new_n219), .B2(new_n447), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n241), .A2(new_n800), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n792), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(G143), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n836), .A2(G58), .B1(new_n890), .B2(G137), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n855), .A2(new_n1072), .B1(new_n1073), .B2(KEYINPUT116), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1073), .A2(KEYINPUT116), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n324), .B1(new_n824), .B2(new_n403), .C1(new_n903), .C2(new_n823), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n819), .A2(new_n271), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n832), .A2(new_n204), .ZN(new_n1078));
  OR4_X1    g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1074), .B(new_n1079), .C1(new_n901), .C2(new_n897), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n823), .A2(new_n850), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n265), .B1(new_n824), .B2(new_n849), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(G317), .C2(new_n890), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n836), .A2(G116), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT46), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n830), .A2(G311), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n852), .A2(G107), .B1(new_n833), .B2(new_n566), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G294), .B2(new_n897), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1080), .A2(new_n1089), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT47), .Z(new_n1091));
  AOI21_X1  g0891(.A(new_n1071), .B1(new_n1091), .B2(new_n808), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n806), .B2(new_n1021), .ZN(new_n1093));
  XOR2_X1   g0893(.A(new_n1093), .B(KEYINPUT117), .Z(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1068), .A2(new_n1095), .ZN(G387));
  NAND3_X1  g0896(.A1(new_n785), .A2(new_n1061), .A3(new_n1060), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n733), .A3(new_n1063), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n265), .B1(new_n815), .B2(new_n856), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n852), .A2(G283), .B1(new_n836), .B2(G294), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n889), .A2(G317), .B1(new_n847), .B2(G303), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n855), .B2(new_n844), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n897), .B2(G311), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1100), .B1(new_n1103), .B2(KEYINPUT48), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(KEYINPUT48), .B2(new_n1103), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT49), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1099), .B(new_n1106), .C1(G116), .C2(new_n833), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n324), .B1(new_n824), .B2(new_n271), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G150), .B2(new_n890), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n836), .A2(G77), .B1(new_n833), .B2(G97), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(new_n332), .C2(new_n840), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n819), .A2(new_n447), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G50), .B2(new_n889), .ZN(new_n1113));
  XOR2_X1   g0913(.A(new_n1113), .B(KEYINPUT119), .Z(new_n1114));
  AOI211_X1 g0914(.A(new_n1111), .B(new_n1114), .C1(G159), .C2(new_n830), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n808), .B1(new_n1107), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n719), .A2(new_n806), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n795), .A2(new_n737), .B1(new_n207), .B2(new_n732), .ZN(new_n1118));
  AOI211_X1 g0918(.A(G45), .B(new_n737), .C1(G68), .C2(G77), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n250), .A2(G50), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(KEYINPUT50), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1120), .A2(KEYINPUT50), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1119), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n799), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n238), .A2(new_n295), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1118), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1126), .A2(KEYINPUT118), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n810), .B1(new_n1126), .B2(KEYINPUT118), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n793), .B(new_n1117), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1062), .A2(new_n791), .B1(new_n1116), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT120), .B1(new_n1098), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1098), .A2(KEYINPUT120), .A3(new_n1130), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(G393));
  AND3_X1   g0934(.A1(new_n1045), .A2(new_n722), .A3(new_n1055), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1063), .B1(new_n1135), .B2(new_n1056), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1066), .A2(new_n1136), .A3(new_n733), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1015), .A2(new_n807), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT121), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n248), .A2(new_n800), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n809), .B1(new_n219), .B2(new_n482), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n830), .A2(G317), .B1(G311), .B2(new_n889), .ZN(new_n1142));
  XOR2_X1   g0942(.A(new_n1142), .B(KEYINPUT52), .Z(new_n1143));
  INV_X1    g0943(.A(G294), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n265), .B1(new_n815), .B2(new_n844), .C1(new_n1144), .C2(new_n824), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n834), .B1(new_n849), .B2(new_n835), .C1(new_n736), .C2(new_n819), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1145), .B(new_n1146), .C1(new_n897), .C2(G303), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n324), .B1(new_n815), .B2(new_n1072), .C1(new_n250), .C2(new_n824), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n887), .B1(new_n271), .B2(new_n835), .C1(new_n204), .C2(new_n819), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(new_n897), .C2(G50), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n830), .A2(G150), .B1(G159), .B2(new_n889), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(KEYINPUT122), .B(KEYINPUT51), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1143), .A2(new_n1147), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n792), .B1(new_n1140), .B2(new_n1141), .C1(new_n1154), .C2(new_n884), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1139), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1135), .A2(new_n1056), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n791), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1137), .A2(new_n1158), .ZN(G390));
  NAND3_X1  g0959(.A1(new_n745), .A2(new_n749), .A3(new_n877), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n876), .A3(new_n977), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n992), .A2(new_n965), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n963), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n977), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n979), .B1(new_n978), .B2(new_n980), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n873), .A2(KEYINPUT108), .A3(new_n877), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1164), .B1(new_n1168), .B2(new_n965), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n878), .B1(new_n779), .B2(new_n782), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n977), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1163), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n993), .A2(G330), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n994), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n1163), .B2(new_n1169), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n791), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n792), .B1(new_n251), .B2(new_n885), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n898), .A2(new_n207), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n837), .B1(new_n271), .B2(new_n832), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G77), .B2(new_n852), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n824), .A2(new_n482), .B1(new_n815), .B2(new_n1144), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n324), .B(new_n1182), .C1(G116), .C2(new_n889), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1181), .B(new_n1183), .C1(new_n849), .C2(new_n855), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n898), .A2(new_n904), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n830), .A2(G128), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n835), .A2(new_n903), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n1187), .B(KEYINPUT53), .ZN(new_n1188));
  INV_X1    g0988(.A(G125), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n823), .A2(new_n909), .B1(new_n815), .B2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT54), .B(G143), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n324), .B1(new_n824), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n852), .A2(G159), .B1(new_n833), .B2(G50), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1186), .A2(new_n1188), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n1179), .A2(new_n1184), .B1(new_n1185), .B2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1178), .B1(new_n1196), .B2(new_n808), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n963), .B2(new_n804), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1177), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1174), .B1(new_n1170), .B2(new_n977), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1173), .A2(new_n877), .A3(new_n876), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n1160), .A2(new_n876), .B1(new_n1165), .B2(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1200), .A2(new_n1201), .B1(new_n1203), .B2(new_n1171), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n465), .A2(new_n1173), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n930), .A2(new_n678), .A3(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT123), .B1(new_n1176), .B2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1163), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1163), .A2(new_n1169), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1209), .B1(new_n1210), .B2(new_n1174), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1203), .A2(new_n1171), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AND3_X1   g1014(.A1(new_n930), .A2(new_n678), .A3(new_n1205), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT123), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1211), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1208), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n734), .B1(new_n1176), .B2(new_n1207), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1199), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(G378));
  INV_X1    g1022(.A(KEYINPUT124), .ZN(new_n1223));
  INV_X1    g1023(.A(G330), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n428), .A2(new_n433), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n430), .A2(new_n702), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1227), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n428), .A2(new_n433), .A3(new_n1229), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1228), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1231), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1229), .B1(new_n428), .B2(new_n433), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n432), .B(new_n1227), .C1(new_n425), .C2(new_n427), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1232), .A2(new_n1236), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n992), .A2(KEYINPUT113), .A3(new_n995), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n998), .B1(new_n997), .B2(new_n960), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1225), .B(new_n1237), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1237), .B1(new_n1000), .B2(new_n1225), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n984), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1225), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1237), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n966), .A2(new_n983), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1246), .A2(new_n1247), .A3(new_n1240), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1223), .B1(new_n1243), .B2(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT124), .B1(new_n1250), .B2(new_n1247), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1206), .B1(new_n1176), .B2(new_n1207), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n733), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(KEYINPUT125), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT125), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1256), .B(new_n733), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1215), .B1(new_n1211), .B2(new_n1216), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1243), .A2(new_n1248), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT57), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1255), .A2(new_n1257), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n791), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n792), .B1(G50), .B2(new_n885), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n403), .B1(G33), .B2(G41), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n265), .B2(new_n294), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1077), .B1(G77), .B2(new_n836), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n270), .B2(new_n832), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n294), .B(new_n265), .C1(new_n823), .C2(new_n207), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n824), .A2(new_n447), .B1(new_n815), .B2(new_n849), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1271), .B1(new_n206), .B2(new_n840), .C1(new_n736), .C2(new_n855), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT58), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1266), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n835), .A2(new_n1191), .ZN(new_n1275));
  INV_X1    g1075(.A(G128), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n823), .A2(new_n1276), .B1(new_n824), .B2(new_n904), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n1275), .B(new_n1277), .C1(G150), .C2(new_n852), .ZN(new_n1278));
  OAI221_X1 g1078(.A(new_n1278), .B1(new_n1189), .B2(new_n855), .C1(new_n909), .C2(new_n840), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(KEYINPUT59), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(KEYINPUT59), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n901), .A2(new_n833), .ZN(new_n1282));
  AOI211_X1 g1082(.A(G33), .B(G41), .C1(new_n890), .C2(G124), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  OAI221_X1 g1084(.A(new_n1274), .B1(new_n1273), .B2(new_n1272), .C1(new_n1280), .C2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1264), .B1(new_n1285), .B2(new_n808), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n1245), .B2(new_n804), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1263), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1262), .A2(new_n1289), .ZN(G375));
  INV_X1    g1090(.A(new_n1040), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1216), .A2(new_n1291), .A3(new_n1292), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n792), .B1(G68), .B2(new_n885), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n898), .A2(new_n1191), .ZN(new_n1295));
  OAI22_X1  g1095(.A1(new_n823), .A2(new_n904), .B1(new_n824), .B2(new_n903), .ZN(new_n1296));
  AOI211_X1 g1096(.A(new_n265), .B(new_n1296), .C1(G128), .C2(new_n890), .ZN(new_n1297));
  INV_X1    g1097(.A(G159), .ZN(new_n1298));
  OAI22_X1  g1098(.A1(new_n270), .A2(new_n832), .B1(new_n835), .B2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(G50), .B2(new_n852), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1297), .B(new_n1300), .C1(new_n909), .C2(new_n855), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n898), .A2(new_n736), .ZN(new_n1302));
  OAI22_X1  g1102(.A1(new_n824), .A2(new_n207), .B1(new_n815), .B2(new_n850), .ZN(new_n1303));
  AOI211_X1 g1103(.A(new_n324), .B(new_n1303), .C1(G283), .C2(new_n889), .ZN(new_n1304));
  AOI211_X1 g1104(.A(new_n1078), .B(new_n1112), .C1(G97), .C2(new_n836), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1304), .B(new_n1305), .C1(new_n1144), .C2(new_n855), .ZN(new_n1306));
  OAI22_X1  g1106(.A1(new_n1295), .A2(new_n1301), .B1(new_n1302), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1294), .B1(new_n1307), .B2(new_n808), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1308), .B1(new_n977), .B2(new_n804), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1309), .B1(new_n1204), .B2(new_n790), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1293), .A2(new_n1311), .ZN(G381));
  NOR3_X1   g1112(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1313), .A2(new_n1095), .A3(new_n1068), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1260), .B1(new_n1254), .B2(KEYINPUT125), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1288), .B1(new_n1315), .B2(new_n1257), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1133), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1317), .A2(G396), .A3(new_n1131), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1314), .A2(new_n1316), .A3(new_n1221), .A4(new_n1318), .ZN(G407));
  NAND2_X1  g1119(.A1(new_n703), .A2(G213), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1316), .A2(new_n1221), .A3(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(G407), .A2(G213), .A3(new_n1322), .ZN(G409));
  NAND2_X1  g1123(.A1(new_n1292), .A2(KEYINPUT126), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT60), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1292), .A2(KEYINPUT126), .A3(KEYINPUT60), .ZN(new_n1327));
  AND2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1216), .A2(new_n733), .ZN(new_n1329));
  OAI211_X1 g1129(.A(G384), .B(new_n1311), .C1(new_n1328), .C2(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1329), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n919), .B(new_n883), .C1(new_n1331), .C2(new_n1310), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  AOI211_X1 g1134(.A(new_n1221), .B(new_n1288), .C1(new_n1315), .C2(new_n1257), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1258), .A2(new_n1291), .A3(new_n1259), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n791), .B1(new_n1249), .B2(new_n1251), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1336), .A2(new_n1287), .A3(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(new_n1221), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1320), .B(new_n1334), .C1(new_n1335), .C2(new_n1340), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(KEYINPUT62), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT61), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1262), .A2(G378), .A3(new_n1289), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1321), .B1(new_n1344), .B2(new_n1339), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT62), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1345), .A2(new_n1346), .A3(new_n1334), .ZN(new_n1347));
  INV_X1    g1147(.A(G2897), .ZN(new_n1348));
  OAI211_X1 g1148(.A(new_n1330), .B(new_n1332), .C1(new_n1348), .C2(new_n1320), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1320), .A2(new_n1348), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1333), .A2(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1340), .B1(new_n1316), .B2(G378), .ZN(new_n1352));
  OAI211_X1 g1152(.A(new_n1349), .B(new_n1351), .C1(new_n1352), .C2(new_n1321), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1342), .A2(new_n1343), .A3(new_n1347), .A4(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(G390), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1356));
  NOR3_X1   g1156(.A1(new_n1135), .A2(new_n1056), .A3(new_n1063), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1291), .B1(new_n1357), .B2(new_n785), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n1356), .B1(new_n1358), .B2(new_n790), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1355), .B1(new_n1359), .B2(new_n1094), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n864), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1361));
  NOR2_X1   g1161(.A1(new_n1361), .A2(new_n1318), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1068), .A2(new_n1095), .A3(G390), .ZN(new_n1363));
  AND3_X1   g1163(.A1(new_n1360), .A2(new_n1362), .A3(new_n1363), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1362), .B1(new_n1360), .B2(new_n1363), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(new_n1364), .A2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1366), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1354), .A2(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1351), .A2(new_n1349), .ZN(new_n1369));
  OAI211_X1 g1169(.A(new_n1366), .B(new_n1343), .C1(new_n1345), .C2(new_n1369), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1370), .ZN(new_n1371));
  INV_X1    g1171(.A(KEYINPUT127), .ZN(new_n1372));
  AOI211_X1 g1172(.A(new_n1321), .B(new_n1333), .C1(new_n1344), .C2(new_n1339), .ZN(new_n1373));
  OAI21_X1  g1173(.A(new_n1372), .B1(new_n1373), .B2(KEYINPUT63), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1373), .A2(KEYINPUT63), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT63), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1341), .A2(KEYINPUT127), .A3(new_n1376), .ZN(new_n1377));
  NAND4_X1  g1177(.A1(new_n1371), .A2(new_n1374), .A3(new_n1375), .A4(new_n1377), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1368), .A2(new_n1378), .ZN(G405));
  NAND2_X1  g1179(.A1(G375), .A2(new_n1221), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1380), .A2(new_n1344), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1381), .A2(new_n1334), .ZN(new_n1382));
  NAND3_X1  g1182(.A1(new_n1380), .A2(new_n1344), .A3(new_n1333), .ZN(new_n1383));
  NAND2_X1  g1183(.A1(new_n1382), .A2(new_n1383), .ZN(new_n1384));
  XNOR2_X1  g1184(.A(new_n1384), .B(new_n1367), .ZN(G402));
endmodule


