//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n735, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971;
  NAND2_X1  g000(.A1(G29gat), .A2(G36gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g003(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G43gat), .ZN(new_n208));
  INV_X1    g007(.A(G43gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G50gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT15), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT15), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n209), .A2(G50gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n207), .A2(G43gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(new_n202), .A3(new_n211), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT14), .ZN(new_n219));
  INV_X1    g018(.A(G29gat), .ZN(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT86), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n205), .A2(KEYINPUT86), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n204), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n213), .B1(new_n218), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT87), .ZN(new_n228));
  INV_X1    g027(.A(G22gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G15gat), .ZN(new_n230));
  INV_X1    g029(.A(G15gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G22gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT88), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G1gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n230), .A2(new_n232), .A3(new_n233), .A4(G1gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT16), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n230), .A2(new_n232), .A3(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G8gat), .ZN(new_n241));
  INV_X1    g040(.A(G8gat), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n236), .A2(new_n242), .A3(new_n237), .A4(new_n239), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT87), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n245), .B(new_n213), .C1(new_n218), .C2(new_n226), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT89), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n228), .A2(new_n244), .A3(KEYINPUT89), .A4(new_n246), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(KEYINPUT17), .B(new_n213), .C1(new_n218), .C2(new_n226), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(new_n244), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT17), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n228), .A2(new_n255), .A3(new_n246), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n254), .A2(new_n256), .B1(G229gat), .B2(G233gat), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n251), .A2(new_n257), .A3(KEYINPUT18), .ZN(new_n258));
  XNOR2_X1  g057(.A(G113gat), .B(G141gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(G197gat), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT11), .B(G169gat), .Z(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT12), .ZN(new_n263));
  INV_X1    g062(.A(new_n244), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n228), .A2(new_n246), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n249), .A2(new_n250), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G229gat), .A2(G233gat), .ZN(new_n267));
  XOR2_X1   g066(.A(new_n267), .B(KEYINPUT13), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n258), .B(new_n263), .C1(new_n266), .C2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(KEYINPUT18), .B1(new_n251), .B2(new_n257), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT90), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI211_X1 g072(.A(KEYINPUT90), .B(KEYINPUT18), .C1(new_n251), .C2(new_n257), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n270), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n251), .A2(KEYINPUT18), .A3(new_n257), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n265), .A2(new_n264), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n269), .B1(new_n251), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n271), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n263), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G78gat), .B(G106gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G22gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G228gat), .ZN(new_n286));
  INV_X1    g085(.A(G233gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT22), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n290), .A2(KEYINPUT76), .B1(G211gat), .B2(G218gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(KEYINPUT76), .B2(new_n290), .ZN(new_n292));
  XNOR2_X1  g091(.A(G197gat), .B(G204gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT77), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G211gat), .B(G218gat), .Z(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n294), .B(KEYINPUT77), .ZN(new_n299));
  INV_X1    g098(.A(new_n297), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(KEYINPUT78), .B(KEYINPUT29), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  INV_X1    g104(.A(G155gat), .ZN(new_n306));
  INV_X1    g105(.A(G162gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G141gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(G148gat), .ZN(new_n310));
  INV_X1    g109(.A(G148gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(G141gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n305), .B(new_n308), .C1(new_n313), .C2(KEYINPUT2), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n305), .B1(new_n308), .B2(KEYINPUT2), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT79), .B1(new_n309), .B2(G148gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n316), .B1(G141gat), .B2(new_n311), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n309), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n304), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n289), .B1(new_n302), .B2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT3), .B1(new_n302), .B2(new_n303), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n324), .B1(new_n326), .B2(new_n320), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT29), .B1(new_n298), .B2(new_n301), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n320), .B1(new_n328), .B2(KEYINPUT3), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n302), .A2(new_n323), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n289), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT31), .B(G50gat), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n327), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n333), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n302), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n321), .B1(new_n337), .B2(new_n322), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n288), .B1(new_n338), .B2(new_n330), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n331), .B(new_n289), .C1(new_n321), .C2(new_n325), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n335), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n285), .B1(new_n334), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n333), .B1(new_n327), .B2(new_n332), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n339), .A2(new_n340), .A3(new_n335), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(new_n344), .A3(new_n284), .ZN(new_n345));
  INV_X1    g144(.A(G227gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(new_n287), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT25), .ZN(new_n349));
  XOR2_X1   g148(.A(KEYINPUT66), .B(G190gat), .Z(new_n350));
  INV_X1    g149(.A(G183gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n349), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n358), .A2(KEYINPUT23), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n358), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  OAI221_X1 g162(.A(new_n355), .B1(G183gat), .B2(G190gat), .C1(new_n353), .C2(KEYINPUT64), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n353), .A2(KEYINPUT64), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT25), .B1(new_n366), .B2(new_n361), .ZN(new_n367));
  XOR2_X1   g166(.A(KEYINPUT27), .B(G183gat), .Z(new_n368));
  INV_X1    g167(.A(KEYINPUT28), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT66), .B(G190gat), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT67), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT27), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(G183gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT27), .B(G183gat), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n350), .B(new_n374), .C1(new_n372), .C2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n371), .B1(new_n369), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(G169gat), .B2(G176gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n380), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT68), .ZN(new_n383));
  OAI22_X1  g182(.A1(new_n363), .A2(new_n367), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G113gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT69), .B(G120gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT70), .B(G113gat), .ZN(new_n387));
  INV_X1    g186(.A(G120gat), .ZN(new_n388));
  OAI22_X1  g187(.A1(new_n385), .A2(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G127gat), .B(G134gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT71), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT71), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT1), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n389), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n385), .A2(new_n388), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT1), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(G113gat), .B2(G120gat), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n391), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n395), .A2(new_n399), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n383), .A2(new_n377), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n361), .B1(new_n365), .B2(new_n364), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n349), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n362), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n402), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n348), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT74), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT34), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n384), .A2(new_n400), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n403), .A2(new_n402), .A3(new_n406), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n347), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n410), .A2(new_n411), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G71gat), .B(G99gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT72), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(G15gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(G43gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n413), .A2(new_n347), .A3(new_n414), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(KEYINPUT32), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n421), .B(KEYINPUT32), .C1(new_n422), .C2(new_n420), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n408), .A2(KEYINPUT74), .A3(new_n409), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n416), .A2(new_n425), .A3(new_n426), .A4(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n425), .A2(new_n426), .ZN(new_n429));
  INV_X1    g228(.A(new_n409), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n411), .B1(new_n415), .B2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n427), .B(new_n431), .C1(KEYINPUT34), .C2(new_n408), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n342), .A2(new_n345), .A3(new_n428), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(G226gat), .A2(G233gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n383), .A2(new_n377), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n404), .A2(new_n349), .B1(new_n357), .B2(new_n361), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n435), .B1(new_n438), .B2(KEYINPUT29), .ZN(new_n439));
  INV_X1    g238(.A(new_n435), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n384), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(new_n441), .A3(new_n302), .ZN(new_n442));
  INV_X1    g241(.A(new_n302), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n440), .B1(new_n384), .B2(new_n303), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n435), .B1(new_n403), .B2(new_n406), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G8gat), .B(G36gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(G64gat), .B(G92gat), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n448), .B(new_n449), .Z(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n442), .A2(new_n446), .A3(new_n450), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(KEYINPUT30), .A3(new_n453), .ZN(new_n454));
  OR3_X1    g253(.A1(new_n447), .A2(KEYINPUT30), .A3(new_n451), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n434), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g257(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n459));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n400), .A2(new_n460), .A3(new_n321), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT80), .B1(new_n402), .B2(new_n320), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n402), .A2(new_n320), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(G225gat), .A2(G233gat), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n459), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT4), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n461), .A2(new_n468), .A3(new_n462), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n321), .A2(new_n322), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n320), .A2(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n402), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n402), .A2(new_n320), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT4), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n469), .A2(new_n465), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n467), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n461), .A2(KEYINPUT4), .A3(new_n462), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT82), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n473), .A2(new_n478), .A3(new_n468), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n400), .A2(new_n468), .A3(new_n321), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT82), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n472), .A2(new_n465), .A3(new_n459), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n476), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n486));
  XNOR2_X1  g285(.A(G1gat), .B(G29gat), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT0), .ZN(new_n488));
  XNOR2_X1  g287(.A(G57gat), .B(G85gat), .ZN(new_n489));
  XOR2_X1   g288(.A(new_n488), .B(new_n489), .Z(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n485), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n475), .A2(new_n467), .B1(new_n482), .B2(new_n483), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT85), .B1(new_n493), .B2(new_n490), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT6), .B1(new_n493), .B2(new_n490), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n485), .A2(KEYINPUT6), .A3(new_n491), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT35), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n458), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n485), .B2(new_n491), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n493), .A2(new_n490), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n503), .A2(new_n456), .A3(KEYINPUT83), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT83), .B1(new_n503), .B2(new_n456), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n504), .A2(new_n505), .A3(new_n434), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT35), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n499), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND4_X1   g307(.A1(new_n455), .A2(new_n454), .A3(new_n492), .A4(new_n494), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n461), .A2(new_n462), .A3(new_n465), .A4(new_n463), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT84), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n482), .A2(new_n472), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT39), .B(new_n511), .C1(new_n512), .C2(new_n465), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n465), .B1(new_n482), .B2(new_n472), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT39), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n491), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n513), .A2(KEYINPUT40), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT40), .B1(new_n513), .B2(new_n516), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n509), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n451), .B1(new_n447), .B2(KEYINPUT37), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT37), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n440), .B1(new_n384), .B2(new_n336), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n524), .A2(new_n445), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n523), .B1(new_n525), .B2(new_n443), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n302), .B1(new_n444), .B2(new_n445), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT38), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n447), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n522), .A2(new_n528), .B1(new_n529), .B2(new_n450), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n523), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT38), .B1(new_n531), .B2(new_n521), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n530), .A2(new_n497), .A3(new_n496), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n342), .A2(new_n345), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n534), .B1(new_n504), .B2(new_n505), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT75), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT36), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(KEYINPUT75), .A2(KEYINPUT36), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n429), .A2(new_n432), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n416), .A2(new_n427), .B1(new_n425), .B2(new_n426), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n540), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n428), .A2(new_n433), .A3(new_n538), .A4(new_n539), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n536), .A2(new_n537), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n282), .B1(new_n508), .B2(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G57gat), .B(G64gat), .Z(new_n550));
  OR2_X1    g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(G71gat), .A2(G78gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT9), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n552), .B(new_n551), .C1(new_n557), .C2(new_n554), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G231gat), .A2(G233gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n564), .B(KEYINPUT91), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n563), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G127gat), .B(G155gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n566), .A2(new_n567), .ZN(new_n570));
  XOR2_X1   g369(.A(G183gat), .B(G211gat), .Z(new_n571));
  NOR3_X1   g370(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n264), .B1(new_n560), .B2(new_n559), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n574), .B(new_n575), .Z(new_n576));
  OAI21_X1  g375(.A(new_n571), .B1(new_n569), .B2(new_n570), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n576), .ZN(new_n579));
  INV_X1    g378(.A(new_n571), .ZN(new_n580));
  INV_X1    g379(.A(new_n570), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(new_n568), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n579), .B1(new_n582), .B2(new_n572), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585));
  INV_X1    g384(.A(G85gat), .ZN(new_n586));
  INV_X1    g385(.A(G92gat), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n585), .B(KEYINPUT7), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT7), .ZN(new_n589));
  OAI211_X1 g388(.A(G85gat), .B(G92gat), .C1(new_n589), .C2(KEYINPUT94), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G99gat), .B(G106gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n593), .B1(new_n586), .B2(new_n587), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n592), .B1(new_n591), .B2(new_n594), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n228), .A2(new_n246), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n597), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n256), .A2(new_n252), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT95), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G134gat), .B(G162gat), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n605), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n600), .A2(new_n610), .A3(new_n602), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n606), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n609), .B1(new_n606), .B2(new_n611), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n591), .A2(new_n594), .ZN(new_n615));
  INV_X1    g414(.A(new_n592), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n617), .A2(new_n558), .A3(new_n556), .A4(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n559), .B1(new_n595), .B2(new_n596), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n558), .A4(new_n556), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n619), .B2(new_n620), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n627), .A2(KEYINPUT96), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n619), .A2(new_n620), .ZN(new_n629));
  INV_X1    g428(.A(new_n625), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(KEYINPUT96), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n626), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n633), .B(new_n634), .Z(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n632), .B(new_n636), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n584), .A2(new_n614), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n549), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(new_n503), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT97), .B(G1gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(G1324gat));
  NAND3_X1  g441(.A1(new_n549), .A2(new_n457), .A3(new_n638), .ZN(new_n643));
  XNOR2_X1  g442(.A(KEYINPUT16), .B(G8gat), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n645), .A2(new_n646), .A3(KEYINPUT42), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT42), .B1(new_n645), .B2(new_n646), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n643), .A2(G8gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(KEYINPUT99), .ZN(new_n650));
  AND2_X1   g449(.A1(new_n649), .A2(KEYINPUT99), .ZN(new_n651));
  OAI22_X1  g450(.A1(new_n647), .A2(new_n648), .B1(new_n650), .B2(new_n651), .ZN(G1325gat));
  OR2_X1    g451(.A1(new_n547), .A2(KEYINPUT100), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n547), .A2(KEYINPUT100), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(G15gat), .B1(new_n639), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n428), .A2(new_n433), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n231), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n656), .B1(new_n639), .B2(new_n659), .ZN(G1326gat));
  NOR2_X1   g459(.A1(new_n639), .A2(new_n535), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT43), .B(G22gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  INV_X1    g462(.A(new_n637), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n549), .A2(new_n584), .A3(new_n614), .A4(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(G29gat), .A3(new_n503), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT45), .Z(new_n667));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n508), .A2(new_n548), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n668), .B1(new_n669), .B2(new_n614), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n614), .A2(KEYINPUT103), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(new_n612), .B2(new_n613), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n668), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n537), .A2(KEYINPUT102), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n534), .B1(new_n509), .B2(new_n519), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n546), .B1(new_n677), .B2(new_n533), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n679), .B(new_n534), .C1(new_n504), .C2(new_n505), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n676), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n675), .B1(new_n681), .B2(new_n508), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n670), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n584), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n275), .B2(new_n281), .ZN(new_n686));
  INV_X1    g485(.A(new_n263), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n258), .B1(new_n266), .B2(new_n269), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(new_n271), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n271), .B(new_n272), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n689), .B(KEYINPUT101), .C1(new_n690), .C2(new_n270), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n684), .A2(new_n692), .A3(new_n637), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n683), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n503), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n667), .B1(new_n697), .B2(new_n220), .ZN(G1328gat));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n221), .B1(new_n699), .B2(KEYINPUT104), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n665), .A2(new_n456), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(KEYINPUT104), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n683), .A2(new_n693), .ZN(new_n704));
  OAI21_X1  g503(.A(G36gat), .B1(new_n704), .B2(new_n456), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(G1329gat));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707));
  INV_X1    g506(.A(new_n655), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n209), .B1(new_n694), .B2(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n665), .A2(G43gat), .A3(new_n657), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n710), .A2(KEYINPUT105), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n707), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(KEYINPUT47), .B(G43gat), .C1(new_n704), .C2(new_n547), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n710), .B1(KEYINPUT105), .B2(new_n707), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(G1330gat));
  NOR3_X1   g515(.A1(new_n665), .A2(G50gat), .A3(new_n535), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n683), .A2(new_n534), .A3(new_n693), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(G50gat), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1331gat));
  INV_X1    g520(.A(new_n614), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n684), .A2(new_n692), .A3(new_n722), .A4(new_n637), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(new_n681), .B2(new_n508), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n695), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n457), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n727), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT49), .B(G64gat), .Z(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(G1333gat));
  NAND2_X1  g529(.A1(new_n724), .A2(new_n708), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n657), .A2(G71gat), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n731), .A2(G71gat), .B1(new_n724), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g533(.A1(new_n724), .A2(new_n534), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g535(.A1(new_n681), .A2(new_n508), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n738));
  INV_X1    g537(.A(new_n692), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n684), .A2(new_n739), .A3(new_n722), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n737), .A2(new_n738), .A3(KEYINPUT51), .A4(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n740), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n742), .B1(new_n681), .B2(new_n508), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(KEYINPUT51), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n738), .B1(new_n743), .B2(KEYINPUT51), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n746), .A2(new_n586), .A3(new_n695), .A4(new_n637), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n684), .A2(new_n739), .A3(new_n664), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n683), .A2(new_n695), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n747), .B1(new_n750), .B2(new_n586), .ZN(G1336gat));
  NOR3_X1   g550(.A1(new_n456), .A2(G92gat), .A3(new_n664), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n752), .B1(new_n744), .B2(new_n745), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n457), .B(new_n748), .C1(new_n670), .C2(new_n682), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT52), .B1(new_n754), .B2(G92gat), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(G92gat), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n743), .A2(KEYINPUT51), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n743), .A2(KEYINPUT51), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n752), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n757), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(KEYINPUT108), .B1(new_n756), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n753), .A2(new_n755), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n758), .A2(new_n761), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n764), .B(new_n765), .C1(new_n766), .C2(new_n757), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(new_n767), .ZN(G1337gat));
  NOR3_X1   g567(.A1(new_n657), .A2(G99gat), .A3(new_n664), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n746), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n683), .A2(new_n748), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT109), .B1(new_n771), .B2(new_n655), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G99gat), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n771), .A2(KEYINPUT109), .A3(new_n655), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n770), .B1(new_n773), .B2(new_n774), .ZN(G1338gat));
  NOR3_X1   g574(.A1(new_n535), .A2(G106gat), .A3(new_n664), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n744), .B2(new_n745), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT53), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n534), .B(new_n748), .C1(new_n670), .C2(new_n682), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT110), .B(G106gat), .Z(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n777), .A2(new_n778), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n777), .A2(KEYINPUT111), .A3(new_n778), .A4(new_n781), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n776), .B1(new_n759), .B2(new_n760), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n781), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n784), .B(new_n785), .C1(new_n778), .C2(new_n787), .ZN(G1339gat));
  NOR2_X1   g587(.A1(new_n626), .A2(KEYINPUT54), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n789), .A2(new_n635), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n624), .B2(new_n625), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n622), .A2(new_n623), .A3(new_n630), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n793), .B1(new_n792), .B2(new_n794), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n790), .B(KEYINPUT55), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n632), .A2(new_n636), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n626), .A2(KEYINPUT54), .A3(new_n794), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT112), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT55), .B1(new_n803), .B2(new_n790), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n686), .A2(new_n691), .A3(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n275), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n266), .A2(new_n269), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n254), .A2(new_n256), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n267), .B1(new_n251), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n262), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n637), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n674), .B1(new_n806), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n671), .A2(new_n673), .ZN(new_n814));
  OR2_X1    g613(.A1(new_n799), .A2(new_n804), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n807), .A2(new_n811), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n584), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n638), .A2(new_n692), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n503), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n458), .ZN(new_n821));
  OR3_X1    g620(.A1(new_n821), .A2(new_n387), .A3(new_n692), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n457), .A2(new_n657), .A3(new_n503), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n818), .A2(new_n819), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT113), .B1(new_n824), .B2(new_n535), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n826));
  AOI211_X1 g625(.A(new_n826), .B(new_n534), .C1(new_n818), .C2(new_n819), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n823), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(KEYINPUT114), .ZN(new_n829));
  INV_X1    g628(.A(new_n282), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n831), .B(new_n823), .C1(new_n825), .C2(new_n827), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n822), .B1(new_n833), .B2(new_n385), .ZN(G1340gat));
  OR3_X1    g633(.A1(new_n821), .A2(new_n386), .A3(new_n664), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n829), .A2(new_n637), .A3(new_n832), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n388), .ZN(G1341gat));
  NAND4_X1  g636(.A1(new_n829), .A2(G127gat), .A3(new_n684), .A4(new_n832), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n820), .A2(new_n458), .A3(new_n684), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n842), .A2(KEYINPUT116), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(KEYINPUT116), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n843), .A2(new_n844), .A3(G127gat), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n840), .A2(new_n841), .A3(new_n845), .ZN(G1342gat));
  NAND3_X1  g645(.A1(new_n829), .A2(new_n614), .A3(new_n832), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(G134gat), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n821), .A2(G134gat), .A3(new_n722), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT56), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n848), .A2(KEYINPUT117), .A3(new_n850), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1343gat));
  NOR3_X1   g654(.A1(new_n546), .A2(new_n503), .A3(new_n457), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT118), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT57), .B1(new_n824), .B2(new_n534), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n534), .A2(KEYINPUT57), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n830), .A2(new_n805), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n614), .B1(new_n860), .B2(new_n812), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n584), .B1(new_n861), .B2(new_n817), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n859), .B1(new_n862), .B2(new_n819), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n857), .B1(new_n858), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G141gat), .B1(new_n864), .B2(new_n282), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n820), .A2(new_n655), .A3(new_n456), .A4(new_n534), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n282), .A2(G141gat), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT58), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n864), .A2(new_n692), .ZN(new_n871));
  AOI22_X1  g670(.A1(new_n871), .A2(G141gat), .B1(new_n867), .B2(new_n868), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(G1344gat));
  XOR2_X1   g673(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n875));
  NAND3_X1  g674(.A1(new_n824), .A2(KEYINPUT57), .A3(new_n534), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n815), .A2(new_n816), .A3(new_n722), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n584), .B1(new_n861), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n638), .A2(new_n282), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n535), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n876), .B1(KEYINPUT57), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n637), .A3(new_n857), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n875), .B1(new_n883), .B2(new_n311), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n311), .A2(KEYINPUT59), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n885), .B1(new_n864), .B2(new_n664), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n867), .A2(new_n311), .A3(new_n637), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1345gat));
  OAI21_X1  g691(.A(G155gat), .B1(new_n864), .B2(new_n584), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n867), .A2(new_n306), .A3(new_n684), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1346gat));
  NOR3_X1   g694(.A1(new_n864), .A2(new_n307), .A3(new_n814), .ZN(new_n896));
  AOI21_X1  g695(.A(G162gat), .B1(new_n867), .B2(new_n614), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(G1347gat));
  AOI21_X1  g697(.A(new_n695), .B1(new_n818), .B2(new_n819), .ZN(new_n899));
  AND4_X1   g698(.A1(new_n457), .A2(new_n899), .A3(new_n535), .A4(new_n658), .ZN(new_n900));
  INV_X1    g699(.A(G169gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n739), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT121), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n900), .A2(new_n904), .A3(new_n901), .A4(new_n739), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n824), .A2(new_n535), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n826), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n824), .A2(KEYINPUT113), .A3(new_n535), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n695), .A2(new_n657), .A3(new_n456), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n830), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G169gat), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n906), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT122), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n906), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1348gat));
  INV_X1    g717(.A(G176gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n900), .A2(new_n919), .A3(new_n637), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n910), .A2(new_n637), .A3(new_n911), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n920), .B1(new_n922), .B2(new_n919), .ZN(G1349gat));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(KEYINPUT60), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n924), .A2(KEYINPUT60), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n910), .A2(KEYINPUT123), .A3(new_n684), .A4(new_n911), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n684), .B(new_n911), .C1(new_n825), .C2(new_n827), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n927), .A2(new_n930), .A3(G183gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n900), .A2(new_n375), .A3(new_n684), .ZN(new_n932));
  AOI211_X1 g731(.A(new_n925), .B(new_n926), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  AND4_X1   g732(.A1(new_n924), .A2(new_n931), .A3(KEYINPUT60), .A4(new_n932), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(new_n934), .ZN(G1350gat));
  NAND3_X1  g734(.A1(new_n900), .A2(new_n350), .A3(new_n674), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n614), .B(new_n911), .C1(new_n825), .C2(new_n827), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n937), .A2(new_n938), .A3(G190gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n937), .B2(G190gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT125), .ZN(G1351gat));
  NOR3_X1   g741(.A1(new_n708), .A2(new_n456), .A3(new_n535), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n899), .ZN(new_n944));
  NOR4_X1   g743(.A1(new_n944), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n692), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n695), .A2(new_n456), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n655), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT127), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n881), .A3(new_n830), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G197gat), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952));
  INV_X1    g751(.A(new_n944), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n692), .A2(G197gat), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n945), .B1(new_n951), .B2(new_n955), .ZN(G1352gat));
  NOR3_X1   g755(.A1(new_n944), .A2(G204gat), .A3(new_n664), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n881), .A2(new_n637), .ZN(new_n961));
  OAI21_X1  g760(.A(G204gat), .B1(new_n948), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(G1353gat));
  OR3_X1    g762(.A1(new_n944), .A2(G211gat), .A3(new_n584), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n881), .A2(new_n684), .A3(new_n655), .A4(new_n946), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(G1354gat));
  AOI21_X1  g767(.A(G218gat), .B1(new_n953), .B2(new_n674), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n949), .A2(new_n881), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n614), .A2(G218gat), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(G1355gat));
endmodule


