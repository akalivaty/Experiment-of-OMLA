//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n188), .A2(G107), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT74), .A3(G101), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n189), .A2(new_n192), .A3(new_n196), .A4(new_n193), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(KEYINPUT74), .B1(new_n194), .B2(G101), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT75), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n199), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n197), .A2(KEYINPUT4), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT75), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .A4(new_n195), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n200), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT4), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n194), .A2(new_n206), .A3(G101), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  XNOR2_X1  g023(.A(G143), .B(G146), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n211), .A2(KEYINPUT0), .A3(G128), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n211), .B1(KEYINPUT0), .B2(G128), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n209), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  INV_X1    g031(.A(G143), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n213), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n208), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n205), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n191), .A2(KEYINPUT76), .A3(G104), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT76), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n188), .B2(G107), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n191), .A2(G104), .ZN(new_n229));
  OAI211_X1 g043(.A(G101), .B(new_n226), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT1), .B1(new_n218), .B2(G146), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n218), .A2(G146), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n216), .A2(G143), .ZN(new_n233));
  OAI211_X1 g047(.A(G128), .B(new_n231), .C1(new_n232), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G128), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n217), .B(new_n219), .C1(KEYINPUT1), .C2(new_n235), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n230), .A2(new_n234), .A3(new_n197), .A4(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT10), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT77), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(KEYINPUT77), .A3(new_n238), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT78), .B1(new_n230), .B2(new_n197), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n230), .A2(new_n197), .A3(KEYINPUT78), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n234), .A2(new_n236), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(new_n238), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n240), .A2(new_n241), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT11), .ZN(new_n249));
  INV_X1    g063(.A(G134), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n249), .B1(new_n250), .B2(G137), .ZN(new_n251));
  INV_X1    g065(.A(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT11), .A3(G134), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(G137), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G131), .ZN(new_n256));
  INV_X1    g070(.A(G131), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n251), .A2(new_n253), .A3(new_n257), .A4(new_n254), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n225), .A2(new_n248), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n244), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n247), .B1(new_n262), .B2(new_n242), .ZN(new_n263));
  INV_X1    g077(.A(new_n241), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n264), .B2(new_n239), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n223), .B1(new_n200), .B2(new_n204), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n259), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(G110), .B(G140), .ZN(new_n268));
  INV_X1    g082(.A(G953), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n269), .A2(G227), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n268), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n261), .A2(new_n267), .A3(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n265), .A2(new_n266), .ZN(new_n274));
  AND4_X1   g088(.A1(new_n236), .A2(new_n230), .A3(new_n234), .A4(new_n197), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n197), .A2(new_n230), .B1(new_n234), .B2(new_n236), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT80), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n230), .A2(new_n197), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n246), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT80), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(new_n237), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n277), .A2(new_n259), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT12), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT79), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n256), .B2(new_n258), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n285), .B(new_n286), .C1(new_n275), .C2(new_n276), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n279), .A2(new_n237), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n285), .B1(new_n289), .B2(new_n286), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n274), .A2(new_n260), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  OAI211_X1 g106(.A(G469), .B(new_n273), .C1(new_n292), .C2(new_n272), .ZN(new_n293));
  NAND2_X1  g107(.A1(G469), .A2(G902), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n284), .A2(new_n291), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n261), .A3(new_n272), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n261), .A2(new_n267), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n297), .A2(new_n298), .B1(new_n299), .B2(new_n271), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n296), .A2(new_n261), .A3(KEYINPUT81), .A4(new_n272), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G469), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n295), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT9), .B(G234), .ZN(new_n305));
  OAI21_X1  g119(.A(G221), .B1(new_n305), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n187), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n297), .A2(new_n298), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n299), .A2(new_n271), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n301), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n303), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n295), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(KEYINPUT82), .A3(new_n306), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n308), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G217), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n305), .A2(new_n318), .A3(G953), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT13), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(new_n235), .B2(G143), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n235), .A2(G143), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT87), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT87), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n218), .A2(G128), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n218), .A2(G128), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n324), .B(new_n325), .C1(new_n326), .C2(new_n320), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n322), .A2(KEYINPUT13), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT88), .A3(G134), .ZN(new_n330));
  XNOR2_X1  g144(.A(G116), .B(G122), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G107), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n191), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n322), .A2(new_n326), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n333), .A2(new_n334), .B1(new_n250), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n330), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT88), .B1(new_n329), .B2(G134), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT89), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n329), .A2(G134), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT88), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT89), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n342), .A2(new_n343), .A3(new_n330), .A4(new_n336), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n335), .B(new_n250), .ZN(new_n346));
  INV_X1    g160(.A(G116), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(KEYINPUT14), .A3(G122), .ZN(new_n348));
  OAI211_X1 g162(.A(G107), .B(new_n348), .C1(new_n332), .C2(KEYINPUT14), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n334), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n319), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n350), .ZN(new_n352));
  INV_X1    g166(.A(new_n319), .ZN(new_n353));
  AOI211_X1 g167(.A(new_n352), .B(new_n353), .C1(new_n339), .C2(new_n344), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n312), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G478), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(KEYINPUT15), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g172(.A(G113), .B(G122), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n359), .B(new_n188), .ZN(new_n360));
  XNOR2_X1  g174(.A(G125), .B(G140), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(new_n216), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  AND4_X1   g177(.A1(G143), .A2(new_n363), .A3(new_n269), .A4(G214), .ZN(new_n364));
  NOR2_X1   g178(.A1(G237), .A2(G953), .ZN(new_n365));
  AOI21_X1  g179(.A(G143), .B1(new_n365), .B2(G214), .ZN(new_n366));
  OAI211_X1 g180(.A(KEYINPUT18), .B(G131), .C1(new_n364), .C2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(new_n269), .A3(G214), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n218), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n365), .A2(G143), .A3(G214), .ZN(new_n370));
  NAND2_X1  g184(.A1(KEYINPUT18), .A2(G131), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n362), .A2(new_n367), .A3(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(G131), .B1(new_n364), .B2(new_n366), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT17), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n369), .A2(new_n257), .A3(new_n370), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G125), .ZN(new_n380));
  INV_X1    g194(.A(G125), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G140), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT16), .ZN(new_n383));
  OR3_X1    g197(.A1(new_n381), .A2(KEYINPUT16), .A3(G140), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n216), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n383), .A2(new_n384), .A3(G146), .ZN(new_n387));
  OAI211_X1 g201(.A(KEYINPUT17), .B(G131), .C1(new_n364), .C2(new_n366), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n360), .B(new_n373), .C1(new_n378), .C2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n377), .A2(new_n386), .A3(new_n387), .A4(new_n388), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n360), .B1(new_n392), .B2(new_n373), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n312), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT86), .B(G475), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G952), .ZN(new_n397));
  AOI211_X1 g211(.A(G953), .B(new_n397), .C1(G234), .C2(G237), .ZN(new_n398));
  AOI211_X1 g212(.A(new_n312), .B(new_n269), .C1(G234), .C2(G237), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT21), .B(G898), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n374), .A2(new_n376), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n380), .A2(new_n382), .A3(KEYINPUT19), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT19), .B1(new_n380), .B2(new_n382), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n216), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n387), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n373), .ZN(new_n409));
  INV_X1    g223(.A(new_n360), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(new_n390), .ZN(new_n412));
  NOR2_X1   g226(.A1(G475), .A2(G902), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n403), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n413), .ZN(new_n415));
  AOI211_X1 g229(.A(KEYINPUT20), .B(new_n415), .C1(new_n411), .C2(new_n390), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n396), .B(new_n402), .C1(new_n414), .C2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  OAI221_X1 g232(.A(new_n312), .B1(KEYINPUT15), .B2(new_n356), .C1(new_n351), .C2(new_n354), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n358), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT90), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT90), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n358), .A2(new_n418), .A3(new_n419), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G214), .B1(G237), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(KEYINPUT2), .A2(G113), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT68), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OR2_X1    g245(.A1(KEYINPUT2), .A2(G113), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G119), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G116), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n347), .A2(G119), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT5), .ZN(new_n439));
  OAI21_X1  g253(.A(G113), .B1(new_n435), .B2(KEYINPUT5), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n245), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G110), .B(G122), .ZN(new_n444));
  AND2_X1   g258(.A1(new_n200), .A2(new_n204), .ZN(new_n445));
  INV_X1    g259(.A(new_n437), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n431), .B2(new_n432), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n208), .B1(new_n447), .B2(new_n438), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n443), .B(new_n444), .C1(new_n445), .C2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n444), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n448), .B1(new_n200), .B2(new_n204), .ZN(new_n451));
  INV_X1    g265(.A(new_n443), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n449), .A2(new_n453), .A3(KEYINPUT6), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n246), .A2(new_n381), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n213), .A2(new_n221), .A3(G125), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G224), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G953), .ZN(new_n459));
  XOR2_X1   g273(.A(new_n459), .B(KEYINPUT83), .Z(new_n460));
  XNOR2_X1  g274(.A(new_n457), .B(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n462), .B(new_n450), .C1(new_n451), .C2(new_n452), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n454), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n442), .A2(new_n278), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n444), .B(KEYINPUT8), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n439), .A2(KEYINPUT84), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(new_n440), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n439), .A2(KEYINPUT84), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n438), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n465), .B(new_n466), .C1(new_n470), .C2(new_n278), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n456), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT7), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n457), .B(new_n473), .C1(new_n474), .C2(new_n459), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n473), .B1(new_n474), .B2(new_n459), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n456), .A3(new_n455), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n471), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(G902), .B1(new_n478), .B2(new_n449), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n464), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G210), .B1(G237), .B2(G902), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n464), .A2(new_n479), .A3(new_n481), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n426), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n424), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT32), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n259), .A2(new_n222), .ZN(new_n489));
  INV_X1    g303(.A(new_n254), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n250), .A2(G137), .ZN(new_n491));
  OAI21_X1  g305(.A(G131), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(new_n234), .A3(new_n236), .A4(new_n258), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n489), .A2(KEYINPUT30), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT66), .ZN(new_n495));
  INV_X1    g309(.A(new_n209), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT0), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n235), .A3(KEYINPUT65), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n220), .B2(new_n498), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n209), .A2(new_n214), .B1(new_n217), .B2(new_n219), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n213), .A2(new_n221), .A3(KEYINPUT66), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n259), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT67), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT67), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n501), .A2(new_n505), .A3(new_n502), .A4(new_n259), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n493), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n494), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n433), .B(new_n446), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT31), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT26), .B(G101), .Z(new_n514));
  NAND2_X1  g328(.A1(new_n365), .A2(G210), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n510), .A2(new_n489), .A3(new_n493), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n512), .A2(new_n513), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n507), .A2(new_n511), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(KEYINPUT28), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT28), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n510), .A2(new_n489), .A3(new_n525), .A4(new_n493), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n518), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT71), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n507), .A2(new_n511), .B1(new_n524), .B2(new_n526), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT71), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n531), .A2(new_n532), .A3(new_n518), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n522), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT70), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n520), .B1(new_n509), .B2(new_n511), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(new_n513), .ZN(new_n537));
  AOI211_X1 g351(.A(new_n510), .B(new_n494), .C1(new_n507), .C2(new_n508), .ZN(new_n538));
  OAI211_X1 g352(.A(KEYINPUT70), .B(KEYINPUT31), .C1(new_n538), .C2(new_n520), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n534), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(G472), .A2(G902), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n488), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n489), .A2(new_n493), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n511), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n527), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT29), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n518), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n528), .A2(KEYINPUT29), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n312), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n529), .A2(new_n519), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n512), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n553), .A2(KEYINPUT29), .ZN(new_n554));
  OAI21_X1  g368(.A(G472), .B1(new_n550), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n537), .A2(new_n539), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n528), .A2(KEYINPUT71), .A3(new_n529), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n532), .B1(new_n531), .B2(new_n518), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n557), .A2(new_n558), .B1(new_n536), .B2(new_n513), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(KEYINPUT32), .A3(new_n541), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n543), .A2(new_n555), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT23), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n434), .B2(G128), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n235), .A2(KEYINPUT23), .A3(G119), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n564), .B(new_n565), .C1(G119), .C2(new_n235), .ZN(new_n566));
  XNOR2_X1  g380(.A(G119), .B(G128), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT24), .B(G110), .Z(new_n568));
  AOI22_X1  g382(.A1(new_n566), .A2(G110), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n387), .ZN(new_n570));
  AOI21_X1  g384(.A(G146), .B1(new_n383), .B2(new_n384), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI22_X1  g386(.A1(new_n566), .A2(G110), .B1(new_n567), .B2(new_n568), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n361), .A2(new_n216), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n573), .A2(new_n387), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT22), .B(G137), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n269), .A2(G221), .A3(G234), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n572), .A2(new_n575), .A3(new_n579), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n312), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(KEYINPUT73), .A2(KEYINPUT25), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n584), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n581), .A2(new_n312), .A3(new_n582), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(KEYINPUT73), .A2(KEYINPUT25), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G234), .ZN(new_n590));
  OAI21_X1  g404(.A(G217), .B1(new_n590), .B2(G902), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT72), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n581), .A2(new_n582), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(G902), .B1(new_n590), .B2(G217), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n317), .A2(new_n487), .A3(new_n562), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(KEYINPUT91), .B(G101), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(G3));
  NOR2_X1   g416(.A1(new_n356), .A2(new_n312), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n345), .A2(new_n350), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n353), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n345), .A2(new_n350), .A3(new_n319), .ZN(new_n606));
  AOI21_X1  g420(.A(G902), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n603), .B1(new_n607), .B2(new_n356), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n605), .A2(new_n609), .A3(new_n606), .ZN(new_n610));
  OAI21_X1  g424(.A(KEYINPUT33), .B1(new_n351), .B2(new_n354), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n610), .A2(new_n611), .A3(G478), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n396), .B1(new_n414), .B2(new_n416), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n483), .A2(KEYINPUT93), .A3(new_n484), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n464), .A2(new_n618), .A3(new_n479), .A4(new_n481), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n619), .A2(new_n425), .ZN(new_n620));
  AND4_X1   g434(.A1(new_n402), .A2(new_n616), .A3(new_n617), .A4(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(G902), .B1(new_n556), .B2(new_n559), .ZN(new_n622));
  INV_X1    g436(.A(G472), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(KEYINPUT92), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  AOI211_X1 g440(.A(G902), .B(new_n624), .C1(new_n556), .C2(new_n559), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n626), .A2(new_n627), .A3(new_n598), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n317), .A2(new_n621), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT34), .B(G104), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n629), .B(new_n630), .ZN(G6));
  AOI21_X1  g445(.A(new_n614), .B1(new_n358), .B2(new_n419), .ZN(new_n632));
  AND4_X1   g446(.A1(new_n402), .A2(new_n617), .A3(new_n620), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n317), .A2(new_n628), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  OAI21_X1  g450(.A(new_n576), .B1(KEYINPUT36), .B2(new_n580), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT36), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n572), .A2(new_n575), .A3(new_n638), .A4(new_n579), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n637), .A2(new_n596), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT94), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT94), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n637), .A2(new_n642), .A3(new_n596), .A4(new_n639), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n589), .B2(new_n592), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n626), .A2(new_n627), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n317), .A2(new_n487), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT95), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT37), .B(G110), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  NAND2_X1  g464(.A1(new_n617), .A2(new_n620), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT32), .B1(new_n560), .B2(new_n541), .ZN(new_n652));
  AOI211_X1 g466(.A(new_n488), .B(new_n542), .C1(new_n556), .C2(new_n559), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n651), .B1(new_n654), .B2(new_n555), .ZN(new_n655));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n399), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n398), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n632), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n645), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n308), .B2(new_n316), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n655), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  XNOR2_X1  g479(.A(new_n659), .B(KEYINPUT39), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n317), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n529), .B1(new_n512), .B2(new_n519), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n552), .A2(new_n545), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n312), .ZN(new_n672));
  OAI21_X1  g486(.A(G472), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT96), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n543), .A2(new_n561), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n483), .A2(new_n484), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT38), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n615), .B1(new_n358), .B2(new_n419), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n679), .A2(new_n425), .A3(new_n645), .A4(new_n680), .ZN(new_n681));
  NOR4_X1   g495(.A1(new_n668), .A2(new_n669), .A3(new_n677), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n218), .ZN(G45));
  NAND4_X1  g497(.A1(new_n608), .A2(new_n614), .A3(new_n612), .A4(new_n659), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n645), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n655), .A2(new_n317), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  NAND2_X1  g501(.A1(new_n311), .A2(new_n312), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G469), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n306), .A3(new_n313), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n621), .A2(new_n562), .A3(new_n599), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND4_X1  g508(.A1(new_n562), .A2(new_n633), .A3(new_n691), .A4(new_n599), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NOR2_X1   g510(.A1(new_n690), .A2(new_n651), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(new_n562), .A3(new_n424), .A4(new_n661), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  NAND4_X1  g513(.A1(new_n689), .A2(new_n306), .A3(new_n313), .A4(new_n402), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n546), .A2(KEYINPUT97), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n529), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n546), .A2(KEYINPUT97), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n522), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n536), .A2(new_n513), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n541), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n599), .B(new_n706), .C1(new_n622), .C2(new_n623), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n617), .A2(new_n620), .A3(new_n680), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  OAI211_X1 g525(.A(new_n661), .B(new_n706), .C1(new_n622), .C2(new_n623), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n684), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n697), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  AOI21_X1  g529(.A(new_n598), .B1(new_n654), .B2(new_n555), .ZN(new_n716));
  INV_X1    g530(.A(new_n684), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n294), .B(KEYINPUT98), .Z(new_n718));
  NAND2_X1  g532(.A1(new_n293), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n302), .B2(new_n303), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n483), .A2(new_n425), .A3(new_n484), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n720), .A2(new_n721), .A3(new_n307), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n716), .A2(new_n717), .A3(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT99), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n724), .A2(KEYINPUT42), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n723), .A2(new_n725), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G131), .ZN(G33));
  OR2_X1    g544(.A1(new_n660), .A2(KEYINPUT100), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n660), .A2(KEYINPUT100), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n716), .A2(new_n722), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  NAND3_X1  g548(.A1(new_n608), .A2(new_n615), .A3(new_n612), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n735), .B(KEYINPUT43), .Z(new_n736));
  OAI211_X1 g550(.A(new_n736), .B(new_n661), .C1(new_n627), .C2(new_n626), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n721), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n738), .B2(new_n737), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n273), .B1(new_n292), .B2(new_n272), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n303), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n742), .B2(new_n741), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(KEYINPUT101), .ZN(new_n745));
  INV_X1    g559(.A(new_n718), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(KEYINPUT46), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n313), .B1(new_n747), .B2(KEYINPUT46), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n306), .B(new_n666), .C1(new_n748), .C2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n740), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n252), .ZN(G39));
  OAI21_X1  g566(.A(new_n306), .B1(new_n748), .B2(new_n749), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT47), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n562), .A2(new_n599), .A3(new_n684), .A4(new_n721), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(KEYINPUT102), .B(G140), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G42));
  NAND2_X1  g575(.A1(new_n689), .A2(new_n313), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT49), .Z(new_n763));
  NOR3_X1   g577(.A1(new_n598), .A2(new_n307), .A3(new_n426), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT103), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n679), .A2(new_n765), .A3(new_n735), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(new_n766), .A3(new_n677), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n713), .A2(new_n722), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n358), .A2(new_n419), .A3(new_n615), .A4(new_n659), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(KEYINPUT106), .Z(new_n770));
  INV_X1    g584(.A(new_n721), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n562), .A2(new_n770), .A3(new_n661), .A4(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n317), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n768), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n728), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n733), .B(new_n775), .C1(new_n776), .C2(new_n726), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n616), .A2(new_n632), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n485), .A2(new_n402), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n317), .A2(new_n628), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  AND4_X1   g596(.A1(KEYINPUT105), .A2(new_n600), .A3(new_n782), .A4(new_n647), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n486), .B1(new_n308), .B2(new_n316), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n716), .B2(new_n646), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT105), .B1(new_n785), .B2(new_n782), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n692), .A2(new_n698), .A3(new_n695), .A4(new_n710), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n778), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT109), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT82), .B1(new_n315), .B2(new_n306), .ZN(new_n793));
  AOI211_X1 g607(.A(new_n187), .B(new_n307), .C1(new_n313), .C2(new_n314), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n660), .B(new_n661), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n651), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n562), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n714), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n644), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n593), .A2(new_n799), .A3(new_n659), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT107), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT107), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n645), .A2(new_n802), .A3(new_n659), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n720), .A2(new_n804), .A3(new_n307), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n676), .A2(new_n709), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n685), .B1(new_n793), .B2(new_n794), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n806), .B1(new_n807), .B2(new_n797), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT52), .B1(new_n798), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT108), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n798), .B2(new_n808), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n655), .A2(new_n663), .B1(new_n697), .B2(new_n713), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(KEYINPUT108), .A3(new_n686), .A4(new_n806), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n792), .B(new_n809), .C1(new_n814), .C2(KEYINPUT52), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT52), .B1(new_n811), .B2(new_n813), .ZN(new_n816));
  INV_X1    g630(.A(new_n809), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT109), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n791), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n811), .A2(new_n813), .A3(KEYINPUT52), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n816), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n788), .A2(KEYINPUT104), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n424), .A2(new_n661), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n823), .B1(new_n654), .B2(new_n555), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n824), .A2(new_n697), .B1(new_n709), .B2(new_n708), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT104), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n825), .A2(new_n826), .A3(new_n692), .A4(new_n695), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n822), .B(new_n827), .C1(new_n783), .C2(new_n786), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n777), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT53), .B1(new_n821), .B2(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n819), .A2(new_n830), .A3(KEYINPUT54), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n821), .A2(new_n829), .A3(KEYINPUT53), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT110), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n821), .A2(new_n829), .A3(KEYINPUT110), .A4(KEYINPUT53), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n828), .B(new_n777), .C1(new_n815), .C2(new_n818), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(KEYINPUT53), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n831), .B1(new_n837), .B2(KEYINPUT54), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n691), .A2(new_n426), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT111), .ZN(new_n840));
  INV_X1    g654(.A(new_n679), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n736), .A2(new_n398), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n707), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n690), .A2(new_n721), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n677), .A2(new_n599), .A3(new_n398), .A4(new_n847), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n848), .A2(KEYINPUT115), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(KEYINPUT115), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n849), .A2(new_n615), .A3(new_n613), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n847), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n842), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(KEYINPUT113), .ZN(new_n854));
  INV_X1    g668(.A(new_n712), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n856), .A2(KEYINPUT114), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT114), .B1(new_n854), .B2(new_n855), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n846), .B(new_n851), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n755), .B(new_n756), .C1(new_n306), .C2(new_n762), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n860), .A2(new_n771), .A3(new_n843), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n849), .A2(new_n616), .A3(new_n850), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n397), .B(G953), .C1(new_n843), .C2(new_n697), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT48), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n854), .A2(new_n866), .A3(new_n716), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n866), .B1(new_n854), .B2(new_n716), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n864), .B(new_n865), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT116), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n862), .B1(new_n859), .B2(new_n861), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n838), .A2(new_n863), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n767), .B1(new_n872), .B2(new_n873), .ZN(G75));
  NOR2_X1   g688(.A1(new_n269), .A2(G952), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT119), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n815), .A2(new_n818), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n787), .A3(new_n778), .A4(new_n790), .ZN(new_n879));
  INV_X1    g693(.A(new_n830), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n312), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(G210), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT56), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n454), .A2(new_n463), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT117), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT118), .Z(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(new_n461), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n884), .A2(new_n889), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n877), .B1(new_n890), .B2(new_n891), .ZN(G51));
  NAND2_X1  g706(.A1(new_n879), .A2(new_n880), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT54), .ZN(new_n894));
  INV_X1    g708(.A(new_n831), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  XOR2_X1   g711(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n898));
  XNOR2_X1  g712(.A(new_n718), .B(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n311), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n881), .A2(new_n745), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n875), .B1(new_n900), .B2(new_n901), .ZN(G54));
  NAND3_X1  g716(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .ZN(new_n903));
  INV_X1    g717(.A(new_n412), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n905), .A2(new_n906), .A3(new_n875), .ZN(G60));
  INV_X1    g721(.A(KEYINPUT122), .ZN(new_n908));
  XOR2_X1   g722(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n603), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n834), .A2(new_n835), .ZN(new_n911));
  AOI21_X1  g725(.A(KEYINPUT53), .B1(new_n878), .B2(new_n829), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT54), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n910), .B1(new_n913), .B2(new_n895), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n610), .A2(new_n611), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n908), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n915), .ZN(new_n917));
  OAI211_X1 g731(.A(KEYINPUT122), .B(new_n917), .C1(new_n838), .C2(new_n910), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n910), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n877), .B1(new_n896), .B2(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n916), .A2(new_n918), .A3(new_n920), .ZN(G63));
  AND2_X1   g735(.A1(new_n637), .A2(new_n639), .ZN(new_n922));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n893), .A2(new_n922), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n924), .B1(new_n879), .B2(new_n880), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n926), .B(new_n876), .C1(new_n595), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT61), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n928), .A2(new_n929), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n893), .A2(new_n925), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n877), .B1(new_n934), .B2(new_n594), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n935), .A2(new_n930), .A3(new_n931), .A4(new_n926), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n933), .A2(new_n936), .ZN(G66));
  NAND2_X1  g751(.A1(new_n828), .A2(new_n269), .ZN(new_n938));
  OAI21_X1  g752(.A(G953), .B1(new_n400), .B2(new_n458), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n938), .A2(KEYINPUT124), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(KEYINPUT124), .B2(new_n938), .ZN(new_n941));
  INV_X1    g755(.A(G898), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n886), .B1(new_n942), .B2(G953), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(G69));
  XNOR2_X1  g758(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n716), .A2(new_n771), .A3(new_n779), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(new_n667), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n751), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n812), .A2(new_n686), .ZN(new_n950));
  OR3_X1    g764(.A1(new_n682), .A2(KEYINPUT62), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(KEYINPUT62), .B1(new_n682), .B2(new_n950), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n759), .A2(new_n949), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n269), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n405), .A2(new_n406), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT125), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n509), .B(new_n956), .Z(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(G900), .A2(G953), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n751), .A2(new_n950), .ZN(new_n961));
  INV_X1    g775(.A(new_n733), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n727), .B2(new_n728), .ZN(new_n963));
  INV_X1    g777(.A(new_n750), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n964), .A2(new_n716), .A3(new_n709), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n759), .A2(new_n961), .A3(new_n963), .A4(new_n965), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n957), .B(new_n960), .C1(new_n966), .C2(G953), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n269), .B1(G227), .B2(G900), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n959), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n969), .B1(new_n959), .B2(new_n967), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n946), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n972), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n945), .A3(new_n970), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n975), .ZN(G72));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT63), .Z(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n953), .B2(new_n828), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n670), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n966), .A2(new_n828), .ZN(new_n981));
  INV_X1    g795(.A(new_n978), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI221_X1 g797(.A(new_n980), .B1(G952), .B2(new_n269), .C1(new_n983), .C2(new_n553), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n982), .B(new_n670), .C1(new_n512), .C2(new_n552), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n984), .B1(new_n837), .B2(new_n985), .ZN(G57));
endmodule


