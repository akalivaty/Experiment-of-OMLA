//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n533, new_n534, new_n535,
    new_n536, new_n539, new_n540, new_n541, new_n542, new_n544, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1135, new_n1136,
    new_n1137, new_n1138;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT65), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g040(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(KEYINPUT3), .B1(KEYINPUT66), .B2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G137), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(new_n470), .ZN(G160));
  INV_X1    g046(.A(KEYINPUT67), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n472), .B1(new_n466), .B2(new_n467), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT66), .A2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(KEYINPUT66), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(KEYINPUT67), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n473), .A2(new_n478), .A3(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n473), .A2(new_n478), .A3(new_n461), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND3_X1  g063(.A1(new_n462), .A2(G138), .A3(new_n461), .ZN(new_n489));
  OAI21_X1  g064(.A(G126), .B1(new_n466), .B2(new_n467), .ZN(new_n490));
  NAND2_X1  g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n461), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(KEYINPUT4), .B(G138), .C1(new_n466), .C2(new_n467), .ZN(new_n495));
  NAND2_X1  g070(.A1(G102), .A2(G2104), .ZN(new_n496));
  AOI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n501), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(KEYINPUT68), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT6), .A3(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n515), .A2(new_n506), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n509), .A2(G651), .B1(new_n516), .B2(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT69), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR3_X1    g095(.A1(new_n518), .A2(KEYINPUT69), .A3(new_n519), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n517), .A2(new_n520), .A3(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  XNOR2_X1  g098(.A(new_n518), .B(KEYINPUT72), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n524), .A2(G51), .B1(G89), .B2(new_n516), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT71), .ZN(new_n527));
  XOR2_X1   g102(.A(KEYINPUT73), .B(KEYINPUT7), .Z(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n525), .A2(new_n527), .A3(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(new_n524), .A2(G52), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n511), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n516), .A2(G90), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AND2_X1   g113(.A1(new_n516), .A2(G81), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n511), .ZN(new_n541));
  AOI211_X1 g116(.A(new_n539), .B(new_n541), .C1(new_n524), .C2(G43), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(G188));
  NAND2_X1  g123(.A1(new_n516), .A2(G91), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT76), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n549), .B(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n511), .ZN(new_n553));
  NAND2_X1  g128(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n554));
  NAND2_X1  g129(.A1(G53), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n515), .A2(new_n554), .A3(new_n558), .ZN(new_n559));
  AOI211_X1 g134(.A(new_n556), .B(new_n555), .C1(new_n512), .C2(new_n514), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n560), .B2(new_n554), .ZN(new_n561));
  AND2_X1   g136(.A1(new_n553), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n551), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT77), .ZN(G299));
  INV_X1    g139(.A(new_n518), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G49), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n516), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(new_n506), .A2(G61), .ZN(new_n570));
  INV_X1    g145(.A(G73), .ZN(new_n571));
  OAI21_X1  g146(.A(KEYINPUT78), .B1(new_n571), .B2(new_n503), .ZN(new_n572));
  OR3_X1    g147(.A1(new_n571), .A2(new_n503), .A3(KEYINPUT78), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n565), .A2(G48), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n516), .A2(G86), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n524), .A2(G47), .B1(G85), .B2(new_n516), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT79), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n511), .B2(new_n581), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n516), .A2(G92), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT10), .Z(new_n585));
  NAND2_X1  g160(.A1(new_n524), .A2(G54), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  XNOR2_X1  g162(.A(KEYINPUT80), .B(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n507), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n583), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n583), .B1(new_n592), .B2(G868), .ZN(G321));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n563), .B(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n595), .B1(new_n597), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n595), .B1(new_n597), .B2(G868), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n592), .B1(new_n600), .B2(G860), .ZN(G148));
  NOR2_X1   g176(.A1(new_n591), .A2(G559), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g181(.A1(new_n480), .A2(G123), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n483), .A2(G135), .ZN(new_n608));
  OR2_X1    g183(.A1(G99), .A2(G2105), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n609), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(new_n611), .B(G2096), .Z(new_n612));
  NAND3_X1  g187(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n612), .A2(new_n616), .ZN(G156));
  XNOR2_X1  g192(.A(KEYINPUT15), .B(G2430), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2435), .ZN(new_n619));
  XOR2_X1   g194(.A(G2427), .B(G2438), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(KEYINPUT14), .ZN(new_n622));
  XOR2_X1   g197(.A(G2451), .B(G2454), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT16), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n622), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G1341), .B(G1348), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n627), .B(new_n628), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G14), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(G401));
  XOR2_X1   g206(.A(G2084), .B(G2090), .Z(new_n632));
  XNOR2_X1  g207(.A(G2072), .B(G2078), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2067), .B(G2678), .Z(new_n635));
  AOI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n633), .B(KEYINPUT17), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n636), .B1(new_n638), .B2(new_n635), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT81), .Z(new_n640));
  INV_X1    g215(.A(new_n635), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n641), .A2(new_n633), .A3(new_n632), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT18), .Z(new_n643));
  NAND3_X1  g218(.A1(new_n638), .A2(new_n632), .A3(new_n635), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n640), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT82), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2096), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(G2100), .Z(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G227));
  XNOR2_X1  g224(.A(G1971), .B(G1976), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT83), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT19), .Z(new_n652));
  XOR2_X1   g227(.A(G1956), .B(G2474), .Z(new_n653));
  XOR2_X1   g228(.A(G1961), .B(G1966), .Z(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n653), .A2(new_n654), .ZN(new_n658));
  AOI22_X1  g233(.A1(new_n656), .A2(new_n657), .B1(new_n652), .B2(new_n658), .ZN(new_n659));
  OR3_X1    g234(.A1(new_n652), .A2(new_n655), .A3(new_n658), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n659), .B(new_n660), .C1(new_n657), .C2(new_n656), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1991), .B(G1996), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G1981), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n661), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT84), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G229));
  XOR2_X1   g243(.A(KEYINPUT96), .B(KEYINPUT23), .Z(new_n669));
  INV_X1    g244(.A(G16), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(G20), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(new_n597), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G1956), .ZN(new_n674));
  INV_X1    g249(.A(G29), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G35), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(G162), .B2(new_n675), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT29), .Z(new_n678));
  INV_X1    g253(.A(G2090), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n681), .A2(KEYINPUT97), .ZN(new_n682));
  NOR2_X1   g257(.A1(G4), .A2(G16), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n592), .B2(G16), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(G1348), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(G1348), .ZN(new_n687));
  OAI21_X1  g262(.A(G29), .B1(new_n465), .B2(new_n470), .ZN(new_n688));
  INV_X1    g263(.A(G34), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n689), .A2(KEYINPUT24), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(KEYINPUT24), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n675), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(G2084), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT95), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT30), .B(G28), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n695), .B1(new_n675), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT31), .B(G11), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n687), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n611), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(G29), .B2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G1341), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n542), .A2(G16), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G16), .B2(G19), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n686), .B(new_n701), .C1(new_n702), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(G168), .A2(G16), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G16), .B2(G21), .ZN(new_n707));
  INV_X1    g282(.A(G1966), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT93), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT94), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G5), .B2(G16), .ZN(new_n712));
  OR3_X1    g287(.A1(new_n711), .A2(G5), .A3(G16), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n712), .B(new_n713), .C1(G301), .C2(new_n670), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1961), .ZN(new_n715));
  NAND2_X1  g290(.A1(G164), .A2(G29), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G27), .B2(G29), .ZN(new_n717));
  INV_X1    g292(.A(G2078), .ZN(new_n718));
  INV_X1    g293(.A(G2072), .ZN(new_n719));
  OR2_X1    g294(.A1(G29), .A2(G33), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n462), .A2(G127), .ZN(new_n721));
  AND2_X1   g296(.A1(G115), .A2(G2104), .ZN(new_n722));
  OAI21_X1  g297(.A(G2105), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT25), .Z(new_n725));
  INV_X1    g300(.A(G139), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n723), .B(new_n725), .C1(new_n482), .C2(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n720), .B1(new_n727), .B2(new_n675), .ZN(new_n728));
  OAI22_X1  g303(.A1(new_n717), .A2(new_n718), .B1(new_n719), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n719), .B2(new_n728), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n710), .A2(new_n715), .A3(new_n730), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n681), .A2(KEYINPUT97), .B1(new_n679), .B2(new_n678), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n707), .A2(new_n708), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n717), .A2(new_n718), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n731), .A2(new_n732), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n675), .A2(G26), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT28), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n480), .A2(G128), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n483), .A2(G140), .ZN(new_n739));
  NOR2_X1   g314(.A1(G104), .A2(G2105), .ZN(new_n740));
  OAI21_X1  g315(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n738), .B(new_n739), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G29), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(KEYINPUT91), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n737), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2067), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n705), .A2(new_n735), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n704), .A2(new_n702), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n480), .A2(G119), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n483), .A2(G131), .ZN(new_n751));
  OR2_X1    g326(.A1(G95), .A2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  MUX2_X1   g329(.A(G25), .B(new_n754), .S(G29), .Z(new_n755));
  XOR2_X1   g330(.A(KEYINPUT35), .B(G1991), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT85), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n755), .B(new_n757), .ZN(new_n758));
  MUX2_X1   g333(.A(G24), .B(G290), .S(G16), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1986), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n758), .B(new_n760), .C1(KEYINPUT90), .C2(KEYINPUT36), .ZN(new_n761));
  NOR2_X1   g336(.A1(G6), .A2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G305), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(G16), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT32), .B(G1981), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n670), .A2(G22), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G166), .B2(new_n670), .ZN(new_n770));
  INV_X1    g345(.A(G1971), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n670), .A2(G23), .ZN(new_n773));
  INV_X1    g348(.A(G288), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n774), .B2(new_n670), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1976), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT88), .B(KEYINPUT33), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n768), .A2(new_n772), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT89), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT34), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n779), .A2(new_n780), .ZN(new_n783));
  AND3_X1   g358(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n782), .B1(new_n781), .B2(new_n783), .ZN(new_n785));
  OAI221_X1 g360(.A(new_n761), .B1(KEYINPUT90), .B2(KEYINPUT36), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n761), .B1(new_n784), .B2(new_n785), .ZN(new_n787));
  NOR2_X1   g362(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n748), .A2(new_n749), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n693), .ZN(new_n791));
  INV_X1    g366(.A(G2084), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n480), .A2(G129), .ZN(new_n794));
  NAND3_X1  g369(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT92), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT26), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n483), .A2(G141), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n794), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n801), .A2(G29), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G29), .B2(G32), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT27), .B(G1996), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NOR3_X1   g380(.A1(new_n790), .A2(new_n793), .A3(new_n805), .ZN(G311));
  AND3_X1   g381(.A1(new_n748), .A2(new_n786), .A3(new_n789), .ZN(new_n807));
  INV_X1    g382(.A(new_n793), .ZN(new_n808));
  INV_X1    g383(.A(new_n805), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n807), .A2(new_n808), .A3(new_n809), .A4(new_n749), .ZN(G150));
  AOI22_X1  g385(.A1(new_n524), .A2(G55), .B1(G93), .B2(new_n516), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n511), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G860), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT98), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT37), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n813), .A2(new_n542), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n813), .A2(new_n542), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n591), .A2(new_n600), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n816), .B1(new_n823), .B2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT99), .Z(G145));
  INV_X1    g400(.A(G142), .ZN(new_n826));
  NOR2_X1   g401(.A1(G106), .A2(G2105), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(new_n461), .B2(G118), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n482), .A2(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(G130), .B2(new_n480), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n800), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT100), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G160), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n727), .B(new_n499), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n614), .B(KEYINPUT101), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n833), .A2(new_n836), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n742), .B(new_n754), .Z(new_n840));
  XOR2_X1   g415(.A(new_n611), .B(new_n487), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT102), .B(G37), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n839), .A2(new_n842), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT103), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n843), .A2(new_n848), .A3(new_n844), .A4(new_n845), .ZN(new_n849));
  AND3_X1   g424(.A1(new_n847), .A2(KEYINPUT40), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT40), .B1(new_n847), .B2(new_n849), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(new_n851), .ZN(G395));
  XNOR2_X1  g427(.A(G290), .B(G288), .ZN(new_n853));
  XNOR2_X1  g428(.A(G303), .B(G305), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n853), .B(new_n854), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT42), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT41), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n597), .A2(new_n591), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n597), .A2(new_n591), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(G299), .A2(new_n592), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(new_n862), .A3(KEYINPUT41), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n819), .B(new_n603), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n859), .A2(new_n860), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(new_n865), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n856), .B(new_n868), .ZN(new_n869));
  MUX2_X1   g444(.A(new_n813), .B(new_n869), .S(G868), .Z(G295));
  MUX2_X1   g445(.A(new_n813), .B(new_n869), .S(G868), .Z(G331));
  INV_X1    g446(.A(new_n864), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n819), .A2(G171), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n817), .A2(G301), .A3(new_n818), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n873), .A2(G168), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(G168), .B1(new_n873), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT104), .B1(new_n872), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n859), .B2(new_n860), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n864), .B(new_n880), .C1(new_n875), .C2(new_n876), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n855), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  INV_X1    g460(.A(new_n855), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n886), .A2(new_n879), .A3(new_n878), .A4(new_n881), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n883), .A2(new_n884), .A3(new_n885), .A4(new_n887), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n888), .A2(KEYINPUT106), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n867), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n864), .B2(KEYINPUT105), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n879), .B1(new_n892), .B2(new_n877), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n855), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n887), .A2(new_n894), .A3(new_n844), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n890), .B1(new_n895), .B2(KEYINPUT43), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n888), .A2(KEYINPUT106), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n889), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n887), .A2(new_n894), .A3(new_n884), .A4(new_n844), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n899), .B1(new_n900), .B2(new_n884), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n890), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n898), .A2(new_n902), .ZN(G397));
  INV_X1    g478(.A(G1384), .ZN(new_n904));
  INV_X1    g479(.A(new_n489), .ZN(new_n905));
  INV_X1    g480(.A(G126), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n906), .B1(new_n476), .B2(new_n477), .ZN(new_n907));
  INV_X1    g482(.A(new_n491), .ZN(new_n908));
  OAI21_X1  g483(.A(G2105), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n905), .B1(new_n909), .B2(KEYINPUT4), .ZN(new_n910));
  OAI211_X1 g485(.A(KEYINPUT45), .B(new_n904), .C1(new_n910), .C2(new_n497), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n904), .B1(new_n910), .B2(new_n497), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT45), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G40), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n465), .A2(new_n470), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n914), .A2(new_n912), .A3(new_n915), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n771), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT111), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n919), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT50), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n914), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n499), .A2(KEYINPUT50), .A3(new_n904), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n679), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n921), .A2(KEYINPUT111), .A3(new_n771), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n924), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT112), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n924), .A2(KEYINPUT112), .A3(new_n930), .A4(new_n931), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(G8), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(G303), .A2(G8), .ZN(new_n937));
  XOR2_X1   g512(.A(new_n937), .B(KEYINPUT55), .Z(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n934), .A2(G8), .A3(new_n938), .A4(new_n935), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n499), .A2(new_n904), .A3(new_n919), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G8), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(G1976), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n945), .B1(new_n946), .B2(G288), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT52), .B1(G288), .B2(new_n946), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(KEYINPUT114), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n949), .B1(KEYINPUT114), .B2(new_n948), .ZN(new_n950));
  OR2_X1    g525(.A1(G305), .A2(G1981), .ZN(new_n951));
  NAND2_X1  g526(.A1(G305), .A2(G1981), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT49), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n951), .A2(KEYINPUT49), .A3(new_n952), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n945), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT113), .B1(new_n947), .B2(KEYINPUT52), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n947), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n950), .B(new_n957), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(KEYINPUT116), .B(G2084), .Z(new_n962));
  NAND2_X1  g537(.A1(new_n929), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n916), .A2(new_n919), .A3(new_n911), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n708), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n944), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n967), .A2(G286), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n940), .A2(new_n941), .A3(new_n961), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT63), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n957), .A2(new_n946), .A3(new_n774), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n951), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT115), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n971), .A2(KEYINPUT115), .A3(new_n951), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n945), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n941), .B2(new_n960), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n970), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n922), .A2(new_n930), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n939), .B1(new_n980), .B2(new_n944), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n961), .A2(new_n981), .A3(new_n941), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT56), .B(G2072), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n917), .A2(new_n919), .A3(new_n920), .A4(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT118), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n561), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n986), .A2(KEYINPUT57), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n563), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n551), .B(new_n562), .C1(new_n986), .C2(KEYINPUT57), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT50), .B1(new_n499), .B2(new_n904), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n926), .B(G1384), .C1(new_n494), .C2(new_n498), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n919), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(KEYINPUT117), .B(G1956), .Z(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n984), .A2(new_n990), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n990), .B1(new_n984), .B2(new_n995), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n942), .A2(G2067), .ZN(new_n998));
  INV_X1    g573(.A(G1348), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(new_n591), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n996), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n984), .A2(new_n995), .ZN(new_n1003));
  INV_X1    g578(.A(new_n990), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(KEYINPUT61), .A3(new_n996), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1005), .A2(KEYINPUT119), .A3(KEYINPUT61), .A4(new_n996), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n998), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n929), .B2(G1348), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT60), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n1012), .A2(new_n1013), .A3(new_n592), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n591), .B1(new_n1000), .B2(KEYINPUT60), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT61), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n984), .A2(new_n990), .A3(new_n995), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1018), .B1(new_n1019), .B2(new_n997), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT58), .B(G1341), .Z(new_n1022));
  NAND2_X1  g597(.A1(new_n942), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n921), .B2(G1996), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1021), .B1(new_n1024), .B2(new_n542), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1024), .A2(new_n1021), .A3(new_n542), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1017), .B(new_n1020), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1002), .B1(new_n1010), .B2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n917), .A2(new_n718), .A3(new_n919), .A4(new_n920), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n916), .A2(new_n919), .A3(new_n911), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n718), .A2(KEYINPUT121), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n718), .A2(KEYINPUT121), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1030), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1961), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n1032), .A2(new_n1035), .B1(new_n993), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1031), .A2(G301), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1030), .A2(G2078), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n916), .A2(new_n919), .A3(new_n911), .A4(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n929), .B2(G1961), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n1030), .B2(new_n1029), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1038), .B1(new_n1042), .B2(G301), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT122), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1031), .A2(G301), .A3(new_n1037), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1032), .A2(new_n1039), .B1(new_n993), .B2(new_n1036), .ZN(new_n1049));
  AOI21_X1  g624(.A(G301), .B1(new_n1031), .B2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1047), .B(new_n1044), .C1(new_n1048), .C2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1031), .A2(new_n1037), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G171), .ZN(new_n1054));
  OAI211_X1 g629(.A(G301), .B(new_n1040), .C1(new_n929), .C2(G1961), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1044), .B1(new_n1056), .B2(new_n1031), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT123), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1054), .A2(new_n1060), .A3(new_n1057), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n1062));
  NOR3_X1   g637(.A1(G168), .A2(new_n1062), .A3(new_n944), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT120), .B1(G286), .B2(G8), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n963), .A2(new_n965), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT51), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  OR2_X1    g643(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1068), .B1(new_n966), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n967), .A2(KEYINPUT51), .A3(new_n1065), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1059), .A2(new_n1061), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1028), .A2(new_n1052), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT63), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n968), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n982), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT124), .B1(new_n979), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(new_n1069), .B2(new_n1066), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1069), .A2(new_n966), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1071), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(KEYINPUT62), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n982), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(KEYINPUT62), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n1050), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n977), .B1(new_n969), .B2(KEYINPUT63), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1075), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1051), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1047), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1054), .A2(new_n1060), .A3(new_n1057), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1060), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1081), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1088), .B1(new_n1095), .B2(new_n1028), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1086), .B(new_n1087), .C1(new_n1096), .C2(new_n982), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1077), .A2(new_n1085), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n916), .A2(new_n925), .ZN(new_n1099));
  INV_X1    g674(.A(G1996), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OR3_X1    g676(.A1(new_n1101), .A2(KEYINPUT107), .A3(new_n800), .ZN(new_n1102));
  INV_X1    g677(.A(G2067), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n742), .B(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1100), .B2(new_n801), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n1099), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT107), .B1(new_n1101), .B2(new_n800), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1102), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT108), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n754), .A2(new_n757), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n754), .A2(new_n757), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1099), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1099), .ZN(new_n1114));
  XOR2_X1   g689(.A(G290), .B(G1986), .Z(new_n1115));
  OAI21_X1  g690(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(new_n1116), .B(KEYINPUT109), .Z(new_n1117));
  NAND2_X1  g692(.A1(new_n1098), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1101), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n1119), .A2(KEYINPUT46), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(KEYINPUT46), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1114), .B1(new_n1104), .B2(new_n801), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n1123), .B(KEYINPUT47), .Z(new_n1124));
  NOR2_X1   g699(.A1(new_n742), .A2(G2067), .ZN(new_n1125));
  XOR2_X1   g700(.A(new_n1110), .B(KEYINPUT125), .Z(new_n1126));
  AOI21_X1  g701(.A(new_n1125), .B1(new_n1109), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1124), .B1(new_n1127), .B2(new_n1114), .ZN(new_n1128));
  NOR3_X1   g703(.A1(G290), .A2(G1986), .A3(new_n1114), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT48), .Z(new_n1130));
  AOI21_X1  g705(.A(new_n1128), .B1(new_n1113), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT126), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1118), .A2(new_n1132), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g708(.A1(G229), .A2(new_n459), .ZN(new_n1135));
  NAND3_X1  g709(.A1(new_n648), .A2(new_n630), .A3(new_n1135), .ZN(new_n1136));
  OR2_X1    g710(.A1(new_n1136), .A2(KEYINPUT127), .ZN(new_n1137));
  NAND2_X1  g711(.A1(new_n1136), .A2(KEYINPUT127), .ZN(new_n1138));
  NAND4_X1  g712(.A1(new_n901), .A2(new_n1137), .A3(new_n846), .A4(new_n1138), .ZN(G225));
  INV_X1    g713(.A(G225), .ZN(G308));
endmodule


