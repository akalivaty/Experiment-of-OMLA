//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1160, new_n1161, new_n1162, new_n1163, new_n1165,
    new_n1166, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT64), .B(G238), .ZN(new_n210));
  AOI21_X1  g0010(.A(new_n209), .B1(G68), .B2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AND2_X1   g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n203), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT65), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n218), .B1(new_n219), .B2(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n220), .B(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(G58), .A2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n206), .B(new_n222), .C1(new_n225), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(KEYINPUT66), .B(G264), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n232), .B(new_n233), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT67), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n235), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(KEYINPUT69), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT69), .ZN(new_n255));
  NAND2_X1  g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n254), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G222), .ZN(new_n260));
  INV_X1    g0060(.A(G223), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n258), .B(new_n260), .C1(new_n261), .C2(new_n259), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n262), .B(new_n263), .C1(G77), .C2(new_n258), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT68), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n265), .B(KEYINPUT68), .C1(G41), .C2(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n263), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G226), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n264), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G190), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT74), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n278), .B1(G200), .B2(new_n275), .ZN(new_n279));
  NAND2_X1  g0079(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n223), .ZN(new_n282));
  XOR2_X1   g0082(.A(KEYINPUT8), .B(G58), .Z(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n224), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(G20), .B1(new_n227), .B2(G50), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n282), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g0092(.A(new_n292), .B(KEYINPUT70), .Z(new_n293));
  AOI21_X1  g0093(.A(new_n282), .B1(new_n265), .B2(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G50), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n293), .B(new_n295), .C1(G50), .C2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT9), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n279), .A2(new_n280), .A3(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT75), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n299), .B(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n276), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n297), .B(new_n305), .C1(G169), .C2(new_n276), .ZN(new_n306));
  INV_X1    g0106(.A(new_n282), .ZN(new_n307));
  NAND2_X1  g0107(.A1(G58), .A2(G68), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n227), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G159), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n309), .A2(new_n224), .B1(new_n310), .B2(new_n290), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n254), .A2(new_n256), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT7), .ZN(new_n313));
  NOR3_X1   g0113(.A1(new_n312), .A2(new_n313), .A3(G20), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n249), .A2(new_n250), .ZN(new_n315));
  AOI21_X1  g0115(.A(KEYINPUT7), .B1(new_n315), .B2(new_n224), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n311), .B1(new_n317), .B2(G68), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n307), .B1(new_n318), .B2(KEYINPUT16), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT16), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n251), .A2(new_n257), .A3(new_n224), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n314), .B1(new_n313), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G68), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n320), .B1(new_n324), .B2(new_n311), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n270), .A2(G232), .ZN(new_n327));
  INV_X1    g0127(.A(G41), .ZN(new_n328));
  OAI211_X1 g0128(.A(G1), .B(G13), .C1(new_n253), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n261), .A2(new_n259), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n312), .B(new_n330), .C1(G226), .C2(new_n259), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G87), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NOR3_X1   g0133(.A1(new_n327), .A2(new_n333), .A3(new_n273), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G200), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(G190), .ZN(new_n337));
  INV_X1    g0137(.A(new_n296), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n283), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n294), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(new_n283), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n326), .A2(new_n336), .A3(new_n337), .A4(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n343), .A2(new_n344), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n334), .A2(G179), .ZN(new_n347));
  INV_X1    g0147(.A(G169), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(new_n334), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT81), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n347), .B(KEYINPUT81), .C1(new_n348), .C2(new_n334), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n326), .A2(new_n342), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n353), .A2(KEYINPUT18), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT18), .B1(new_n353), .B2(new_n354), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n345), .B(new_n346), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n210), .A2(G1698), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n258), .B(new_n359), .C1(new_n237), .C2(G1698), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(new_n263), .C1(G107), .C2(new_n258), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n270), .A2(G244), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n274), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n348), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n283), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT15), .B(G87), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT71), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n367), .B2(new_n285), .ZN(new_n368));
  INV_X1    g0168(.A(G77), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n368), .A2(new_n282), .B1(new_n369), .B2(new_n338), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(new_n369), .B2(new_n340), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n364), .A2(new_n371), .A3(KEYINPUT73), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT73), .B1(new_n364), .B2(new_n371), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n363), .A2(G179), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n303), .A2(new_n306), .A3(new_n358), .A4(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G50), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n290), .A2(new_n378), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n285), .A2(new_n369), .B1(new_n224), .B2(G68), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n282), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT11), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT79), .B1(new_n338), .B2(new_n323), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT12), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n323), .B2(new_n340), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G97), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n237), .B1(new_n251), .B2(new_n257), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(G1698), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n259), .A2(G226), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT69), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n255), .B1(new_n254), .B2(new_n256), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT76), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT76), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n258), .A2(new_n397), .A3(new_n392), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n391), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT77), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n391), .A2(new_n396), .A3(KEYINPUT77), .A4(new_n398), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n263), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n273), .B1(new_n270), .B2(G238), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT13), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT13), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n387), .B1(new_n409), .B2(G200), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(G190), .A3(new_n408), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT78), .ZN(new_n412));
  AND3_X1   g0212(.A1(new_n403), .A2(new_n407), .A3(new_n404), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT78), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(new_n416), .A3(G190), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n410), .A2(new_n412), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT14), .B1(new_n415), .B2(new_n348), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT14), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n420), .B(G169), .C1(new_n413), .C2(new_n414), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT80), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n415), .B2(G179), .ZN(new_n423));
  NOR4_X1   g0223(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT80), .A4(new_n304), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n419), .B(new_n421), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n418), .B1(new_n387), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n371), .B1(G200), .B2(new_n363), .ZN(new_n428));
  XOR2_X1   g0228(.A(new_n428), .B(KEYINPUT72), .Z(new_n429));
  INV_X1    g0229(.A(G190), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n363), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n377), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G283), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(new_n224), .C1(G33), .C2(new_n214), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n436), .B(new_n282), .C1(new_n224), .C2(G116), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT20), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n437), .B(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G116), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n338), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n307), .B(new_n296), .C1(G1), .C2(new_n253), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G116), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n439), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT88), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT88), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n439), .A2(new_n447), .A3(new_n441), .A4(new_n444), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n251), .A2(new_n257), .A3(G303), .ZN(new_n450));
  OAI211_X1 g0250(.A(G257), .B(new_n259), .C1(new_n249), .C2(new_n250), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT87), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT87), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n312), .A2(new_n453), .A3(G257), .A4(new_n259), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n312), .A2(G264), .A3(G1698), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n450), .A2(new_n452), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n263), .ZN(new_n457));
  INV_X1    g0257(.A(G45), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G1), .ZN(new_n459));
  NOR2_X1   g0259(.A1(KEYINPUT5), .A2(G41), .ZN(new_n460));
  AND2_X1   g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n459), .B(G274), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n459), .B1(new_n461), .B2(new_n460), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n329), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G270), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n457), .A2(new_n462), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n449), .B1(G190), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G200), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n467), .ZN(new_n470));
  INV_X1    g0270(.A(new_n467), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n449), .A2(G169), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT21), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n449), .A2(G179), .A3(new_n467), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n449), .A2(KEYINPUT21), .A3(G169), .A4(new_n471), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT89), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n258), .A2(new_n478), .A3(new_n224), .A4(G87), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT22), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT69), .B1(new_n480), .B2(KEYINPUT89), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n312), .A2(G87), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n224), .ZN(new_n486));
  INV_X1    g0286(.A(G107), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G20), .ZN(new_n488));
  XOR2_X1   g0288(.A(new_n488), .B(KEYINPUT23), .Z(new_n489));
  NAND3_X1  g0289(.A1(new_n481), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n490), .B(KEYINPUT24), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n282), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n443), .A2(G107), .ZN(new_n493));
  INV_X1    g0293(.A(G13), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n488), .A2(G1), .A3(new_n494), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n495), .B(KEYINPUT25), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n312), .B1(G257), .B2(new_n259), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G250), .A2(G1698), .ZN(new_n499));
  INV_X1    g0299(.A(G294), .ZN(new_n500));
  OAI22_X1  g0300(.A1(new_n498), .A2(new_n499), .B1(new_n253), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n501), .A2(new_n263), .B1(G264), .B2(new_n465), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n462), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(G179), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n504), .B1(new_n348), .B2(new_n503), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n477), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n312), .A2(G244), .A3(G1698), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT85), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n312), .A2(G238), .A3(new_n259), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n312), .A2(KEYINPUT85), .A3(G244), .A4(G1698), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n509), .A2(new_n484), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n263), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n459), .A2(G274), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n329), .B(G250), .C1(G1), .C2(new_n458), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n348), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n224), .B1(new_n388), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(G97), .A2(G107), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n212), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT86), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n518), .B1(new_n285), .B2(new_n214), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n312), .A2(new_n224), .A3(G68), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT86), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n519), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n523), .A2(new_n524), .A3(new_n525), .A4(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n528), .A2(new_n282), .B1(new_n338), .B2(new_n367), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n367), .B2(new_n442), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n517), .B(new_n530), .C1(G179), .C2(new_n516), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n516), .A2(G200), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n443), .A2(G87), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(new_n534), .C1(new_n430), .C2(new_n516), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n487), .A2(KEYINPUT6), .A3(G97), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n214), .A2(new_n487), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(new_n520), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n540), .B2(KEYINPUT6), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(G20), .B1(G77), .B2(new_n289), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n322), .B2(new_n487), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n282), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n338), .A2(G97), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n442), .B2(G97), .ZN(new_n548));
  XOR2_X1   g0348(.A(new_n548), .B(KEYINPUT83), .Z(new_n549));
  NAND3_X1  g0349(.A1(new_n543), .A2(KEYINPUT82), .A3(new_n282), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT4), .B1(new_n312), .B2(G244), .ZN(new_n552));
  INV_X1    g0352(.A(G244), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n251), .B2(new_n257), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT4), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(G1698), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n552), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n555), .B1(new_n258), .B2(G250), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n557), .B(new_n435), .C1(new_n259), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n263), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n462), .B1(new_n464), .B2(new_n215), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT84), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT84), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n563), .B(new_n462), .C1(new_n464), .C2(new_n215), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n348), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n565), .B1(new_n559), .B2(new_n263), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n304), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n551), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(new_n546), .A2(new_n550), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(G200), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n569), .A2(G190), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n572), .A2(new_n549), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n537), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n503), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G190), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n492), .A2(new_n493), .A3(new_n496), .A4(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n577), .A2(new_n469), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  AND4_X1   g0382(.A1(new_n434), .A2(new_n470), .A3(new_n506), .A4(new_n582), .ZN(G372));
  NAND2_X1  g0383(.A1(new_n346), .A2(new_n345), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n425), .A2(new_n387), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n410), .A2(new_n417), .A3(new_n412), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n375), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n584), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n354), .A2(new_n349), .ZN(new_n589));
  XOR2_X1   g0389(.A(new_n589), .B(KEYINPUT18), .Z(new_n590));
  NOR2_X1   g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n591), .B(KEYINPUT90), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n303), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n593), .A2(new_n306), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT26), .ZN(new_n595));
  OR3_X1    g0395(.A1(new_n536), .A2(new_n571), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n536), .B2(new_n571), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n492), .A2(new_n496), .ZN(new_n599));
  INV_X1    g0399(.A(new_n580), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n599), .A2(new_n493), .A3(new_n600), .A4(new_n578), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n575), .A2(new_n571), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n601), .A2(new_n602), .A3(new_n537), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n531), .B(new_n598), .C1(new_n603), .C2(new_n506), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n434), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n594), .A2(new_n605), .ZN(G369));
  NAND2_X1  g0406(.A1(new_n497), .A2(new_n505), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n265), .A2(new_n224), .A3(G13), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n608), .A2(KEYINPUT27), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(KEYINPUT27), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(G213), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(G343), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n497), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n601), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n616), .B2(new_n607), .ZN(new_n617));
  INV_X1    g0417(.A(new_n613), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n477), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(new_n607), .B2(new_n613), .ZN(new_n621));
  XNOR2_X1  g0421(.A(new_n621), .B(KEYINPUT91), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n449), .A2(new_n613), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n477), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n477), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(new_n470), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G330), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n617), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n622), .A2(new_n629), .ZN(G399));
  INV_X1    g0430(.A(new_n204), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n631), .A2(G41), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n521), .A2(G116), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G1), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n228), .B2(new_n633), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n636), .B(KEYINPUT28), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n604), .A2(new_n618), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT29), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n638), .A2(KEYINPUT94), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT94), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n604), .B2(new_n618), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n640), .B1(new_n645), .B2(new_n639), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT31), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n457), .A2(G179), .A3(new_n462), .A4(new_n466), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n516), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n560), .A2(new_n566), .A3(new_n502), .ZN(new_n650));
  OAI21_X1  g0450(.A(KEYINPUT30), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n516), .A2(new_n648), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT30), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n652), .A2(new_n569), .A3(new_n653), .A4(new_n502), .ZN(new_n654));
  NOR4_X1   g0454(.A1(new_n569), .A2(new_n577), .A3(new_n467), .A4(G179), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n651), .A2(new_n654), .B1(new_n655), .B2(new_n516), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT92), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n613), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n651), .A2(new_n654), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n655), .A2(new_n516), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n660), .A3(new_n657), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n647), .B1(new_n658), .B2(new_n662), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT93), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT93), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n582), .A2(new_n506), .A3(new_n470), .A4(new_n618), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n659), .A2(new_n660), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(KEYINPUT31), .A3(new_n613), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n664), .A2(new_n665), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n646), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n637), .B1(new_n671), .B2(G1), .ZN(G364));
  AOI21_X1  g0472(.A(new_n223), .B1(G20), .B2(new_n348), .ZN(new_n673));
  NOR2_X1   g0473(.A1(G13), .A2(G33), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G20), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n258), .A2(new_n204), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT96), .Z(new_n678));
  NAND2_X1  g0478(.A1(new_n244), .A2(G45), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n631), .A2(new_n312), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n458), .B2(new_n229), .ZN(new_n682));
  AOI22_X1  g0482(.A1(new_n678), .A2(G355), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n631), .A2(new_n440), .ZN(new_n684));
  AOI211_X1 g0484(.A(new_n673), .B(new_n676), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n494), .A2(G20), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT95), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n265), .B1(new_n687), .B2(G45), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n632), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AOI211_X1 g0491(.A(new_n685), .B(new_n691), .C1(new_n626), .C2(new_n676), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n224), .A2(new_n430), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n304), .A2(G200), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n224), .A2(G190), .ZN(new_n697));
  NOR2_X1   g0497(.A1(G179), .A2(G200), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI22_X1  g0500(.A1(G322), .A2(new_n696), .B1(new_n700), .B2(G329), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n469), .A2(G179), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n693), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G303), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n258), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n304), .A2(new_n469), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n697), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  XNOR2_X1  g0510(.A(KEYINPUT33), .B(G317), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G283), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n697), .A2(new_n702), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n707), .B(new_n712), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n708), .A2(new_n693), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  XNOR2_X1  g0517(.A(KEYINPUT97), .B(G326), .ZN(new_n718));
  AOI211_X1 g0518(.A(new_n706), .B(new_n715), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n224), .B1(new_n698), .B2(G190), .ZN(new_n720));
  INV_X1    g0520(.A(G311), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n697), .A2(new_n694), .ZN(new_n722));
  OAI221_X1 g0522(.A(new_n719), .B1(new_n500), .B2(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n720), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G97), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n212), .B2(new_n703), .ZN(new_n726));
  OAI22_X1  g0526(.A1(new_n369), .A2(new_n722), .B1(new_n714), .B2(new_n487), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n710), .A2(G68), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n699), .A2(new_n310), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT32), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n707), .B1(G58), .B2(new_n696), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n728), .A2(new_n729), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n716), .A2(new_n378), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n723), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n673), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n692), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n628), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n626), .A2(new_n627), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n738), .A2(new_n691), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n737), .A2(new_n740), .ZN(G396));
  NAND2_X1  g0541(.A1(new_n371), .A2(new_n613), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n432), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n375), .B(KEYINPUT98), .Z(new_n744));
  OAI22_X1  g0544(.A1(new_n743), .A2(new_n744), .B1(new_n376), .B2(new_n742), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n638), .B(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(new_n670), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n691), .ZN(new_n748));
  OR2_X1    g0548(.A1(new_n745), .A2(new_n675), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n673), .A2(new_n674), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n369), .ZN(new_n751));
  INV_X1    g0551(.A(G303), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n725), .B1(new_n487), .B2(new_n703), .C1(new_n752), .C2(new_n716), .ZN(new_n753));
  INV_X1    g0553(.A(new_n722), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(G116), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n714), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G87), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n700), .A2(G311), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n709), .A2(new_n713), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n258), .B(new_n759), .C1(G294), .C2(new_n696), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n755), .A2(new_n757), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(G143), .A2(new_n696), .B1(new_n754), .B2(G159), .ZN(new_n762));
  INV_X1    g0562(.A(G137), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n762), .B1(new_n763), .B2(new_n716), .C1(new_n288), .C2(new_n709), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT34), .Z(new_n765));
  AOI21_X1  g0565(.A(new_n765), .B1(G50), .B2(new_n704), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n724), .A2(G58), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n756), .A2(G68), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G132), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n312), .B1(new_n699), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n761), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n673), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n749), .A2(new_n690), .A3(new_n751), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n748), .A2(new_n774), .ZN(G384));
  INV_X1    g0575(.A(new_n387), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n618), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n585), .A2(new_n586), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT101), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n426), .A2(KEYINPUT101), .A3(new_n778), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n420), .B1(new_n409), .B2(G169), .ZN(new_n783));
  INV_X1    g0583(.A(new_n421), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(KEYINPUT80), .B1(new_n409), .B2(new_n304), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n415), .A2(new_n422), .A3(G179), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n785), .A2(new_n586), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n777), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(KEYINPUT102), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT102), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n789), .A2(new_n792), .A3(new_n777), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n781), .A2(new_n782), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n667), .A2(KEYINPUT92), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n795), .A2(KEYINPUT31), .A3(new_n613), .A4(new_n661), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT105), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n618), .B1(new_n667), .B2(KEYINPUT92), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n799), .A2(KEYINPUT105), .A3(KEYINPUT31), .A4(new_n661), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n798), .A2(new_n666), .A3(new_n663), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n745), .ZN(new_n802));
  OAI21_X1  g0602(.A(KEYINPUT106), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(KEYINPUT101), .B1(new_n426), .B2(new_n778), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n776), .B1(new_n785), .B2(new_n788), .ZN(new_n805));
  NOR4_X1   g0605(.A1(new_n805), .A2(new_n780), .A3(new_n418), .A4(new_n777), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n792), .B1(new_n789), .B2(new_n777), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n789), .A2(new_n792), .A3(new_n777), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n804), .A2(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n802), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT106), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n353), .A2(new_n354), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT104), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  INV_X1    g0616(.A(new_n611), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n354), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n343), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n353), .A2(KEYINPUT104), .A3(new_n354), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n815), .A2(new_n816), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(KEYINPUT37), .B1(new_n819), .B2(new_n589), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n590), .A2(new_n584), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n825), .B2(new_n818), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n319), .B1(KEYINPUT16), .B2(new_n318), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n342), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n349), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n817), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n831), .A2(new_n832), .A3(new_n343), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT37), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n822), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n832), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n357), .A2(KEYINPUT103), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT103), .B1(new_n357), .B2(new_n836), .ZN(new_n838));
  OAI211_X1 g0638(.A(KEYINPUT38), .B(new_n835), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n828), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n803), .A2(new_n812), .A3(KEYINPUT40), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT107), .ZN(new_n842));
  INV_X1    g0642(.A(new_n840), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n809), .A2(new_n810), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n843), .B1(new_n844), .B2(KEYINPUT106), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT40), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n781), .A2(new_n782), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n791), .A2(new_n793), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n802), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n846), .B1(new_n849), .B2(new_n811), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT107), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n845), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n842), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n835), .B1(new_n837), .B2(new_n838), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n827), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n839), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n849), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n846), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n434), .A2(new_n801), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n859), .B(new_n860), .Z(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(G330), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT39), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n840), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n855), .A2(KEYINPUT39), .A3(new_n839), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n585), .A2(new_n613), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n590), .A2(new_n611), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n744), .A2(new_n618), .ZN(new_n870));
  INV_X1    g0670(.A(new_n638), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(new_n871), .B2(new_n745), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n794), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n873), .A2(new_n856), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT108), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n434), .B(new_n640), .C1(new_n645), .C2(new_n639), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n594), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n876), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n862), .B(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n265), .B2(new_n687), .ZN(new_n881));
  OAI211_X1 g0681(.A(G116), .B(new_n225), .C1(new_n541), .C2(KEYINPUT35), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT99), .Z(new_n883));
  NAND2_X1  g0683(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT36), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n308), .A2(G77), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n228), .A2(new_n887), .B1(G50), .B2(new_n323), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(G1), .A3(new_n494), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(KEYINPUT100), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n881), .A2(new_n886), .A3(new_n890), .ZN(G367));
  AOI22_X1  g0691(.A1(G143), .A2(new_n717), .B1(new_n704), .B2(G58), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n892), .B1(new_n323), .B2(new_n720), .C1(new_n763), .C2(new_n699), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n707), .B(new_n893), .C1(G159), .C2(new_n710), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n894), .B1(new_n369), .B2(new_n714), .C1(new_n288), .C2(new_n695), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n722), .A2(new_n378), .ZN(new_n896));
  INV_X1    g0696(.A(G317), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n714), .A2(new_n214), .B1(new_n699), .B2(new_n897), .ZN(new_n898));
  OAI221_X1 g0698(.A(new_n315), .B1(new_n720), .B2(new_n487), .C1(new_n752), .C2(new_n695), .ZN(new_n899));
  AOI211_X1 g0699(.A(new_n898), .B(new_n899), .C1(G283), .C2(new_n754), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n704), .A2(G116), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT46), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n900), .B(new_n902), .C1(new_n500), .C2(new_n709), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n716), .A2(new_n721), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n895), .A2(new_n896), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT47), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n673), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n234), .A2(new_n680), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n676), .A2(new_n673), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n908), .B(new_n909), .C1(new_n204), .C2(new_n367), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n907), .A2(new_n690), .A3(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n534), .A2(new_n618), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n537), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n531), .B2(new_n912), .ZN(new_n914));
  INV_X1    g0714(.A(new_n676), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n551), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n602), .B1(new_n918), .B2(new_n618), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n571), .A2(new_n618), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR3_X1    g0721(.A1(new_n622), .A2(KEYINPUT44), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT44), .B1(new_n622), .B2(new_n921), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n622), .A2(new_n921), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT45), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT45), .B1(new_n622), .B2(new_n921), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n924), .B(new_n629), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n629), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n927), .A2(new_n928), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n922), .A2(new_n923), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n617), .B(new_n619), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(new_n628), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n671), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n929), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n671), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n632), .B(KEYINPUT41), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT110), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT110), .ZN(new_n941));
  INV_X1    g0741(.A(new_n939), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n941), .B(new_n942), .C1(new_n937), .C2(new_n671), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n688), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n617), .A2(new_n619), .A3(new_n921), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT42), .Z(new_n946));
  OAI21_X1  g0746(.A(new_n571), .B1(new_n919), .B2(new_n607), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n618), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n946), .A2(new_n948), .B1(KEYINPUT43), .B2(new_n914), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT109), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n930), .A2(new_n921), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n951), .B(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n950), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n917), .B1(new_n944), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(G387));
  NAND2_X1  g0756(.A1(new_n935), .A2(new_n689), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n681), .B1(new_n240), .B2(G45), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n323), .A2(new_n369), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT50), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n283), .A2(new_n960), .A3(new_n378), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT50), .B1(new_n284), .B2(G50), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n961), .A2(new_n458), .A3(new_n634), .A4(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n958), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n634), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n678), .A2(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n964), .B(new_n966), .C1(G107), .C2(new_n204), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n967), .A2(KEYINPUT111), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n909), .B1(new_n967), .B2(KEYINPUT111), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n690), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT112), .Z(new_n971));
  OAI22_X1  g0771(.A1(new_n714), .A2(new_n214), .B1(new_n699), .B2(new_n288), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n315), .B(new_n972), .C1(G68), .C2(new_n754), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n367), .A2(new_n720), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G159), .A2(new_n717), .B1(new_n710), .B2(new_n283), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G50), .A2(new_n696), .B1(new_n704), .B2(G77), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT113), .Z(new_n978));
  AOI22_X1  g0778(.A1(G322), .A2(new_n717), .B1(new_n710), .B2(G311), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n979), .B1(new_n752), .B2(new_n722), .C1(new_n897), .C2(new_n695), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT48), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n713), .B2(new_n720), .C1(new_n500), .C2(new_n703), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT49), .Z(new_n983));
  INV_X1    g0783(.A(new_n718), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n315), .B1(new_n714), .B2(new_n440), .C1(new_n984), .C2(new_n699), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n978), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n673), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n971), .B(new_n987), .C1(new_n617), .C2(new_n915), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n632), .B1(new_n671), .B2(new_n935), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n957), .B(new_n988), .C1(new_n936), .C2(new_n989), .ZN(G393));
  OAI221_X1 g0790(.A(new_n909), .B1(new_n214), .B2(new_n204), .C1(new_n247), .C2(new_n681), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(KEYINPUT114), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n690), .B1(new_n991), .B2(KEYINPUT114), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n716), .A2(new_n897), .B1(new_n695), .B2(new_n721), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT52), .Z(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G294), .B2(new_n754), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n703), .A2(new_n713), .B1(new_n714), .B2(new_n487), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n258), .B(new_n997), .C1(G322), .C2(new_n700), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n440), .B2(new_n720), .C1(new_n752), .C2(new_n709), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G68), .A2(new_n704), .B1(new_n754), .B2(new_n283), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n700), .A2(G143), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1001), .B(new_n1002), .C1(new_n378), .C2(new_n709), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G77), .B2(new_n724), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n716), .A2(new_n288), .B1(new_n695), .B2(new_n310), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT51), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1004), .A2(new_n312), .A3(new_n757), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1000), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n993), .B1(new_n1008), .B2(new_n673), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n992), .B(new_n1009), .C1(new_n921), .C2(new_n915), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n929), .A2(new_n933), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1010), .B1(new_n1011), .B2(new_n688), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n936), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n633), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1012), .B1(new_n1014), .B2(new_n937), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(G390));
  XOR2_X1   g0816(.A(new_n866), .B(KEYINPUT115), .Z(new_n1017));
  AOI21_X1  g0817(.A(new_n870), .B1(new_n644), .B2(new_n745), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n840), .B(new_n1017), .C1(new_n1018), .C2(new_n794), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n864), .A2(new_n865), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n873), .B2(new_n866), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n810), .A2(G330), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(new_n794), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n669), .A2(G330), .A3(new_n745), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1027), .A2(new_n794), .A3(KEYINPUT116), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT116), .B1(new_n1027), .B2(new_n794), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1019), .A2(new_n1021), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1026), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(KEYINPUT118), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n434), .A2(G330), .A3(new_n801), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n877), .A2(new_n593), .A3(new_n306), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1023), .A2(new_n794), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1030), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1018), .B(new_n1036), .C1(new_n1037), .C2(new_n1028), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n872), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1027), .A2(new_n794), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1039), .B1(new_n1024), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1035), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT118), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1026), .A2(new_n1044), .A3(new_n1031), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1033), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(KEYINPUT119), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1032), .A2(new_n1042), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(KEYINPUT117), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT117), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1032), .A2(new_n1042), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT119), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1033), .A2(new_n1043), .A3(new_n1053), .A4(new_n1045), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1047), .A2(new_n1052), .A3(new_n632), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1032), .A2(new_n689), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1020), .A2(new_n674), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n750), .A2(new_n284), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n717), .A2(G128), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n710), .A2(G137), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n258), .B1(new_n378), .B2(new_n714), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT120), .Z(new_n1062));
  NOR2_X1   g0862(.A1(new_n703), .A2(new_n288), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1063), .B(KEYINPUT53), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n700), .A2(G125), .ZN(new_n1065));
  AND4_X1   g0865(.A1(new_n1060), .A2(new_n1062), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n724), .A2(G159), .ZN(new_n1067));
  XOR2_X1   g0867(.A(KEYINPUT54), .B(G143), .Z(new_n1068));
  AOI22_X1  g0868(.A1(G132), .A2(new_n696), .B1(new_n754), .B2(new_n1068), .ZN(new_n1069));
  AND4_X1   g0869(.A1(new_n1059), .A2(new_n1066), .A3(new_n1067), .A4(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n717), .A2(G283), .B1(new_n724), .B2(G77), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1071), .B(new_n768), .C1(new_n440), .C2(new_n695), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n707), .B1(new_n212), .B2(new_n703), .C1(new_n487), .C2(new_n709), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n699), .A2(new_n500), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n722), .A2(new_n214), .ZN(new_n1075));
  NOR4_X1   g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n673), .B1(new_n1070), .B2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1057), .A2(new_n690), .A3(new_n1058), .A4(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1055), .A2(new_n1056), .A3(new_n1078), .ZN(G378));
  INV_X1    g0879(.A(new_n1035), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1051), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1050), .B1(new_n1032), .B2(new_n1042), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1080), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n841), .A2(KEYINPUT107), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n851), .B1(new_n845), .B2(new_n850), .ZN(new_n1085));
  OAI211_X1 g0885(.A(G330), .B(new_n858), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n303), .A2(new_n306), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1088));
  XNOR2_X1  g0888(.A(new_n1087), .B(new_n1088), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n297), .A2(new_n817), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1089), .B(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n853), .A2(G330), .A3(new_n858), .A4(new_n1091), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n875), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1093), .A2(new_n875), .A3(new_n1094), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1083), .B(KEYINPUT57), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1035), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1098));
  OAI21_X1  g0898(.A(KEYINPUT121), .B1(new_n1096), .B2(new_n1095), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n875), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT121), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1098), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n632), .B(new_n1097), .C1(new_n1105), .C2(KEYINPUT57), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1092), .A2(new_n674), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n750), .A2(new_n378), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n328), .B1(new_n720), .B2(new_n323), .C1(new_n369), .C2(new_n703), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(G58), .A2(new_n756), .B1(new_n700), .B2(G283), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1110), .B(new_n315), .C1(new_n214), .C2(new_n709), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(G116), .C2(new_n717), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n1112), .B1(new_n487), .B2(new_n695), .C1(new_n367), .C2(new_n722), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT58), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n378), .B1(new_n249), .B2(G41), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G128), .A2(new_n696), .B1(new_n754), .B2(G137), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n704), .A2(new_n1068), .B1(new_n724), .B2(G150), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n717), .A2(G125), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G132), .B2(new_n710), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT59), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(G41), .B1(new_n700), .B2(G124), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n253), .A3(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G159), .B2(new_n756), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n1121), .B2(new_n1120), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1114), .A2(new_n1115), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n691), .B1(new_n1127), .B2(new_n673), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1107), .A2(new_n1108), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n689), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1106), .A2(new_n1132), .ZN(G375));
  AOI21_X1  g0933(.A(new_n688), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT122), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n794), .A2(new_n674), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n750), .A2(new_n323), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n974), .B1(new_n369), .B2(new_n714), .C1(new_n500), .C2(new_n716), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n258), .B(new_n1138), .C1(G283), .C2(new_n696), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(G107), .A2(new_n754), .B1(new_n700), .B2(G303), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(new_n214), .C2(new_n703), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G116), .B2(new_n710), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n704), .A2(G159), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G132), .A2(new_n717), .B1(new_n710), .B2(new_n1068), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n763), .B2(new_n695), .ZN(new_n1145));
  OR2_X1    g0945(.A1(new_n1145), .A2(KEYINPUT123), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n315), .B1(new_n756), .B2(G58), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1145), .A2(KEYINPUT123), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(G150), .A2(new_n754), .B1(new_n724), .B2(G50), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1146), .A2(new_n1147), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G128), .B2(new_n700), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1142), .B1(new_n1143), .B2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT124), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n673), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1136), .A2(new_n690), .A3(new_n1137), .A4(new_n1154), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1135), .A2(new_n1155), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1038), .A2(new_n1035), .A3(new_n1041), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1157), .A2(new_n942), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1156), .B1(new_n1042), .B2(new_n1158), .ZN(G381));
  NAND2_X1  g0959(.A1(new_n955), .A2(new_n1015), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n1160), .A2(G396), .A3(G393), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(G375), .A2(G378), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(G381), .A2(G384), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(G407));
  INV_X1    g0964(.A(G213), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1162), .B2(new_n612), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(G407), .ZN(G409));
  INV_X1    g0967(.A(KEYINPUT61), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1165), .A2(G343), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1106), .A2(G378), .A3(new_n1132), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1093), .A2(new_n875), .A3(new_n1094), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1103), .B1(new_n1102), .B2(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1095), .A2(KEYINPUT121), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n939), .B(new_n1083), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n689), .B1(new_n1096), .B2(new_n1095), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(new_n1129), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(G378), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1169), .B1(new_n1170), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n633), .B1(new_n1157), .B2(KEYINPUT60), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n1043), .C1(KEYINPUT60), .C2(new_n1157), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1156), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1182), .A2(new_n748), .A3(new_n774), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1156), .A2(new_n1181), .A3(G384), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(G2897), .B(new_n1169), .C1(new_n1185), .C2(KEYINPUT125), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1169), .A2(G2897), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1169), .A2(KEYINPUT125), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1183), .A2(new_n1184), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1168), .B1(new_n1179), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT63), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1170), .A2(new_n1178), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1169), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1193), .B1(new_n1196), .B2(new_n1185), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1160), .A2(KEYINPUT126), .ZN(new_n1198));
  XOR2_X1   g0998(.A(G393), .B(G396), .Z(new_n1199));
  NOR2_X1   g0999(.A1(new_n955), .A2(new_n1015), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1199), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1200), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT126), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n955), .B2(new_n1015), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1202), .B1(new_n1203), .B2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1201), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1185), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1179), .A2(KEYINPUT63), .A3(new_n1208), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1192), .A2(new_n1197), .A3(new_n1207), .A4(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT62), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1179), .A2(new_n1211), .A3(new_n1208), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1179), .B2(new_n1208), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1212), .A2(new_n1191), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1210), .B1(new_n1214), .B2(new_n1207), .ZN(G405));
  NAND2_X1  g1015(.A1(G375), .A2(new_n1177), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT127), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1217), .A3(new_n1170), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(G375), .A2(KEYINPUT127), .A3(new_n1177), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1218), .A2(new_n1185), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1185), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1199), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1203), .A2(new_n1205), .A3(new_n1202), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1220), .A2(new_n1221), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1170), .A2(new_n1217), .ZN(new_n1226));
  AOI21_X1  g1026(.A(G378), .B1(new_n1106), .B2(new_n1132), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1219), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1208), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1218), .A2(new_n1185), .A3(new_n1219), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1207), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1225), .A2(new_n1232), .ZN(G402));
endmodule


