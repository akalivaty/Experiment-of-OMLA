

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U550 ( .A(n603), .B(n602), .ZN(n633) );
  NOR2_X2 U551 ( .A1(n976), .A2(n633), .ZN(n605) );
  OR2_X1 U552 ( .A1(n597), .A2(n650), .ZN(n599) );
  XNOR2_X1 U553 ( .A(n593), .B(KEYINPUT64), .ZN(n650) );
  NAND2_X1 U554 ( .A1(n793), .A2(G138), .ZN(n583) );
  INV_X1 U555 ( .A(KEYINPUT98), .ZN(n602) );
  NOR2_X1 U556 ( .A1(n650), .A2(G2084), .ZN(n651) );
  NOR2_X1 U557 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  INV_X1 U558 ( .A(KEYINPUT17), .ZN(n527) );
  NAND2_X1 U559 ( .A1(n755), .A2(n754), .ZN(n756) );
  AND2_X1 U560 ( .A1(n642), .A2(G1341), .ZN(n513) );
  NOR2_X1 U561 ( .A1(n513), .A2(n969), .ZN(n616) );
  AND2_X1 U562 ( .A1(n617), .A2(n616), .ZN(n629) );
  INV_X1 U563 ( .A(G168), .ZN(n654) );
  AND2_X1 U564 ( .A1(n655), .A2(n654), .ZN(n656) );
  AND2_X1 U565 ( .A1(n658), .A2(n657), .ZN(n660) );
  OR2_X1 U566 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U567 ( .A1(n757), .A2(G1384), .ZN(n688) );
  INV_X1 U568 ( .A(KEYINPUT87), .ZN(n582) );
  XNOR2_X1 U569 ( .A(n583), .B(n582), .ZN(n585) );
  NOR2_X1 U570 ( .A1(G651), .A2(n564), .ZN(n816) );
  AND2_X1 U571 ( .A1(n532), .A2(G2104), .ZN(n794) );
  NOR2_X1 U572 ( .A1(G651), .A2(G543), .ZN(n810) );
  NOR2_X1 U573 ( .A1(n536), .A2(n535), .ZN(G160) );
  NAND2_X1 U574 ( .A1(G89), .A2(n810), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n514), .B(KEYINPUT4), .ZN(n515) );
  XNOR2_X1 U576 ( .A(n515), .B(KEYINPUT72), .ZN(n517) );
  XOR2_X1 U577 ( .A(KEYINPUT0), .B(G543), .Z(n564) );
  INV_X1 U578 ( .A(G651), .ZN(n519) );
  NOR2_X1 U579 ( .A1(n564), .A2(n519), .ZN(n815) );
  NAND2_X1 U580 ( .A1(G76), .A2(n815), .ZN(n516) );
  NAND2_X1 U581 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(KEYINPUT5), .ZN(n525) );
  NOR2_X1 U583 ( .A1(G543), .A2(n519), .ZN(n520) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n520), .Z(n812) );
  NAND2_X1 U585 ( .A1(G63), .A2(n812), .ZN(n522) );
  NAND2_X1 U586 ( .A1(G51), .A2(n816), .ZN(n521) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U588 ( .A(KEYINPUT6), .B(n523), .Z(n524) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X2 U591 ( .A(n528), .B(n527), .ZN(n793) );
  NAND2_X1 U592 ( .A1(n793), .A2(G137), .ZN(n531) );
  INV_X1 U593 ( .A(G2105), .ZN(n532) );
  NAND2_X1 U594 ( .A1(G101), .A2(n794), .ZN(n529) );
  XOR2_X1 U595 ( .A(KEYINPUT23), .B(n529), .Z(n530) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n536) );
  AND2_X1 U597 ( .A1(G2105), .A2(G2104), .ZN(n798) );
  NAND2_X1 U598 ( .A1(G113), .A2(n798), .ZN(n534) );
  NOR2_X1 U599 ( .A1(G2104), .A2(n532), .ZN(n799) );
  NAND2_X1 U600 ( .A1(G125), .A2(n799), .ZN(n533) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U602 ( .A1(G64), .A2(n812), .ZN(n538) );
  NAND2_X1 U603 ( .A1(G52), .A2(n816), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n544) );
  NAND2_X1 U605 ( .A1(n815), .A2(G77), .ZN(n539) );
  XNOR2_X1 U606 ( .A(n539), .B(KEYINPUT66), .ZN(n541) );
  NAND2_X1 U607 ( .A1(G90), .A2(n810), .ZN(n540) );
  NAND2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U609 ( .A(KEYINPUT9), .B(n542), .Z(n543) );
  NOR2_X1 U610 ( .A1(n544), .A2(n543), .ZN(G171) );
  NAND2_X1 U611 ( .A1(G65), .A2(n812), .ZN(n546) );
  NAND2_X1 U612 ( .A1(G53), .A2(n816), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(KEYINPUT67), .B(n547), .ZN(n551) );
  NAND2_X1 U615 ( .A1(n815), .A2(G78), .ZN(n549) );
  NAND2_X1 U616 ( .A1(G91), .A2(n810), .ZN(n548) );
  AND2_X1 U617 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(G299) );
  NAND2_X1 U619 ( .A1(G75), .A2(n815), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(KEYINPUT80), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G62), .A2(n812), .ZN(n554) );
  NAND2_X1 U622 ( .A1(G50), .A2(n816), .ZN(n553) );
  NAND2_X1 U623 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U624 ( .A(KEYINPUT78), .B(n555), .ZN(n558) );
  NAND2_X1 U625 ( .A1(G88), .A2(n810), .ZN(n556) );
  XNOR2_X1 U626 ( .A(KEYINPUT79), .B(n556), .ZN(n557) );
  NOR2_X1 U627 ( .A1(n558), .A2(n557), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(G303) );
  XOR2_X1 U629 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U630 ( .A1(G49), .A2(n816), .ZN(n562) );
  NAND2_X1 U631 ( .A1(G74), .A2(G651), .ZN(n561) );
  NAND2_X1 U632 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U633 ( .A1(n812), .A2(n563), .ZN(n567) );
  NAND2_X1 U634 ( .A1(G87), .A2(n564), .ZN(n565) );
  XOR2_X1 U635 ( .A(KEYINPUT77), .B(n565), .Z(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(G288) );
  NAND2_X1 U637 ( .A1(G61), .A2(n812), .ZN(n569) );
  NAND2_X1 U638 ( .A1(G48), .A2(n816), .ZN(n568) );
  NAND2_X1 U639 ( .A1(n569), .A2(n568), .ZN(n572) );
  NAND2_X1 U640 ( .A1(G73), .A2(n815), .ZN(n570) );
  XOR2_X1 U641 ( .A(KEYINPUT2), .B(n570), .Z(n571) );
  NOR2_X1 U642 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n810), .A2(G86), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(G305) );
  NAND2_X1 U645 ( .A1(G72), .A2(n815), .ZN(n576) );
  NAND2_X1 U646 ( .A1(G85), .A2(n810), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U648 ( .A(KEYINPUT65), .B(n577), .ZN(n581) );
  NAND2_X1 U649 ( .A1(G60), .A2(n812), .ZN(n579) );
  NAND2_X1 U650 ( .A1(G47), .A2(n816), .ZN(n578) );
  AND2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U652 ( .A1(n581), .A2(n580), .ZN(G290) );
  INV_X1 U653 ( .A(G303), .ZN(G166) );
  NAND2_X1 U654 ( .A1(G160), .A2(G40), .ZN(n687) );
  INV_X1 U655 ( .A(n687), .ZN(n592) );
  NAND2_X1 U656 ( .A1(n794), .A2(G102), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U658 ( .A(n586), .B(KEYINPUT88), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n798), .A2(G114), .ZN(n587) );
  XNOR2_X1 U660 ( .A(n587), .B(KEYINPUT86), .ZN(n589) );
  NAND2_X1 U661 ( .A1(G126), .A2(n799), .ZN(n588) );
  NAND2_X1 U662 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U663 ( .A1(n591), .A2(n590), .ZN(n757) );
  NAND2_X1 U664 ( .A1(n592), .A2(n688), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n650), .A2(G8), .ZN(n730) );
  BUF_X2 U666 ( .A(n650), .Z(n642) );
  INV_X1 U667 ( .A(n642), .ZN(n625) );
  NOR2_X1 U668 ( .A1(G1961), .A2(n625), .ZN(n595) );
  XOR2_X1 U669 ( .A(KEYINPUT25), .B(G2078), .Z(n952) );
  NOR2_X1 U670 ( .A1(n642), .A2(n952), .ZN(n594) );
  NOR2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U672 ( .A(n596), .B(KEYINPUT97), .ZN(n648) );
  NAND2_X1 U673 ( .A1(n648), .A2(G171), .ZN(n640) );
  INV_X1 U674 ( .A(G299), .ZN(n976) );
  INV_X1 U675 ( .A(G2072), .ZN(n597) );
  INV_X1 U676 ( .A(KEYINPUT27), .ZN(n598) );
  XNOR2_X1 U677 ( .A(n599), .B(n598), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n642), .A2(G1956), .ZN(n600) );
  NAND2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n603) );
  INV_X1 U680 ( .A(KEYINPUT28), .ZN(n604) );
  XNOR2_X1 U681 ( .A(n605), .B(n604), .ZN(n637) );
  NAND2_X1 U682 ( .A1(n625), .A2(G1996), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n606), .B(KEYINPUT26), .ZN(n617) );
  NAND2_X1 U684 ( .A1(G56), .A2(n812), .ZN(n607) );
  XOR2_X1 U685 ( .A(KEYINPUT14), .B(n607), .Z(n613) );
  NAND2_X1 U686 ( .A1(n810), .A2(G81), .ZN(n608) );
  XNOR2_X1 U687 ( .A(n608), .B(KEYINPUT12), .ZN(n610) );
  NAND2_X1 U688 ( .A1(G68), .A2(n815), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U690 ( .A(KEYINPUT13), .B(n611), .Z(n612) );
  NOR2_X1 U691 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n816), .A2(G43), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n969) );
  NAND2_X1 U694 ( .A1(G79), .A2(n815), .ZN(n619) );
  NAND2_X1 U695 ( .A1(G54), .A2(n816), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U697 ( .A1(G66), .A2(n812), .ZN(n621) );
  NAND2_X1 U698 ( .A1(G92), .A2(n810), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U701 ( .A(n624), .B(KEYINPUT15), .ZN(n979) );
  NAND2_X1 U702 ( .A1(G2067), .A2(n625), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n642), .A2(G1348), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n630) );
  NOR2_X1 U705 ( .A1(n979), .A2(n630), .ZN(n628) );
  OR2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n979), .A2(n630), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U709 ( .A1(n976), .A2(n633), .ZN(n634) );
  NAND2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U712 ( .A(n638), .B(KEYINPUT29), .Z(n639) );
  NAND2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n668) );
  INV_X1 U714 ( .A(G8), .ZN(n647) );
  NOR2_X1 U715 ( .A1(G1971), .A2(n730), .ZN(n641) );
  XOR2_X1 U716 ( .A(KEYINPUT101), .B(n641), .Z(n644) );
  NOR2_X1 U717 ( .A1(n642), .A2(G2090), .ZN(n643) );
  NOR2_X1 U718 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n645), .A2(G303), .ZN(n646) );
  OR2_X1 U720 ( .A1(n647), .A2(n646), .ZN(n662) );
  AND2_X1 U721 ( .A1(n668), .A2(n662), .ZN(n661) );
  NOR2_X1 U722 ( .A1(G171), .A2(n648), .ZN(n649) );
  XOR2_X1 U723 ( .A(KEYINPUT100), .B(n649), .Z(n658) );
  NOR2_X1 U724 ( .A1(G1966), .A2(n730), .ZN(n671) );
  XOR2_X1 U725 ( .A(KEYINPUT96), .B(n651), .Z(n669) );
  NAND2_X1 U726 ( .A1(G8), .A2(n669), .ZN(n652) );
  NOR2_X1 U727 ( .A1(n671), .A2(n652), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n653), .B(KEYINPUT30), .ZN(n655) );
  XNOR2_X1 U729 ( .A(KEYINPUT99), .B(n656), .ZN(n657) );
  INV_X1 U730 ( .A(KEYINPUT31), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n660), .B(n659), .ZN(n667) );
  NAND2_X1 U732 ( .A1(n661), .A2(n667), .ZN(n665) );
  INV_X1 U733 ( .A(n662), .ZN(n663) );
  OR2_X1 U734 ( .A1(n663), .A2(G286), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n666), .B(KEYINPUT32), .ZN(n676) );
  AND2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n674) );
  INV_X1 U738 ( .A(n669), .ZN(n670) );
  AND2_X1 U739 ( .A1(n670), .A2(G8), .ZN(n672) );
  OR2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n731) );
  NOR2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n685) );
  NOR2_X1 U743 ( .A1(G1971), .A2(G303), .ZN(n677) );
  NOR2_X1 U744 ( .A1(n685), .A2(n677), .ZN(n973) );
  XNOR2_X1 U745 ( .A(KEYINPUT102), .B(n973), .ZN(n678) );
  NAND2_X1 U746 ( .A1(n731), .A2(n678), .ZN(n679) );
  NAND2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n982) );
  NAND2_X1 U748 ( .A1(n679), .A2(n982), .ZN(n680) );
  XOR2_X1 U749 ( .A(KEYINPUT103), .B(n680), .Z(n681) );
  NOR2_X1 U750 ( .A1(n730), .A2(n681), .ZN(n682) );
  NOR2_X1 U751 ( .A1(KEYINPUT33), .A2(n682), .ZN(n684) );
  INV_X1 U752 ( .A(KEYINPUT104), .ZN(n683) );
  XNOR2_X1 U753 ( .A(n684), .B(n683), .ZN(n724) );
  NAND2_X1 U754 ( .A1(n685), .A2(KEYINPUT33), .ZN(n686) );
  NOR2_X1 U755 ( .A1(n730), .A2(n686), .ZN(n722) );
  XOR2_X1 U756 ( .A(G1981), .B(G305), .Z(n984) );
  NOR2_X1 U757 ( .A1(n688), .A2(n687), .ZN(n750) );
  NAND2_X1 U758 ( .A1(G140), .A2(n793), .ZN(n690) );
  NAND2_X1 U759 ( .A1(G104), .A2(n794), .ZN(n689) );
  NAND2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  XNOR2_X1 U761 ( .A(KEYINPUT34), .B(n691), .ZN(n696) );
  NAND2_X1 U762 ( .A1(G116), .A2(n798), .ZN(n693) );
  NAND2_X1 U763 ( .A1(G128), .A2(n799), .ZN(n692) );
  NAND2_X1 U764 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U765 ( .A(n694), .B(KEYINPUT35), .Z(n695) );
  NOR2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U767 ( .A(KEYINPUT36), .B(n697), .Z(n698) );
  XNOR2_X1 U768 ( .A(KEYINPUT91), .B(n698), .ZN(n807) );
  XNOR2_X1 U769 ( .A(G2067), .B(KEYINPUT37), .ZN(n747) );
  NOR2_X1 U770 ( .A1(n807), .A2(n747), .ZN(n699) );
  XNOR2_X1 U771 ( .A(n699), .B(KEYINPUT92), .ZN(n932) );
  NAND2_X1 U772 ( .A1(n750), .A2(n932), .ZN(n745) );
  XOR2_X1 U773 ( .A(KEYINPUT89), .B(G1986), .Z(n700) );
  XNOR2_X1 U774 ( .A(G290), .B(n700), .ZN(n971) );
  NAND2_X1 U775 ( .A1(n971), .A2(n750), .ZN(n701) );
  XNOR2_X1 U776 ( .A(n701), .B(KEYINPUT90), .ZN(n718) );
  NAND2_X1 U777 ( .A1(G117), .A2(n798), .ZN(n703) );
  NAND2_X1 U778 ( .A1(G141), .A2(n793), .ZN(n702) );
  NAND2_X1 U779 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U780 ( .A1(n794), .A2(G105), .ZN(n704) );
  XOR2_X1 U781 ( .A(KEYINPUT38), .B(n704), .Z(n705) );
  NOR2_X1 U782 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U783 ( .A1(n799), .A2(G129), .ZN(n707) );
  NAND2_X1 U784 ( .A1(n708), .A2(n707), .ZN(n780) );
  NAND2_X1 U785 ( .A1(G1996), .A2(n780), .ZN(n716) );
  NAND2_X1 U786 ( .A1(G107), .A2(n798), .ZN(n710) );
  NAND2_X1 U787 ( .A1(G131), .A2(n793), .ZN(n709) );
  NAND2_X1 U788 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U789 ( .A1(G119), .A2(n799), .ZN(n712) );
  NAND2_X1 U790 ( .A1(G95), .A2(n794), .ZN(n711) );
  NAND2_X1 U791 ( .A1(n712), .A2(n711), .ZN(n713) );
  OR2_X1 U792 ( .A1(n714), .A2(n713), .ZN(n785) );
  NAND2_X1 U793 ( .A1(G1991), .A2(n785), .ZN(n715) );
  NAND2_X1 U794 ( .A1(n716), .A2(n715), .ZN(n928) );
  NAND2_X1 U795 ( .A1(n928), .A2(n750), .ZN(n717) );
  AND2_X1 U796 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U797 ( .A1(n745), .A2(n719), .ZN(n740) );
  INV_X1 U798 ( .A(n740), .ZN(n720) );
  NAND2_X1 U799 ( .A1(n984), .A2(n720), .ZN(n721) );
  NOR2_X1 U800 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U801 ( .A1(n724), .A2(n723), .ZN(n755) );
  NOR2_X1 U802 ( .A1(G1981), .A2(G305), .ZN(n727) );
  XNOR2_X1 U803 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n725) );
  XNOR2_X1 U804 ( .A(n725), .B(KEYINPUT24), .ZN(n726) );
  XNOR2_X1 U805 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U806 ( .A1(n730), .A2(n728), .ZN(n729) );
  XOR2_X1 U807 ( .A(KEYINPUT95), .B(n729), .Z(n738) );
  INV_X1 U808 ( .A(n730), .ZN(n736) );
  INV_X1 U809 ( .A(n731), .ZN(n734) );
  NAND2_X1 U810 ( .A1(G8), .A2(G166), .ZN(n732) );
  NOR2_X1 U811 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U812 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U813 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U814 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U815 ( .A1(n740), .A2(n739), .ZN(n753) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n780), .ZN(n921) );
  NOR2_X1 U817 ( .A1(G1986), .A2(G290), .ZN(n741) );
  NOR2_X1 U818 ( .A1(G1991), .A2(n785), .ZN(n924) );
  NOR2_X1 U819 ( .A1(n741), .A2(n924), .ZN(n742) );
  NOR2_X1 U820 ( .A1(n928), .A2(n742), .ZN(n743) );
  NOR2_X1 U821 ( .A1(n921), .A2(n743), .ZN(n744) );
  XNOR2_X1 U822 ( .A(KEYINPUT39), .B(n744), .ZN(n746) );
  NAND2_X1 U823 ( .A1(n746), .A2(n745), .ZN(n748) );
  NAND2_X1 U824 ( .A1(n747), .A2(n807), .ZN(n934) );
  NAND2_X1 U825 ( .A1(n748), .A2(n934), .ZN(n749) );
  NAND2_X1 U826 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U827 ( .A(n751), .B(KEYINPUT105), .ZN(n752) );
  NOR2_X1 U828 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U829 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  BUF_X1 U830 ( .A(n757), .Z(G164) );
  NAND2_X1 U831 ( .A1(G124), .A2(n799), .ZN(n758) );
  XOR2_X1 U832 ( .A(KEYINPUT115), .B(n758), .Z(n759) );
  XNOR2_X1 U833 ( .A(n759), .B(KEYINPUT44), .ZN(n761) );
  NAND2_X1 U834 ( .A1(G112), .A2(n798), .ZN(n760) );
  NAND2_X1 U835 ( .A1(n761), .A2(n760), .ZN(n765) );
  NAND2_X1 U836 ( .A1(G136), .A2(n793), .ZN(n763) );
  NAND2_X1 U837 ( .A1(G100), .A2(n794), .ZN(n762) );
  NAND2_X1 U838 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U839 ( .A1(n765), .A2(n764), .ZN(G162) );
  NAND2_X1 U840 ( .A1(G111), .A2(n798), .ZN(n767) );
  NAND2_X1 U841 ( .A1(G135), .A2(n793), .ZN(n766) );
  NAND2_X1 U842 ( .A1(n767), .A2(n766), .ZN(n770) );
  NAND2_X1 U843 ( .A1(n799), .A2(G123), .ZN(n768) );
  XOR2_X1 U844 ( .A(KEYINPUT18), .B(n768), .Z(n769) );
  NOR2_X1 U845 ( .A1(n770), .A2(n769), .ZN(n772) );
  NAND2_X1 U846 ( .A1(n794), .A2(G99), .ZN(n771) );
  NAND2_X1 U847 ( .A1(n772), .A2(n771), .ZN(n925) );
  NAND2_X1 U848 ( .A1(G118), .A2(n798), .ZN(n774) );
  NAND2_X1 U849 ( .A1(G130), .A2(n799), .ZN(n773) );
  NAND2_X1 U850 ( .A1(n774), .A2(n773), .ZN(n779) );
  NAND2_X1 U851 ( .A1(G142), .A2(n793), .ZN(n776) );
  NAND2_X1 U852 ( .A1(G106), .A2(n794), .ZN(n775) );
  NAND2_X1 U853 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U854 ( .A(n777), .B(KEYINPUT45), .Z(n778) );
  NOR2_X1 U855 ( .A1(n779), .A2(n778), .ZN(n781) );
  XNOR2_X1 U856 ( .A(n781), .B(n780), .ZN(n789) );
  XOR2_X1 U857 ( .A(KEYINPUT117), .B(KEYINPUT48), .Z(n783) );
  XNOR2_X1 U858 ( .A(KEYINPUT120), .B(KEYINPUT119), .ZN(n782) );
  XNOR2_X1 U859 ( .A(n783), .B(n782), .ZN(n784) );
  XNOR2_X1 U860 ( .A(KEYINPUT116), .B(n784), .ZN(n787) );
  XNOR2_X1 U861 ( .A(n785), .B(KEYINPUT46), .ZN(n786) );
  XNOR2_X1 U862 ( .A(n787), .B(n786), .ZN(n788) );
  XOR2_X1 U863 ( .A(n789), .B(n788), .Z(n791) );
  XNOR2_X1 U864 ( .A(G164), .B(G162), .ZN(n790) );
  XNOR2_X1 U865 ( .A(n791), .B(n790), .ZN(n792) );
  XNOR2_X1 U866 ( .A(n925), .B(n792), .ZN(n806) );
  NAND2_X1 U867 ( .A1(G139), .A2(n793), .ZN(n796) );
  NAND2_X1 U868 ( .A1(G103), .A2(n794), .ZN(n795) );
  NAND2_X1 U869 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U870 ( .A(KEYINPUT118), .B(n797), .ZN(n804) );
  NAND2_X1 U871 ( .A1(G115), .A2(n798), .ZN(n801) );
  NAND2_X1 U872 ( .A1(G127), .A2(n799), .ZN(n800) );
  NAND2_X1 U873 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U874 ( .A(KEYINPUT47), .B(n802), .Z(n803) );
  NOR2_X1 U875 ( .A1(n804), .A2(n803), .ZN(n937) );
  XNOR2_X1 U876 ( .A(G160), .B(n937), .ZN(n805) );
  XNOR2_X1 U877 ( .A(n806), .B(n805), .ZN(n808) );
  XOR2_X1 U878 ( .A(n808), .B(n807), .Z(n809) );
  NOR2_X1 U879 ( .A1(G37), .A2(n809), .ZN(G395) );
  XNOR2_X1 U880 ( .A(G286), .B(n979), .ZN(n829) );
  NAND2_X1 U881 ( .A1(G93), .A2(n810), .ZN(n811) );
  XNOR2_X1 U882 ( .A(n811), .B(KEYINPUT76), .ZN(n814) );
  NAND2_X1 U883 ( .A1(n812), .A2(G67), .ZN(n813) );
  NAND2_X1 U884 ( .A1(n814), .A2(n813), .ZN(n820) );
  NAND2_X1 U885 ( .A1(G80), .A2(n815), .ZN(n818) );
  NAND2_X1 U886 ( .A1(G55), .A2(n816), .ZN(n817) );
  NAND2_X1 U887 ( .A1(n818), .A2(n817), .ZN(n819) );
  OR2_X1 U888 ( .A1(n820), .A2(n819), .ZN(n902) );
  XNOR2_X1 U889 ( .A(KEYINPUT19), .B(KEYINPUT82), .ZN(n822) );
  XNOR2_X1 U890 ( .A(G290), .B(KEYINPUT81), .ZN(n821) );
  XNOR2_X1 U891 ( .A(n822), .B(n821), .ZN(n823) );
  XNOR2_X1 U892 ( .A(G166), .B(n823), .ZN(n825) );
  XNOR2_X1 U893 ( .A(G288), .B(n976), .ZN(n824) );
  XNOR2_X1 U894 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U895 ( .A(n902), .B(n826), .Z(n827) );
  XNOR2_X1 U896 ( .A(n827), .B(G305), .ZN(n828) );
  XNOR2_X1 U897 ( .A(n969), .B(n828), .ZN(n899) );
  XNOR2_X1 U898 ( .A(n829), .B(n899), .ZN(n830) );
  XOR2_X1 U899 ( .A(G171), .B(n830), .Z(n831) );
  NOR2_X1 U900 ( .A1(G37), .A2(n831), .ZN(G397) );
  XOR2_X1 U901 ( .A(G2096), .B(KEYINPUT43), .Z(n833) );
  XNOR2_X1 U902 ( .A(G2090), .B(KEYINPUT42), .ZN(n832) );
  XNOR2_X1 U903 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U904 ( .A(n834), .B(G2678), .Z(n836) );
  XNOR2_X1 U905 ( .A(G2067), .B(G2072), .ZN(n835) );
  XNOR2_X1 U906 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U907 ( .A(KEYINPUT112), .B(G2100), .Z(n838) );
  XNOR2_X1 U908 ( .A(G2078), .B(G2084), .ZN(n837) );
  XNOR2_X1 U909 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U910 ( .A(n840), .B(n839), .ZN(G227) );
  XOR2_X1 U911 ( .A(KEYINPUT114), .B(G1961), .Z(n842) );
  XNOR2_X1 U912 ( .A(G1981), .B(G1966), .ZN(n841) );
  XNOR2_X1 U913 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U914 ( .A(n843), .B(KEYINPUT41), .Z(n845) );
  XNOR2_X1 U915 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U916 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U917 ( .A(G1986), .B(G1971), .Z(n847) );
  XNOR2_X1 U918 ( .A(G1976), .B(G1956), .ZN(n846) );
  XNOR2_X1 U919 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U920 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U921 ( .A(KEYINPUT113), .B(G2474), .ZN(n850) );
  XNOR2_X1 U922 ( .A(n851), .B(n850), .ZN(G229) );
  XNOR2_X1 U923 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U924 ( .A(G57), .ZN(G237) );
  XOR2_X1 U925 ( .A(KEYINPUT83), .B(KEYINPUT22), .Z(n853) );
  NAND2_X1 U926 ( .A1(G132), .A2(G82), .ZN(n852) );
  XNOR2_X1 U927 ( .A(n853), .B(n852), .ZN(n854) );
  NOR2_X1 U928 ( .A1(n854), .A2(G218), .ZN(n855) );
  NAND2_X1 U929 ( .A1(G96), .A2(n855), .ZN(n918) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n918), .ZN(n859) );
  NAND2_X1 U931 ( .A1(G69), .A2(G120), .ZN(n856) );
  NOR2_X1 U932 ( .A1(G237), .A2(n856), .ZN(n857) );
  NAND2_X1 U933 ( .A1(G108), .A2(n857), .ZN(n919) );
  NAND2_X1 U934 ( .A1(G567), .A2(n919), .ZN(n858) );
  NAND2_X1 U935 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U936 ( .A(KEYINPUT84), .B(n860), .ZN(n911) );
  XNOR2_X1 U937 ( .A(KEYINPUT111), .B(n911), .ZN(G319) );
  XNOR2_X1 U938 ( .A(G2443), .B(G2454), .ZN(n870) );
  XOR2_X1 U939 ( .A(G2430), .B(KEYINPUT106), .Z(n862) );
  XNOR2_X1 U940 ( .A(G2446), .B(KEYINPUT107), .ZN(n861) );
  XNOR2_X1 U941 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U942 ( .A(G2451), .B(G2427), .Z(n864) );
  XNOR2_X1 U943 ( .A(G1341), .B(G1348), .ZN(n863) );
  XNOR2_X1 U944 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U945 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U946 ( .A(G2438), .B(G2435), .ZN(n867) );
  XNOR2_X1 U947 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U948 ( .A(n870), .B(n869), .ZN(n871) );
  NAND2_X1 U949 ( .A1(n871), .A2(G14), .ZN(n912) );
  NOR2_X1 U950 ( .A1(G227), .A2(G229), .ZN(n872) );
  XOR2_X1 U951 ( .A(KEYINPUT49), .B(n872), .Z(n873) );
  NAND2_X1 U952 ( .A1(n912), .A2(n873), .ZN(n874) );
  NOR2_X1 U953 ( .A1(G397), .A2(n874), .ZN(n875) );
  NAND2_X1 U954 ( .A1(n875), .A2(G319), .ZN(n876) );
  OR2_X1 U955 ( .A1(G395), .A2(n876), .ZN(G225) );
  AND2_X1 U956 ( .A1(G452), .A2(G94), .ZN(G173) );
  XNOR2_X1 U957 ( .A(G2096), .B(n925), .ZN(n877) );
  OR2_X1 U958 ( .A1(G2100), .A2(n877), .ZN(G156) );
  NAND2_X1 U959 ( .A1(G7), .A2(G661), .ZN(n878) );
  XNOR2_X1 U960 ( .A(n878), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U961 ( .A(G223), .B(KEYINPUT68), .Z(n913) );
  NAND2_X1 U962 ( .A1(n913), .A2(G567), .ZN(n879) );
  XOR2_X1 U963 ( .A(KEYINPUT11), .B(n879), .Z(G234) );
  INV_X1 U964 ( .A(G860), .ZN(n886) );
  OR2_X1 U965 ( .A1(n969), .A2(n886), .ZN(n880) );
  XOR2_X1 U966 ( .A(KEYINPUT69), .B(n880), .Z(G153) );
  XOR2_X1 U967 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  INV_X1 U968 ( .A(G868), .ZN(n901) );
  NOR2_X1 U969 ( .A1(G301), .A2(n901), .ZN(n882) );
  NOR2_X1 U970 ( .A1(G868), .A2(n979), .ZN(n881) );
  NOR2_X1 U971 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U972 ( .A(KEYINPUT71), .B(n883), .Z(G284) );
  NOR2_X1 U973 ( .A1(G286), .A2(n901), .ZN(n885) );
  NOR2_X1 U974 ( .A1(G868), .A2(G299), .ZN(n884) );
  NOR2_X1 U975 ( .A1(n885), .A2(n884), .ZN(G297) );
  NAND2_X1 U976 ( .A1(n886), .A2(G559), .ZN(n887) );
  INV_X1 U977 ( .A(n979), .ZN(n895) );
  NAND2_X1 U978 ( .A1(n887), .A2(n895), .ZN(n888) );
  XNOR2_X1 U979 ( .A(n888), .B(KEYINPUT16), .ZN(n889) );
  XOR2_X1 U980 ( .A(KEYINPUT73), .B(n889), .Z(G148) );
  NAND2_X1 U981 ( .A1(n895), .A2(G868), .ZN(n890) );
  NOR2_X1 U982 ( .A1(G559), .A2(n890), .ZN(n891) );
  XOR2_X1 U983 ( .A(KEYINPUT75), .B(n891), .Z(n894) );
  NOR2_X1 U984 ( .A1(G868), .A2(n969), .ZN(n892) );
  XNOR2_X1 U985 ( .A(KEYINPUT74), .B(n892), .ZN(n893) );
  NOR2_X1 U986 ( .A1(n894), .A2(n893), .ZN(G282) );
  NAND2_X1 U987 ( .A1(n895), .A2(G559), .ZN(n898) );
  XNOR2_X1 U988 ( .A(n969), .B(n898), .ZN(n896) );
  NOR2_X1 U989 ( .A1(n896), .A2(G860), .ZN(n897) );
  XOR2_X1 U990 ( .A(n897), .B(n902), .Z(G145) );
  XOR2_X1 U991 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U992 ( .A1(n901), .A2(n900), .ZN(n904) );
  NOR2_X1 U993 ( .A1(G868), .A2(n902), .ZN(n903) );
  NOR2_X1 U994 ( .A1(n904), .A2(n903), .ZN(G295) );
  NAND2_X1 U995 ( .A1(G2078), .A2(G2084), .ZN(n905) );
  XOR2_X1 U996 ( .A(KEYINPUT20), .B(n905), .Z(n906) );
  NAND2_X1 U997 ( .A1(G2090), .A2(n906), .ZN(n907) );
  XNOR2_X1 U998 ( .A(KEYINPUT21), .B(n907), .ZN(n908) );
  NAND2_X1 U999 ( .A1(n908), .A2(G2072), .ZN(G158) );
  NAND2_X1 U1000 ( .A1(G661), .A2(G483), .ZN(n909) );
  XOR2_X1 U1001 ( .A(KEYINPUT85), .B(n909), .Z(n910) );
  NOR2_X1 U1002 ( .A1(n911), .A2(n910), .ZN(n917) );
  NAND2_X1 U1003 ( .A1(n917), .A2(G36), .ZN(G176) );
  XOR2_X1 U1004 ( .A(KEYINPUT108), .B(n912), .Z(G401) );
  NAND2_X1 U1005 ( .A1(G2106), .A2(n913), .ZN(G217) );
  AND2_X1 U1006 ( .A1(G15), .A2(G2), .ZN(n914) );
  NAND2_X1 U1007 ( .A1(G661), .A2(n914), .ZN(G259) );
  NAND2_X1 U1008 ( .A1(G3), .A2(G1), .ZN(n915) );
  XOR2_X1 U1009 ( .A(KEYINPUT109), .B(n915), .Z(n916) );
  NAND2_X1 U1010 ( .A1(n917), .A2(n916), .ZN(G188) );
  NOR2_X1 U1011 ( .A1(n919), .A2(n918), .ZN(G325) );
  XOR2_X1 U1012 ( .A(KEYINPUT110), .B(G325), .Z(G261) );
  XNOR2_X1 U1013 ( .A(KEYINPUT121), .B(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G132), .ZN(G219) );
  INV_X1 U1016 ( .A(G120), .ZN(G236) );
  INV_X1 U1017 ( .A(G96), .ZN(G221) );
  INV_X1 U1018 ( .A(G82), .ZN(G220) );
  INV_X1 U1019 ( .A(G69), .ZN(G235) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n920) );
  NOR2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n922) );
  XOR2_X1 U1023 ( .A(KEYINPUT51), .B(n922), .Z(n930) );
  XOR2_X1 U1024 ( .A(G2084), .B(G160), .Z(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(n933), .B(KEYINPUT122), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n943) );
  XNOR2_X1 U1032 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n936) );
  XNOR2_X1 U1033 ( .A(n936), .B(KEYINPUT50), .ZN(n941) );
  XOR2_X1 U1034 ( .A(G2072), .B(n937), .Z(n939) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1037 ( .A(n941), .B(n940), .ZN(n942) );
  NOR2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(KEYINPUT52), .B(n944), .ZN(n945) );
  INV_X1 U1040 ( .A(KEYINPUT55), .ZN(n965) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n965), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n946), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1043 ( .A(KEYINPUT125), .B(G2090), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(n947), .B(G35), .ZN(n963) );
  XNOR2_X1 U1045 ( .A(G2084), .B(G34), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(n948), .B(KEYINPUT54), .ZN(n961) );
  XOR2_X1 U1047 ( .A(G1991), .B(G25), .Z(n949) );
  NAND2_X1 U1048 ( .A1(n949), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(G1996), .B(G32), .ZN(n951) );
  XNOR2_X1 U1050 ( .A(G33), .B(G2072), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n954) );
  XNOR2_X1 U1053 ( .A(G27), .B(n952), .ZN(n953) );
  NOR2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(n959), .B(KEYINPUT53), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(n965), .B(n964), .ZN(n967) );
  INV_X1 U1061 ( .A(G29), .ZN(n966) );
  NAND2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n968), .ZN(n1020) );
  XNOR2_X1 U1064 ( .A(G16), .B(KEYINPUT56), .ZN(n992) );
  XNOR2_X1 U1065 ( .A(G1341), .B(n969), .ZN(n970) );
  NOR2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1067 ( .A1(n973), .A2(n972), .ZN(n975) );
  XOR2_X1 U1068 ( .A(G171), .B(G1961), .Z(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n990) );
  XNOR2_X1 U1070 ( .A(n976), .B(G1956), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(G1971), .A2(G303), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(G1348), .B(n979), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G168), .ZN(n985) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1078 ( .A(KEYINPUT57), .B(n986), .Z(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n1018) );
  INV_X1 U1082 ( .A(G16), .ZN(n1016) );
  XNOR2_X1 U1083 ( .A(KEYINPUT61), .B(KEYINPUT127), .ZN(n1014) );
  XOR2_X1 U1084 ( .A(G1961), .B(G5), .Z(n1002) );
  XNOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT59), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n993), .B(G4), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(G1981), .B(G6), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(G19), .B(G1341), .ZN(n994) );
  NOR2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(G20), .B(G1956), .ZN(n998) );
  NOR2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(KEYINPUT60), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(G21), .B(G1966), .ZN(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(KEYINPUT126), .B(n1005), .ZN(n1012) );
  XOR2_X1 U1098 ( .A(G1976), .B(G23), .Z(n1007) );
  XOR2_X1 U1099 ( .A(G1971), .B(G22), .Z(n1006) );
  NAND2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(G24), .B(G1986), .ZN(n1008) );
  NOR2_X1 U1102 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1104 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1105 ( .A(n1014), .B(n1013), .ZN(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

