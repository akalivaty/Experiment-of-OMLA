

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X2 U555 ( .A1(n751), .A2(n750), .ZN(n764) );
  AND2_X1 U556 ( .A1(n831), .A2(n830), .ZN(n832) );
  AND2_X2 U557 ( .A1(n536), .A2(G2104), .ZN(n889) );
  OR2_X1 U558 ( .A1(n704), .A2(n939), .ZN(n705) );
  NAND2_X1 U559 ( .A1(n784), .A2(n690), .ZN(n692) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n784) );
  NOR2_X1 U561 ( .A1(G651), .A2(n648), .ZN(n651) );
  AND2_X1 U562 ( .A1(n762), .A2(n522), .ZN(n521) );
  AND2_X1 U563 ( .A1(n940), .A2(n761), .ZN(n522) );
  NOR2_X1 U564 ( .A1(n764), .A2(n754), .ZN(n523) );
  BUF_X1 U565 ( .A(n720), .Z(n709) );
  NOR2_X1 U566 ( .A1(n715), .A2(n714), .ZN(n716) );
  INV_X1 U567 ( .A(n952), .ZN(n752) );
  NAND2_X1 U568 ( .A1(n753), .A2(n752), .ZN(n754) );
  INV_X1 U569 ( .A(KEYINPUT32), .ZN(n743) );
  XNOR2_X1 U570 ( .A(n744), .B(n743), .ZN(n751) );
  NOR2_X1 U571 ( .A1(n648), .A2(n527), .ZN(n652) );
  XOR2_X1 U572 ( .A(KEYINPUT70), .B(n533), .Z(G299) );
  XOR2_X1 U573 ( .A(G543), .B(KEYINPUT0), .Z(n648) );
  NAND2_X1 U574 ( .A1(G53), .A2(n651), .ZN(n526) );
  INV_X1 U575 ( .A(G651), .ZN(n527) );
  NOR2_X1 U576 ( .A1(G543), .A2(n527), .ZN(n524) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n524), .Z(n600) );
  NAND2_X1 U578 ( .A1(G65), .A2(n600), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n532) );
  NAND2_X1 U580 ( .A1(G78), .A2(n652), .ZN(n529) );
  NOR2_X1 U581 ( .A1(G543), .A2(G651), .ZN(n653) );
  NAND2_X1 U582 ( .A1(G91), .A2(n653), .ZN(n528) );
  NAND2_X1 U583 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U584 ( .A(KEYINPUT69), .B(n530), .Z(n531) );
  NOR2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U586 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n535) );
  NOR2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n534) );
  XNOR2_X2 U588 ( .A(n535), .B(n534), .ZN(n888) );
  NAND2_X1 U589 ( .A1(n888), .A2(G137), .ZN(n539) );
  INV_X1 U590 ( .A(G2105), .ZN(n536) );
  NAND2_X1 U591 ( .A1(G101), .A2(n889), .ZN(n537) );
  XOR2_X1 U592 ( .A(n537), .B(KEYINPUT23), .Z(n538) );
  NAND2_X1 U593 ( .A1(n539), .A2(n538), .ZN(n543) );
  NOR2_X2 U594 ( .A1(G2104), .A2(n536), .ZN(n898) );
  NAND2_X1 U595 ( .A1(G125), .A2(n898), .ZN(n541) );
  AND2_X1 U596 ( .A1(G2105), .A2(G2104), .ZN(n894) );
  NAND2_X1 U597 ( .A1(G113), .A2(n894), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X2 U599 ( .A1(n543), .A2(n542), .ZN(G160) );
  NAND2_X1 U600 ( .A1(n888), .A2(G138), .ZN(n545) );
  NAND2_X1 U601 ( .A1(G102), .A2(n889), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G126), .A2(n898), .ZN(n547) );
  NAND2_X1 U604 ( .A1(G114), .A2(n894), .ZN(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U606 ( .A1(n549), .A2(n548), .ZN(G164) );
  XOR2_X1 U607 ( .A(G2446), .B(G2430), .Z(n551) );
  XNOR2_X1 U608 ( .A(G2451), .B(KEYINPUT102), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U610 ( .A(n552), .B(G2427), .Z(n554) );
  XNOR2_X1 U611 ( .A(G1341), .B(G1348), .ZN(n553) );
  XNOR2_X1 U612 ( .A(n554), .B(n553), .ZN(n558) );
  XOR2_X1 U613 ( .A(G2443), .B(G2435), .Z(n556) );
  XNOR2_X1 U614 ( .A(G2438), .B(G2454), .ZN(n555) );
  XNOR2_X1 U615 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U616 ( .A(n558), .B(n557), .Z(n559) );
  AND2_X1 U617 ( .A1(G14), .A2(n559), .ZN(G401) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  NAND2_X1 U622 ( .A1(G52), .A2(n651), .ZN(n561) );
  NAND2_X1 U623 ( .A1(G64), .A2(n600), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n653), .A2(G90), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n562), .B(KEYINPUT68), .ZN(n564) );
  NAND2_X1 U627 ( .A1(G77), .A2(n652), .ZN(n563) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U629 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  NOR2_X1 U630 ( .A1(n567), .A2(n566), .ZN(G171) );
  NAND2_X1 U631 ( .A1(G50), .A2(n651), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G62), .A2(n600), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U634 ( .A(KEYINPUT78), .B(n570), .Z(n574) );
  NAND2_X1 U635 ( .A1(n652), .A2(G75), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G88), .A2(n653), .ZN(n571) );
  AND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n574), .A2(n573), .ZN(G303) );
  NAND2_X1 U639 ( .A1(n653), .A2(G89), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT4), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G76), .A2(n652), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(KEYINPUT5), .ZN(n583) );
  NAND2_X1 U644 ( .A1(G51), .A2(n651), .ZN(n580) );
  NAND2_X1 U645 ( .A1(G63), .A2(n600), .ZN(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U647 ( .A(KEYINPUT6), .B(n581), .Z(n582) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U650 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U651 ( .A1(G7), .A2(G661), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n585), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U653 ( .A(G223), .ZN(n833) );
  NAND2_X1 U654 ( .A1(n833), .A2(G567), .ZN(n586) );
  XNOR2_X1 U655 ( .A(n586), .B(KEYINPUT71), .ZN(n587) );
  XNOR2_X1 U656 ( .A(KEYINPUT11), .B(n587), .ZN(G234) );
  NAND2_X1 U657 ( .A1(n653), .A2(G81), .ZN(n588) );
  XNOR2_X1 U658 ( .A(n588), .B(KEYINPUT12), .ZN(n590) );
  NAND2_X1 U659 ( .A1(G68), .A2(n652), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n592) );
  XOR2_X1 U661 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n591) );
  XNOR2_X1 U662 ( .A(n592), .B(n591), .ZN(n595) );
  NAND2_X1 U663 ( .A1(n600), .A2(G56), .ZN(n593) );
  XOR2_X1 U664 ( .A(KEYINPUT14), .B(n593), .Z(n594) );
  NOR2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n651), .A2(G43), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n944) );
  INV_X1 U668 ( .A(G860), .ZN(n626) );
  OR2_X1 U669 ( .A1(n944), .A2(n626), .ZN(G153) );
  INV_X1 U670 ( .A(G171), .ZN(G301) );
  NAND2_X1 U671 ( .A1(G868), .A2(G301), .ZN(n608) );
  NAND2_X1 U672 ( .A1(G79), .A2(n652), .ZN(n599) );
  NAND2_X1 U673 ( .A1(G54), .A2(n651), .ZN(n598) );
  NAND2_X1 U674 ( .A1(n599), .A2(n598), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G92), .A2(n653), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G66), .A2(n600), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U678 ( .A(KEYINPUT73), .B(n603), .Z(n604) );
  NOR2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n606) );
  XOR2_X2 U680 ( .A(KEYINPUT15), .B(n606), .Z(n939) );
  OR2_X1 U681 ( .A1(n939), .A2(G868), .ZN(n607) );
  NAND2_X1 U682 ( .A1(n608), .A2(n607), .ZN(G284) );
  INV_X1 U683 ( .A(G868), .ZN(n670) );
  NOR2_X1 U684 ( .A1(G286), .A2(n670), .ZN(n610) );
  NOR2_X1 U685 ( .A1(G299), .A2(G868), .ZN(n609) );
  NOR2_X1 U686 ( .A1(n610), .A2(n609), .ZN(G297) );
  NAND2_X1 U687 ( .A1(n626), .A2(G559), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n611), .A2(n939), .ZN(n612) );
  XNOR2_X1 U689 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U690 ( .A1(G868), .A2(n944), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G868), .A2(n939), .ZN(n613) );
  NOR2_X1 U692 ( .A1(G559), .A2(n613), .ZN(n614) );
  NOR2_X1 U693 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U694 ( .A1(n898), .A2(G123), .ZN(n616) );
  XNOR2_X1 U695 ( .A(n616), .B(KEYINPUT18), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G111), .A2(n894), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G135), .A2(n888), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G99), .A2(n889), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n1005) );
  XNOR2_X1 U702 ( .A(n1005), .B(G2096), .ZN(n624) );
  INV_X1 U703 ( .A(G2100), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(G156) );
  XOR2_X1 U705 ( .A(KEYINPUT74), .B(KEYINPUT76), .Z(n628) );
  NAND2_X1 U706 ( .A1(G559), .A2(n939), .ZN(n625) );
  XOR2_X1 U707 ( .A(n944), .B(n625), .Z(n668) );
  NAND2_X1 U708 ( .A1(n668), .A2(n626), .ZN(n627) );
  XNOR2_X1 U709 ( .A(n628), .B(n627), .ZN(n636) );
  NAND2_X1 U710 ( .A1(G80), .A2(n652), .ZN(n630) );
  NAND2_X1 U711 ( .A1(G67), .A2(n600), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U713 ( .A1(G93), .A2(n653), .ZN(n631) );
  XNOR2_X1 U714 ( .A(KEYINPUT75), .B(n631), .ZN(n632) );
  NOR2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n651), .A2(G55), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n671) );
  XOR2_X1 U718 ( .A(n636), .B(n671), .Z(G145) );
  NAND2_X1 U719 ( .A1(G86), .A2(n653), .ZN(n638) );
  NAND2_X1 U720 ( .A1(G61), .A2(n600), .ZN(n637) );
  NAND2_X1 U721 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n652), .A2(G73), .ZN(n639) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U724 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n651), .A2(G48), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n643), .A2(n642), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G49), .A2(n651), .ZN(n645) );
  NAND2_X1 U728 ( .A1(G74), .A2(G651), .ZN(n644) );
  NAND2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U730 ( .A(KEYINPUT77), .B(n646), .Z(n647) );
  NOR2_X1 U731 ( .A1(n600), .A2(n647), .ZN(n650) );
  NAND2_X1 U732 ( .A1(n648), .A2(G87), .ZN(n649) );
  NAND2_X1 U733 ( .A1(n650), .A2(n649), .ZN(G288) );
  NAND2_X1 U734 ( .A1(n651), .A2(G47), .ZN(n660) );
  NAND2_X1 U735 ( .A1(G72), .A2(n652), .ZN(n655) );
  NAND2_X1 U736 ( .A1(G85), .A2(n653), .ZN(n654) );
  NAND2_X1 U737 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U738 ( .A1(G60), .A2(n600), .ZN(n656) );
  XOR2_X1 U739 ( .A(KEYINPUT66), .B(n656), .Z(n657) );
  NOR2_X1 U740 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U741 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U742 ( .A(KEYINPUT67), .B(n661), .Z(G290) );
  XNOR2_X1 U743 ( .A(KEYINPUT79), .B(G305), .ZN(n662) );
  XNOR2_X1 U744 ( .A(n662), .B(n671), .ZN(n665) );
  XNOR2_X1 U745 ( .A(G299), .B(G303), .ZN(n663) );
  XNOR2_X1 U746 ( .A(n663), .B(G288), .ZN(n664) );
  XNOR2_X1 U747 ( .A(n665), .B(n664), .ZN(n667) );
  XNOR2_X1 U748 ( .A(G290), .B(KEYINPUT19), .ZN(n666) );
  XNOR2_X1 U749 ( .A(n667), .B(n666), .ZN(n839) );
  XOR2_X1 U750 ( .A(n839), .B(n668), .Z(n669) );
  NOR2_X1 U751 ( .A1(n670), .A2(n669), .ZN(n673) );
  NOR2_X1 U752 ( .A1(G868), .A2(n671), .ZN(n672) );
  NOR2_X1 U753 ( .A1(n673), .A2(n672), .ZN(G295) );
  XOR2_X1 U754 ( .A(KEYINPUT21), .B(KEYINPUT80), .Z(n677) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n674) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U757 ( .A1(n675), .A2(G2090), .ZN(n676) );
  XNOR2_X1 U758 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U759 ( .A(KEYINPUT81), .B(n678), .ZN(n679) );
  NAND2_X1 U760 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U762 ( .A1(G69), .A2(G120), .ZN(n680) );
  NOR2_X1 U763 ( .A1(G237), .A2(n680), .ZN(n681) );
  NAND2_X1 U764 ( .A1(G108), .A2(n681), .ZN(n837) );
  NAND2_X1 U765 ( .A1(n837), .A2(G567), .ZN(n687) );
  NOR2_X1 U766 ( .A1(G220), .A2(G219), .ZN(n682) );
  XNOR2_X1 U767 ( .A(KEYINPUT22), .B(n682), .ZN(n683) );
  NAND2_X1 U768 ( .A1(n683), .A2(G96), .ZN(n684) );
  NOR2_X1 U769 ( .A1(G218), .A2(n684), .ZN(n685) );
  XOR2_X1 U770 ( .A(KEYINPUT82), .B(n685), .Z(n838) );
  NAND2_X1 U771 ( .A1(G2106), .A2(n838), .ZN(n686) );
  NAND2_X1 U772 ( .A1(n687), .A2(n686), .ZN(n915) );
  NAND2_X1 U773 ( .A1(G483), .A2(G661), .ZN(n688) );
  NOR2_X1 U774 ( .A1(n915), .A2(n688), .ZN(n689) );
  XOR2_X1 U775 ( .A(KEYINPUT83), .B(n689), .Z(n836) );
  NAND2_X1 U776 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U777 ( .A1(G160), .A2(G40), .ZN(n783) );
  INV_X1 U778 ( .A(n783), .ZN(n690) );
  INV_X1 U779 ( .A(KEYINPUT64), .ZN(n691) );
  XNOR2_X1 U780 ( .A(n692), .B(n691), .ZN(n720) );
  INV_X1 U781 ( .A(n720), .ZN(n735) );
  NAND2_X1 U782 ( .A1(n735), .A2(G8), .ZN(n769) );
  NOR2_X1 U783 ( .A1(G1981), .A2(G305), .ZN(n693) );
  XOR2_X1 U784 ( .A(n693), .B(KEYINPUT24), .Z(n694) );
  NOR2_X1 U785 ( .A1(n769), .A2(n694), .ZN(n763) );
  NAND2_X1 U786 ( .A1(n720), .A2(G1996), .ZN(n695) );
  XNOR2_X1 U787 ( .A(n695), .B(KEYINPUT26), .ZN(n697) );
  NAND2_X1 U788 ( .A1(n735), .A2(G1341), .ZN(n696) );
  NAND2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U790 ( .A1(n698), .A2(n944), .ZN(n704) );
  NAND2_X1 U791 ( .A1(n704), .A2(n939), .ZN(n703) );
  AND2_X1 U792 ( .A1(n735), .A2(G1348), .ZN(n699) );
  XNOR2_X1 U793 ( .A(n699), .B(KEYINPUT93), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n709), .A2(G2067), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U796 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U798 ( .A(n707), .B(KEYINPUT94), .ZN(n713) );
  NAND2_X1 U799 ( .A1(G2072), .A2(n720), .ZN(n708) );
  XNOR2_X1 U800 ( .A(n708), .B(KEYINPUT27), .ZN(n711) );
  INV_X1 U801 ( .A(G1956), .ZN(n966) );
  NOR2_X1 U802 ( .A1(n709), .A2(n966), .ZN(n710) );
  NOR2_X1 U803 ( .A1(n711), .A2(n710), .ZN(n715) );
  INV_X1 U804 ( .A(G299), .ZN(n714) );
  NAND2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n712) );
  NAND2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n718) );
  XOR2_X1 U807 ( .A(n716), .B(KEYINPUT28), .Z(n717) );
  NAND2_X1 U808 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U809 ( .A(n719), .B(KEYINPUT29), .ZN(n724) );
  XOR2_X1 U810 ( .A(G2078), .B(KEYINPUT25), .Z(n921) );
  NOR2_X1 U811 ( .A1(n735), .A2(n921), .ZN(n722) );
  NOR2_X1 U812 ( .A1(G1961), .A2(n720), .ZN(n721) );
  NOR2_X1 U813 ( .A1(n722), .A2(n721), .ZN(n728) );
  NOR2_X1 U814 ( .A1(G301), .A2(n728), .ZN(n723) );
  NOR2_X1 U815 ( .A1(n724), .A2(n723), .ZN(n733) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n769), .ZN(n749) );
  NOR2_X1 U817 ( .A1(n735), .A2(G2084), .ZN(n746) );
  NOR2_X1 U818 ( .A1(n749), .A2(n746), .ZN(n725) );
  NAND2_X1 U819 ( .A1(G8), .A2(n725), .ZN(n726) );
  XNOR2_X1 U820 ( .A(KEYINPUT30), .B(n726), .ZN(n727) );
  NOR2_X1 U821 ( .A1(G168), .A2(n727), .ZN(n730) );
  AND2_X1 U822 ( .A1(G301), .A2(n728), .ZN(n729) );
  NOR2_X1 U823 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U824 ( .A(n731), .B(KEYINPUT31), .ZN(n732) );
  XNOR2_X1 U825 ( .A(n734), .B(KEYINPUT95), .ZN(n745) );
  NAND2_X1 U826 ( .A1(n745), .A2(G286), .ZN(n742) );
  INV_X1 U827 ( .A(G8), .ZN(n740) );
  NOR2_X1 U828 ( .A1(n735), .A2(G2090), .ZN(n737) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n769), .ZN(n736) );
  NOR2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U831 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U832 ( .A1(n740), .A2(n739), .ZN(n741) );
  AND2_X1 U833 ( .A1(n742), .A2(n741), .ZN(n744) );
  NAND2_X1 U834 ( .A1(G8), .A2(n746), .ZN(n747) );
  NAND2_X1 U835 ( .A1(n745), .A2(n747), .ZN(n748) );
  NOR2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U837 ( .A1(G1971), .A2(G303), .ZN(n951) );
  XOR2_X1 U838 ( .A(n951), .B(KEYINPUT96), .Z(n753) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n952) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n950) );
  INV_X1 U841 ( .A(n769), .ZN(n755) );
  NAND2_X1 U842 ( .A1(n950), .A2(n755), .ZN(n756) );
  NOR2_X1 U843 ( .A1(n523), .A2(n756), .ZN(n757) );
  NOR2_X1 U844 ( .A1(n757), .A2(KEYINPUT33), .ZN(n758) );
  XNOR2_X1 U845 ( .A(n758), .B(KEYINPUT97), .ZN(n762) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n940) );
  NAND2_X1 U847 ( .A1(n952), .A2(KEYINPUT33), .ZN(n759) );
  NOR2_X1 U848 ( .A1(n769), .A2(n759), .ZN(n760) );
  XOR2_X1 U849 ( .A(KEYINPUT98), .B(n760), .Z(n761) );
  NOR2_X1 U850 ( .A1(n763), .A2(n521), .ZN(n817) );
  INV_X1 U851 ( .A(n764), .ZN(n767) );
  NOR2_X1 U852 ( .A1(G2090), .A2(G303), .ZN(n765) );
  NAND2_X1 U853 ( .A1(G8), .A2(n765), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U855 ( .A1(n769), .A2(n768), .ZN(n815) );
  NAND2_X1 U856 ( .A1(G140), .A2(n888), .ZN(n771) );
  NAND2_X1 U857 ( .A1(G104), .A2(n889), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U859 ( .A(KEYINPUT34), .B(n772), .ZN(n779) );
  NAND2_X1 U860 ( .A1(n898), .A2(G128), .ZN(n773) );
  XNOR2_X1 U861 ( .A(n773), .B(KEYINPUT84), .ZN(n775) );
  NAND2_X1 U862 ( .A1(G116), .A2(n894), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U864 ( .A(KEYINPUT85), .B(n776), .ZN(n777) );
  XNOR2_X1 U865 ( .A(KEYINPUT35), .B(n777), .ZN(n778) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U867 ( .A(n780), .B(KEYINPUT36), .Z(n781) );
  XOR2_X1 U868 ( .A(KEYINPUT86), .B(n781), .Z(n905) );
  XNOR2_X1 U869 ( .A(KEYINPUT37), .B(G2067), .ZN(n785) );
  AND2_X1 U870 ( .A1(n905), .A2(n785), .ZN(n782) );
  XNOR2_X1 U871 ( .A(n782), .B(KEYINPUT101), .ZN(n1014) );
  NOR2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n820) );
  NOR2_X1 U873 ( .A1(n905), .A2(n785), .ZN(n1012) );
  NAND2_X1 U874 ( .A1(n820), .A2(n1012), .ZN(n822) );
  XOR2_X1 U875 ( .A(KEYINPUT39), .B(KEYINPUT100), .Z(n811) );
  NAND2_X1 U876 ( .A1(G105), .A2(n889), .ZN(n786) );
  XNOR2_X1 U877 ( .A(n786), .B(KEYINPUT38), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G117), .A2(n894), .ZN(n787) );
  XNOR2_X1 U879 ( .A(n787), .B(KEYINPUT90), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n888), .A2(G141), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U882 ( .A1(G129), .A2(n898), .ZN(n790) );
  XNOR2_X1 U883 ( .A(KEYINPUT89), .B(n790), .ZN(n791) );
  NOR2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n871) );
  NOR2_X1 U886 ( .A1(G1996), .A2(n871), .ZN(n999) );
  NAND2_X1 U887 ( .A1(G1996), .A2(n871), .ZN(n795) );
  XOR2_X1 U888 ( .A(KEYINPUT91), .B(n795), .Z(n805) );
  NAND2_X1 U889 ( .A1(n894), .A2(G107), .ZN(n796) );
  XOR2_X1 U890 ( .A(KEYINPUT87), .B(n796), .Z(n798) );
  NAND2_X1 U891 ( .A1(n898), .A2(G119), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U893 ( .A(KEYINPUT88), .B(n799), .Z(n803) );
  NAND2_X1 U894 ( .A1(G131), .A2(n888), .ZN(n801) );
  NAND2_X1 U895 ( .A1(G95), .A2(n889), .ZN(n800) );
  AND2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n902) );
  NAND2_X1 U898 ( .A1(G1991), .A2(n902), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n1001) );
  AND2_X1 U900 ( .A1(n1001), .A2(n820), .ZN(n823) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n902), .ZN(n806) );
  XOR2_X1 U902 ( .A(KEYINPUT99), .B(n806), .Z(n1004) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n1004), .A2(n807), .ZN(n808) );
  NOR2_X1 U905 ( .A1(n823), .A2(n808), .ZN(n809) );
  NOR2_X1 U906 ( .A1(n999), .A2(n809), .ZN(n810) );
  XOR2_X1 U907 ( .A(n811), .B(n810), .Z(n812) );
  NAND2_X1 U908 ( .A1(n822), .A2(n812), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n1014), .A2(n813), .ZN(n814) );
  NAND2_X1 U910 ( .A1(n814), .A2(n820), .ZN(n818) );
  AND2_X1 U911 ( .A1(n815), .A2(n818), .ZN(n816) );
  NAND2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n831) );
  INV_X1 U913 ( .A(n818), .ZN(n829) );
  XOR2_X1 U914 ( .A(G1986), .B(G290), .Z(n957) );
  NAND2_X1 U915 ( .A1(KEYINPUT92), .A2(n1001), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n957), .A2(n819), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n827) );
  XOR2_X1 U918 ( .A(n822), .B(KEYINPUT92), .Z(n825) );
  INV_X1 U919 ( .A(n823), .ZN(n824) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n826) );
  AND2_X1 U921 ( .A1(n827), .A2(n826), .ZN(n828) );
  OR2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U923 ( .A(n832), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U926 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G69), .ZN(G235) );
  NOR2_X1 U933 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U934 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U935 ( .A(n839), .B(KEYINPUT110), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n944), .B(G286), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n841), .B(n840), .ZN(n843) );
  XOR2_X1 U938 ( .A(n939), .B(G171), .Z(n842) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(n844) );
  NOR2_X1 U940 ( .A1(G37), .A2(n844), .ZN(n845) );
  XOR2_X1 U941 ( .A(KEYINPUT111), .B(n845), .Z(G397) );
  XOR2_X1 U942 ( .A(KEYINPUT103), .B(G2090), .Z(n847) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2084), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U945 ( .A(n848), .B(G2100), .Z(n850) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2072), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U948 ( .A(G2096), .B(KEYINPUT43), .Z(n852) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(G2678), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U951 ( .A(n854), .B(n853), .Z(G227) );
  XOR2_X1 U952 ( .A(G1981), .B(G1961), .Z(n856) );
  XNOR2_X1 U953 ( .A(G1986), .B(G1966), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U955 ( .A(n857), .B(G2474), .Z(n859) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U958 ( .A(KEYINPUT41), .B(G1976), .Z(n861) );
  XNOR2_X1 U959 ( .A(G1956), .B(G1971), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(G229) );
  NAND2_X1 U962 ( .A1(n898), .A2(G124), .ZN(n864) );
  XNOR2_X1 U963 ( .A(n864), .B(KEYINPUT44), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G112), .A2(n894), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n866), .A2(n865), .ZN(n870) );
  NAND2_X1 U966 ( .A1(G136), .A2(n888), .ZN(n868) );
  NAND2_X1 U967 ( .A1(G100), .A2(n889), .ZN(n867) );
  NAND2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U969 ( .A1(n870), .A2(n869), .ZN(G162) );
  XNOR2_X1 U970 ( .A(G162), .B(n871), .ZN(n881) );
  NAND2_X1 U971 ( .A1(G139), .A2(n888), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G103), .A2(n889), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n874), .B(KEYINPUT107), .ZN(n880) );
  XNOR2_X1 U975 ( .A(KEYINPUT108), .B(KEYINPUT47), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G127), .A2(n898), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G115), .A2(n894), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n878), .B(n877), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n1017) );
  XNOR2_X1 U981 ( .A(n881), .B(n1017), .ZN(n885) );
  XOR2_X1 U982 ( .A(KEYINPUT48), .B(KEYINPUT109), .Z(n883) );
  XNOR2_X1 U983 ( .A(n1005), .B(KEYINPUT46), .ZN(n882) );
  XNOR2_X1 U984 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U985 ( .A(n885), .B(n884), .Z(n887) );
  XNOR2_X1 U986 ( .A(G164), .B(G160), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n907) );
  NAND2_X1 U988 ( .A1(G142), .A2(n888), .ZN(n891) );
  NAND2_X1 U989 ( .A1(G106), .A2(n889), .ZN(n890) );
  NAND2_X1 U990 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U991 ( .A(n892), .B(KEYINPUT106), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n893), .B(KEYINPUT45), .ZN(n897) );
  NAND2_X1 U993 ( .A1(G118), .A2(n894), .ZN(n895) );
  XOR2_X1 U994 ( .A(KEYINPUT105), .B(n895), .Z(n896) );
  NAND2_X1 U995 ( .A1(n897), .A2(n896), .ZN(n901) );
  NAND2_X1 U996 ( .A1(n898), .A2(G130), .ZN(n899) );
  XOR2_X1 U997 ( .A(n899), .B(KEYINPUT104), .Z(n900) );
  NOR2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n908), .ZN(G395) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n915), .ZN(n912) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1005 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G397), .A2(n910), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(n913), .A2(G395), .ZN(n914) );
  XNOR2_X1 U1009 ( .A(n914), .B(KEYINPUT112), .ZN(G308) );
  INV_X1 U1010 ( .A(G308), .ZN(G225) );
  INV_X1 U1011 ( .A(G303), .ZN(G166) );
  INV_X1 U1012 ( .A(n915), .ZN(G319) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1014 ( .A(G2090), .B(G35), .Z(n932) );
  XNOR2_X1 U1015 ( .A(G1991), .B(G25), .ZN(n927) );
  XNOR2_X1 U1016 ( .A(G2072), .B(KEYINPUT117), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n916), .B(G33), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(G2067), .B(G26), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(G1996), .B(G32), .ZN(n917) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(G27), .B(n921), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(KEYINPUT118), .B(n922), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(KEYINPUT119), .B(n925), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1027 ( .A1(n928), .A2(G28), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(n929), .B(KEYINPUT120), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(n930), .B(KEYINPUT53), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(G34), .B(G2084), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(KEYINPUT54), .B(n933), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(KEYINPUT55), .B(n936), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(KEYINPUT121), .B(n937), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(G29), .A2(n938), .ZN(n995) );
  XNOR2_X1 U1037 ( .A(G16), .B(KEYINPUT56), .ZN(n965) );
  XNOR2_X1 U1038 ( .A(n939), .B(G1348), .ZN(n963) );
  XNOR2_X1 U1039 ( .A(G1966), .B(G168), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(n942), .B(KEYINPUT57), .ZN(n948) );
  XOR2_X1 U1042 ( .A(G1341), .B(KEYINPUT123), .Z(n943) );
  XNOR2_X1 U1043 ( .A(n944), .B(n943), .ZN(n946) );
  XOR2_X1 U1044 ( .A(G1961), .B(G171), .Z(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n961) );
  NAND2_X1 U1047 ( .A1(G1971), .A2(G303), .ZN(n949) );
  NAND2_X1 U1048 ( .A1(n950), .A2(n949), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G299), .B(n966), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(KEYINPUT122), .B(n959), .ZN(n960) );
  NOR2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n993) );
  INV_X1 U1058 ( .A(G16), .ZN(n991) );
  XNOR2_X1 U1059 ( .A(G1966), .B(G21), .ZN(n977) );
  XOR2_X1 U1060 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n975) );
  XNOR2_X1 U1061 ( .A(G20), .B(n966), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(G1341), .B(G19), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(G6), .B(G1981), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1066 ( .A(KEYINPUT59), .B(G1348), .Z(n971) );
  XNOR2_X1 U1067 ( .A(G4), .B(n971), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n975), .B(n974), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1071 ( .A(KEYINPUT125), .B(n978), .Z(n986) );
  XNOR2_X1 U1072 ( .A(G1971), .B(G22), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(G23), .B(G1976), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1075 ( .A(KEYINPUT126), .B(n981), .Z(n983) );
  XNOR2_X1 U1076 ( .A(G1986), .B(G24), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(KEYINPUT58), .B(n984), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(G5), .B(G1961), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(KEYINPUT61), .B(n989), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(G11), .A2(n996), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(n997), .B(KEYINPUT127), .ZN(n1029) );
  XOR2_X1 U1088 ( .A(G2090), .B(G162), .Z(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1090 ( .A(KEYINPUT51), .B(n1000), .Z(n1010) );
  XNOR2_X1 U1091 ( .A(G160), .B(G2084), .ZN(n1003) );
  INV_X1 U1092 ( .A(n1001), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1008) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(KEYINPUT113), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1099 ( .A(n1013), .B(KEYINPUT114), .ZN(n1015) );
  NAND2_X1 U1100 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1101 ( .A(KEYINPUT115), .B(n1016), .Z(n1023) );
  XOR2_X1 U1102 ( .A(G164), .B(G2078), .Z(n1020) );
  XNOR2_X1 U1103 ( .A(KEYINPUT116), .B(n1017), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(G2072), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1106 ( .A(KEYINPUT50), .B(n1021), .Z(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(KEYINPUT52), .B(n1024), .ZN(n1026) );
  INV_X1 U1109 ( .A(KEYINPUT55), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1111 ( .A1(n1027), .A2(G29), .ZN(n1028) );
  NAND2_X1 U1112 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

