

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U553 ( .A1(n689), .A2(n777), .ZN(n732) );
  NOR2_X1 U554 ( .A1(n702), .A2(n907), .ZN(n697) );
  NOR2_X1 U555 ( .A1(n815), .A2(n754), .ZN(n755) );
  INV_X1 U556 ( .A(KEYINPUT66), .ZN(n533) );
  NAND2_X1 U557 ( .A1(n519), .A2(n758), .ZN(n807) );
  INV_X1 U558 ( .A(KEYINPUT33), .ZN(n758) );
  NAND2_X1 U559 ( .A1(n607), .A2(G113), .ZN(n541) );
  XNOR2_X1 U560 ( .A(n535), .B(n534), .ZN(n538) );
  XNOR2_X1 U561 ( .A(n533), .B(KEYINPUT23), .ZN(n534) );
  AND2_X2 U562 ( .A1(G2105), .A2(G2104), .ZN(n607) );
  XOR2_X1 U563 ( .A(n757), .B(KEYINPUT64), .Z(n519) );
  OR2_X1 U564 ( .A1(n804), .A2(n815), .ZN(n520) );
  INV_X1 U565 ( .A(KEYINPUT96), .ZN(n688) );
  INV_X1 U566 ( .A(n901), .ZN(n754) );
  AND2_X1 U567 ( .A1(n756), .A2(n755), .ZN(n757) );
  INV_X1 U568 ( .A(KEYINPUT17), .ZN(n542) );
  AND2_X1 U569 ( .A1(n805), .A2(n520), .ZN(n806) );
  NOR2_X1 U570 ( .A1(G651), .A2(n629), .ZN(n640) );
  NOR2_X1 U571 ( .A1(G651), .A2(G543), .ZN(n647) );
  NAND2_X1 U572 ( .A1(n647), .A2(G89), .ZN(n521) );
  XNOR2_X1 U573 ( .A(n521), .B(KEYINPUT4), .ZN(n523) );
  XOR2_X1 U574 ( .A(KEYINPUT0), .B(G543), .Z(n629) );
  INV_X1 U575 ( .A(G651), .ZN(n525) );
  NOR2_X1 U576 ( .A1(n629), .A2(n525), .ZN(n643) );
  NAND2_X1 U577 ( .A1(G76), .A2(n643), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U579 ( .A(n524), .B(KEYINPUT5), .ZN(n531) );
  NOR2_X1 U580 ( .A1(G543), .A2(n525), .ZN(n526) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n526), .Z(n639) );
  NAND2_X1 U582 ( .A1(G63), .A2(n639), .ZN(n528) );
  NAND2_X1 U583 ( .A1(G51), .A2(n640), .ZN(n527) );
  NAND2_X1 U584 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U585 ( .A(KEYINPUT6), .B(n529), .Z(n530) );
  NAND2_X1 U586 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U587 ( .A(n532), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U588 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XNOR2_X1 U589 ( .A(G2104), .B(KEYINPUT65), .ZN(n536) );
  NOR2_X1 U590 ( .A1(n536), .A2(G2105), .ZN(n603) );
  NAND2_X1 U591 ( .A1(G101), .A2(n603), .ZN(n535) );
  AND2_X1 U592 ( .A1(n536), .A2(G2105), .ZN(n985) );
  NAND2_X1 U593 ( .A1(G125), .A2(n985), .ZN(n537) );
  NAND2_X1 U594 ( .A1(n538), .A2(n537), .ZN(n540) );
  INV_X1 U595 ( .A(KEYINPUT67), .ZN(n539) );
  XNOR2_X1 U596 ( .A(n540), .B(n539), .ZN(n548) );
  XNOR2_X1 U597 ( .A(n541), .B(KEYINPUT68), .ZN(n545) );
  NOR2_X1 U598 ( .A1(G2105), .A2(G2104), .ZN(n543) );
  XNOR2_X1 U599 ( .A(n543), .B(n542), .ZN(n608) );
  NAND2_X1 U600 ( .A1(n608), .A2(G137), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U602 ( .A(KEYINPUT69), .B(n546), .Z(n547) );
  NOR2_X2 U603 ( .A1(n548), .A2(n547), .ZN(G160) );
  NAND2_X1 U604 ( .A1(G64), .A2(n639), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G52), .A2(n640), .ZN(n549) );
  NAND2_X1 U606 ( .A1(n550), .A2(n549), .ZN(n555) );
  NAND2_X1 U607 ( .A1(G90), .A2(n647), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G77), .A2(n643), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U611 ( .A1(n555), .A2(n554), .ZN(G171) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U613 ( .A(G69), .ZN(G235) );
  INV_X1 U614 ( .A(G120), .ZN(G236) );
  INV_X1 U615 ( .A(G132), .ZN(G219) );
  INV_X1 U616 ( .A(G82), .ZN(G220) );
  NAND2_X1 U617 ( .A1(G88), .A2(n647), .ZN(n557) );
  NAND2_X1 U618 ( .A1(G75), .A2(n643), .ZN(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G62), .A2(n639), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G50), .A2(n640), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U623 ( .A1(n561), .A2(n560), .ZN(G166) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U625 ( .A(n562), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U626 ( .A(G223), .B(KEYINPUT72), .Z(n826) );
  NAND2_X1 U627 ( .A1(n826), .A2(G567), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  XNOR2_X1 U629 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n647), .A2(G81), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G68), .A2(n643), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n639), .A2(G56), .ZN(n569) );
  XOR2_X1 U636 ( .A(KEYINPUT14), .B(n569), .Z(n570) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n640), .A2(G43), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n1004) );
  INV_X1 U640 ( .A(G860), .ZN(n623) );
  OR2_X1 U641 ( .A1(n1004), .A2(n623), .ZN(G153) );
  XOR2_X1 U642 ( .A(G171), .B(KEYINPUT74), .Z(G301) );
  NAND2_X1 U643 ( .A1(n647), .A2(G92), .ZN(n580) );
  NAND2_X1 U644 ( .A1(G66), .A2(n639), .ZN(n575) );
  NAND2_X1 U645 ( .A1(G54), .A2(n640), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n643), .A2(G79), .ZN(n576) );
  XOR2_X1 U648 ( .A(KEYINPUT76), .B(n576), .Z(n577) );
  NOR2_X1 U649 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U651 ( .A(KEYINPUT15), .B(n581), .Z(n907) );
  INV_X1 U652 ( .A(n907), .ZN(n1005) );
  NOR2_X1 U653 ( .A1(n1005), .A2(G868), .ZN(n582) );
  XNOR2_X1 U654 ( .A(KEYINPUT77), .B(n582), .ZN(n585) );
  NAND2_X1 U655 ( .A1(G868), .A2(G301), .ZN(n583) );
  XOR2_X1 U656 ( .A(KEYINPUT75), .B(n583), .Z(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U658 ( .A1(G65), .A2(n639), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G53), .A2(n640), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G91), .A2(n647), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G78), .A2(n643), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n897) );
  INV_X1 U665 ( .A(n897), .ZN(G299) );
  NOR2_X1 U666 ( .A1(G868), .A2(G299), .ZN(n592) );
  XOR2_X1 U667 ( .A(KEYINPUT79), .B(n592), .Z(n595) );
  INV_X1 U668 ( .A(G868), .ZN(n659) );
  NOR2_X1 U669 ( .A1(G286), .A2(n659), .ZN(n593) );
  XNOR2_X1 U670 ( .A(KEYINPUT78), .B(n593), .ZN(n594) );
  NOR2_X1 U671 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U672 ( .A1(n623), .A2(G559), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n596), .A2(n1005), .ZN(n597) );
  XNOR2_X1 U674 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U675 ( .A1(n1005), .A2(G868), .ZN(n598) );
  NOR2_X1 U676 ( .A1(G559), .A2(n598), .ZN(n599) );
  XNOR2_X1 U677 ( .A(n599), .B(KEYINPUT80), .ZN(n601) );
  NOR2_X1 U678 ( .A1(n1004), .A2(G868), .ZN(n600) );
  NOR2_X1 U679 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G123), .A2(n985), .ZN(n602) );
  XNOR2_X1 U681 ( .A(n602), .B(KEYINPUT18), .ZN(n606) );
  BUF_X1 U682 ( .A(n603), .Z(n989) );
  NAND2_X1 U683 ( .A1(G99), .A2(n989), .ZN(n604) );
  XOR2_X1 U684 ( .A(KEYINPUT81), .B(n604), .Z(n605) );
  NAND2_X1 U685 ( .A1(n606), .A2(n605), .ZN(n612) );
  NAND2_X1 U686 ( .A1(G111), .A2(n607), .ZN(n610) );
  BUF_X1 U687 ( .A(n608), .Z(n991) );
  NAND2_X1 U688 ( .A1(G135), .A2(n991), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n980) );
  XNOR2_X1 U691 ( .A(n980), .B(G2096), .ZN(n614) );
  INV_X1 U692 ( .A(G2100), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U694 ( .A1(G67), .A2(n639), .ZN(n616) );
  NAND2_X1 U695 ( .A1(G55), .A2(n640), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U697 ( .A1(G80), .A2(n643), .ZN(n617) );
  XNOR2_X1 U698 ( .A(KEYINPUT83), .B(n617), .ZN(n618) );
  NOR2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U700 ( .A1(n647), .A2(G93), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n660) );
  XNOR2_X1 U702 ( .A(n660), .B(KEYINPUT82), .ZN(n625) );
  NAND2_X1 U703 ( .A1(G559), .A2(n1005), .ZN(n622) );
  XOR2_X1 U704 ( .A(n1004), .B(n622), .Z(n656) );
  NAND2_X1 U705 ( .A1(n656), .A2(n623), .ZN(n624) );
  XNOR2_X1 U706 ( .A(n625), .B(n624), .ZN(G145) );
  NAND2_X1 U707 ( .A1(G49), .A2(n640), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G74), .A2(G651), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U710 ( .A1(n639), .A2(n628), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n629), .A2(G87), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U713 ( .A1(G60), .A2(n639), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G47), .A2(n640), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U716 ( .A1(G85), .A2(n647), .ZN(n635) );
  NAND2_X1 U717 ( .A1(G72), .A2(n643), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U720 ( .A(KEYINPUT70), .B(n638), .Z(G290) );
  NAND2_X1 U721 ( .A1(G61), .A2(n639), .ZN(n642) );
  NAND2_X1 U722 ( .A1(G48), .A2(n640), .ZN(n641) );
  NAND2_X1 U723 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U724 ( .A1(n643), .A2(G73), .ZN(n644) );
  XOR2_X1 U725 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n649) );
  NAND2_X1 U727 ( .A1(n647), .A2(G86), .ZN(n648) );
  NAND2_X1 U728 ( .A1(n649), .A2(n648), .ZN(G305) );
  XNOR2_X1 U729 ( .A(n897), .B(G288), .ZN(n655) );
  XOR2_X1 U730 ( .A(KEYINPUT84), .B(KEYINPUT19), .Z(n651) );
  XNOR2_X1 U731 ( .A(G290), .B(G166), .ZN(n650) );
  XNOR2_X1 U732 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U733 ( .A(n652), .B(G305), .Z(n653) );
  XNOR2_X1 U734 ( .A(n660), .B(n653), .ZN(n654) );
  XNOR2_X1 U735 ( .A(n655), .B(n654), .ZN(n1003) );
  XNOR2_X1 U736 ( .A(n1003), .B(n656), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n657), .A2(G868), .ZN(n658) );
  XNOR2_X1 U738 ( .A(n658), .B(KEYINPUT85), .ZN(n662) );
  AND2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U740 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U741 ( .A(KEYINPUT86), .B(n663), .Z(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n664) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n665), .ZN(n667) );
  XOR2_X1 U745 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n666) );
  XNOR2_X1 U746 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U747 ( .A1(G2072), .A2(n668), .ZN(G158) );
  XNOR2_X1 U748 ( .A(KEYINPUT88), .B(G44), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n669), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U750 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U753 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U754 ( .A1(G96), .A2(n672), .ZN(n951) );
  NAND2_X1 U755 ( .A1(n951), .A2(G2106), .ZN(n677) );
  NOR2_X1 U756 ( .A1(G237), .A2(G236), .ZN(n673) );
  NAND2_X1 U757 ( .A1(G108), .A2(n673), .ZN(n674) );
  NOR2_X1 U758 ( .A1(n674), .A2(G235), .ZN(n675) );
  XNOR2_X1 U759 ( .A(n675), .B(KEYINPUT89), .ZN(n952) );
  NAND2_X1 U760 ( .A1(n952), .A2(G567), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n972) );
  NAND2_X1 U762 ( .A1(G661), .A2(G483), .ZN(n678) );
  XNOR2_X1 U763 ( .A(KEYINPUT90), .B(n678), .ZN(n679) );
  NOR2_X1 U764 ( .A1(n972), .A2(n679), .ZN(n829) );
  NAND2_X1 U765 ( .A1(n829), .A2(G36), .ZN(G176) );
  NAND2_X1 U766 ( .A1(G102), .A2(n989), .ZN(n681) );
  NAND2_X1 U767 ( .A1(G138), .A2(n991), .ZN(n680) );
  NAND2_X1 U768 ( .A1(n681), .A2(n680), .ZN(n686) );
  NAND2_X1 U769 ( .A1(G126), .A2(n985), .ZN(n683) );
  NAND2_X1 U770 ( .A1(G114), .A2(n607), .ZN(n682) );
  NAND2_X1 U771 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U772 ( .A(KEYINPUT91), .B(n684), .Z(n685) );
  NOR2_X1 U773 ( .A1(n686), .A2(n685), .ZN(G164) );
  INV_X1 U774 ( .A(G166), .ZN(G303) );
  INV_X1 U775 ( .A(n1004), .ZN(n692) );
  NAND2_X1 U776 ( .A1(G40), .A2(G160), .ZN(n687) );
  XNOR2_X1 U777 ( .A(n687), .B(KEYINPUT92), .ZN(n778) );
  XNOR2_X1 U778 ( .A(n778), .B(n688), .ZN(n689) );
  NOR2_X1 U779 ( .A1(G164), .A2(G1384), .ZN(n777) );
  NAND2_X1 U780 ( .A1(n732), .A2(G1341), .ZN(n690) );
  XNOR2_X1 U781 ( .A(n690), .B(KEYINPUT102), .ZN(n691) );
  AND2_X1 U782 ( .A1(n692), .A2(n691), .ZN(n696) );
  INV_X1 U783 ( .A(n732), .ZN(n693) );
  NAND2_X1 U784 ( .A1(G1996), .A2(n693), .ZN(n694) );
  XNOR2_X1 U785 ( .A(KEYINPUT26), .B(n694), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n702) );
  XNOR2_X1 U787 ( .A(n697), .B(KEYINPUT103), .ZN(n701) );
  XNOR2_X1 U788 ( .A(KEYINPUT99), .B(n732), .ZN(n705) );
  BUF_X1 U789 ( .A(n705), .Z(n718) );
  NAND2_X1 U790 ( .A1(G2067), .A2(n718), .ZN(n699) );
  NAND2_X1 U791 ( .A1(G1348), .A2(n732), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n704) );
  NAND2_X1 U794 ( .A1(n702), .A2(n907), .ZN(n703) );
  NAND2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n710) );
  NAND2_X1 U796 ( .A1(n705), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U797 ( .A(n706), .B(KEYINPUT27), .ZN(n708) );
  XOR2_X1 U798 ( .A(G1956), .B(KEYINPUT100), .Z(n923) );
  NOR2_X1 U799 ( .A1(n718), .A2(n923), .ZN(n707) );
  NOR2_X1 U800 ( .A1(n708), .A2(n707), .ZN(n711) );
  NAND2_X1 U801 ( .A1(n897), .A2(n711), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n715) );
  NOR2_X1 U803 ( .A1(n897), .A2(n711), .ZN(n713) );
  XNOR2_X1 U804 ( .A(KEYINPUT101), .B(KEYINPUT28), .ZN(n712) );
  XNOR2_X1 U805 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n715), .A2(n714), .ZN(n717) );
  XOR2_X1 U807 ( .A(KEYINPUT29), .B(KEYINPUT104), .Z(n716) );
  XNOR2_X1 U808 ( .A(n717), .B(n716), .ZN(n722) );
  INV_X1 U809 ( .A(G1961), .ZN(n917) );
  NAND2_X1 U810 ( .A1(n917), .A2(n732), .ZN(n720) );
  XNOR2_X1 U811 ( .A(G2078), .B(KEYINPUT25), .ZN(n876) );
  NAND2_X1 U812 ( .A1(n718), .A2(n876), .ZN(n719) );
  NAND2_X1 U813 ( .A1(n720), .A2(n719), .ZN(n726) );
  NAND2_X1 U814 ( .A1(n726), .A2(G171), .ZN(n721) );
  NAND2_X1 U815 ( .A1(n722), .A2(n721), .ZN(n731) );
  NAND2_X1 U816 ( .A1(G8), .A2(n732), .ZN(n815) );
  NOR2_X1 U817 ( .A1(G1966), .A2(n815), .ZN(n745) );
  NOR2_X1 U818 ( .A1(G2084), .A2(n732), .ZN(n741) );
  NOR2_X1 U819 ( .A1(n745), .A2(n741), .ZN(n723) );
  NAND2_X1 U820 ( .A1(G8), .A2(n723), .ZN(n724) );
  XNOR2_X1 U821 ( .A(KEYINPUT30), .B(n724), .ZN(n725) );
  NOR2_X1 U822 ( .A1(G168), .A2(n725), .ZN(n728) );
  NOR2_X1 U823 ( .A1(G171), .A2(n726), .ZN(n727) );
  NOR2_X1 U824 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U825 ( .A(KEYINPUT31), .B(n729), .Z(n730) );
  NAND2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n743) );
  NAND2_X1 U827 ( .A1(n743), .A2(G286), .ZN(n737) );
  NOR2_X1 U828 ( .A1(G1971), .A2(n815), .ZN(n734) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U830 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U831 ( .A1(n735), .A2(G303), .ZN(n736) );
  NAND2_X1 U832 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U833 ( .A(n738), .B(KEYINPUT106), .ZN(n739) );
  NAND2_X1 U834 ( .A1(n739), .A2(G8), .ZN(n740) );
  XNOR2_X1 U835 ( .A(n740), .B(KEYINPUT32), .ZN(n750) );
  NAND2_X1 U836 ( .A1(G8), .A2(n741), .ZN(n742) );
  XNOR2_X1 U837 ( .A(KEYINPUT98), .B(n742), .ZN(n748) );
  INV_X1 U838 ( .A(n743), .ZN(n744) );
  NOR2_X1 U839 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U840 ( .A(KEYINPUT105), .B(n746), .Z(n747) );
  NAND2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U842 ( .A1(n750), .A2(n749), .ZN(n811) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n752) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n751) );
  XOR2_X1 U845 ( .A(KEYINPUT107), .B(n751), .Z(n900) );
  NOR2_X1 U846 ( .A1(n752), .A2(n900), .ZN(n753) );
  NAND2_X1 U847 ( .A1(n811), .A2(n753), .ZN(n756) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n901) );
  XOR2_X1 U849 ( .A(G1981), .B(G305), .Z(n894) );
  NAND2_X1 U850 ( .A1(G117), .A2(n607), .ZN(n760) );
  NAND2_X1 U851 ( .A1(G141), .A2(n991), .ZN(n759) );
  NAND2_X1 U852 ( .A1(n760), .A2(n759), .ZN(n764) );
  NAND2_X1 U853 ( .A1(G105), .A2(n989), .ZN(n761) );
  XNOR2_X1 U854 ( .A(n761), .B(KEYINPUT95), .ZN(n762) );
  XNOR2_X1 U855 ( .A(n762), .B(KEYINPUT38), .ZN(n763) );
  NOR2_X1 U856 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U857 ( .A1(n985), .A2(G129), .ZN(n765) );
  NAND2_X1 U858 ( .A1(n766), .A2(n765), .ZN(n982) );
  NOR2_X1 U859 ( .A1(G1996), .A2(n982), .ZN(n840) );
  INV_X1 U860 ( .A(G1991), .ZN(n869) );
  NAND2_X1 U861 ( .A1(G131), .A2(n991), .ZN(n773) );
  NAND2_X1 U862 ( .A1(G119), .A2(n985), .ZN(n768) );
  NAND2_X1 U863 ( .A1(G107), .A2(n607), .ZN(n767) );
  NAND2_X1 U864 ( .A1(n768), .A2(n767), .ZN(n771) );
  NAND2_X1 U865 ( .A1(G95), .A2(n989), .ZN(n769) );
  XNOR2_X1 U866 ( .A(KEYINPUT93), .B(n769), .ZN(n770) );
  NOR2_X1 U867 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U868 ( .A1(n773), .A2(n772), .ZN(n774) );
  XOR2_X1 U869 ( .A(n774), .B(KEYINPUT94), .Z(n977) );
  NOR2_X1 U870 ( .A1(n869), .A2(n977), .ZN(n776) );
  AND2_X1 U871 ( .A1(n982), .A2(G1996), .ZN(n775) );
  OR2_X1 U872 ( .A1(n776), .A2(n775), .ZN(n838) );
  NOR2_X1 U873 ( .A1(n778), .A2(n777), .ZN(n799) );
  NAND2_X1 U874 ( .A1(n838), .A2(n799), .ZN(n797) );
  INV_X1 U875 ( .A(n797), .ZN(n781) );
  AND2_X1 U876 ( .A1(n869), .A2(n977), .ZN(n844) );
  NOR2_X1 U877 ( .A1(G1986), .A2(G290), .ZN(n779) );
  NOR2_X1 U878 ( .A1(n844), .A2(n779), .ZN(n780) );
  NOR2_X1 U879 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U880 ( .A1(n840), .A2(n782), .ZN(n783) );
  XNOR2_X1 U881 ( .A(n783), .B(KEYINPUT39), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G104), .A2(n989), .ZN(n785) );
  NAND2_X1 U883 ( .A1(G140), .A2(n991), .ZN(n784) );
  NAND2_X1 U884 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U885 ( .A(KEYINPUT34), .B(n786), .ZN(n791) );
  NAND2_X1 U886 ( .A1(G128), .A2(n985), .ZN(n788) );
  NAND2_X1 U887 ( .A1(G116), .A2(n607), .ZN(n787) );
  NAND2_X1 U888 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U889 ( .A(KEYINPUT35), .B(n789), .Z(n790) );
  NOR2_X1 U890 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U891 ( .A(KEYINPUT36), .B(n792), .ZN(n999) );
  XNOR2_X1 U892 ( .A(G2067), .B(KEYINPUT37), .ZN(n794) );
  NOR2_X1 U893 ( .A1(n999), .A2(n794), .ZN(n837) );
  NAND2_X1 U894 ( .A1(n799), .A2(n837), .ZN(n798) );
  NAND2_X1 U895 ( .A1(n793), .A2(n798), .ZN(n795) );
  NAND2_X1 U896 ( .A1(n999), .A2(n794), .ZN(n842) );
  NAND2_X1 U897 ( .A1(n795), .A2(n842), .ZN(n796) );
  NAND2_X1 U898 ( .A1(n796), .A2(n799), .ZN(n819) );
  INV_X1 U899 ( .A(n819), .ZN(n803) );
  NAND2_X1 U900 ( .A1(n798), .A2(n797), .ZN(n801) );
  XNOR2_X1 U901 ( .A(G1986), .B(G290), .ZN(n892) );
  AND2_X1 U902 ( .A1(n892), .A2(n799), .ZN(n800) );
  NOR2_X1 U903 ( .A1(n801), .A2(n800), .ZN(n802) );
  OR2_X1 U904 ( .A1(n803), .A2(n802), .ZN(n808) );
  AND2_X1 U905 ( .A1(n894), .A2(n808), .ZN(n805) );
  NAND2_X1 U906 ( .A1(n900), .A2(KEYINPUT33), .ZN(n804) );
  NAND2_X1 U907 ( .A1(n807), .A2(n806), .ZN(n824) );
  INV_X1 U908 ( .A(n808), .ZN(n822) );
  NOR2_X1 U909 ( .A1(G2090), .A2(G303), .ZN(n809) );
  NAND2_X1 U910 ( .A1(G8), .A2(n809), .ZN(n810) );
  NAND2_X1 U911 ( .A1(n811), .A2(n810), .ZN(n812) );
  AND2_X1 U912 ( .A1(n812), .A2(n815), .ZN(n818) );
  NOR2_X1 U913 ( .A1(G1981), .A2(G305), .ZN(n813) );
  XOR2_X1 U914 ( .A(n813), .B(KEYINPUT24), .Z(n814) );
  NOR2_X1 U915 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U916 ( .A(KEYINPUT97), .B(n816), .Z(n817) );
  NOR2_X1 U917 ( .A1(n818), .A2(n817), .ZN(n820) );
  AND2_X1 U918 ( .A1(n820), .A2(n819), .ZN(n821) );
  OR2_X2 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n826), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U924 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U926 ( .A1(n829), .A2(n828), .ZN(G188) );
  NAND2_X1 U928 ( .A1(G112), .A2(n607), .ZN(n831) );
  NAND2_X1 U929 ( .A1(G136), .A2(n991), .ZN(n830) );
  NAND2_X1 U930 ( .A1(n831), .A2(n830), .ZN(n836) );
  NAND2_X1 U931 ( .A1(G124), .A2(n985), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n832), .B(KEYINPUT44), .ZN(n834) );
  NAND2_X1 U933 ( .A1(n989), .A2(G100), .ZN(n833) );
  NAND2_X1 U934 ( .A1(n834), .A2(n833), .ZN(n835) );
  NOR2_X1 U935 ( .A1(n836), .A2(n835), .ZN(G162) );
  OR2_X1 U936 ( .A1(n838), .A2(n837), .ZN(n851) );
  XOR2_X1 U937 ( .A(G2090), .B(G162), .Z(n839) );
  NOR2_X1 U938 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U939 ( .A(KEYINPUT51), .B(n841), .Z(n849) );
  XNOR2_X1 U940 ( .A(G2084), .B(G160), .ZN(n843) );
  NAND2_X1 U941 ( .A1(n843), .A2(n842), .ZN(n847) );
  NOR2_X1 U942 ( .A1(n980), .A2(n844), .ZN(n845) );
  XNOR2_X1 U943 ( .A(KEYINPUT117), .B(n845), .ZN(n846) );
  NOR2_X1 U944 ( .A1(n847), .A2(n846), .ZN(n848) );
  NAND2_X1 U945 ( .A1(n849), .A2(n848), .ZN(n850) );
  NOR2_X1 U946 ( .A1(n851), .A2(n850), .ZN(n852) );
  XNOR2_X1 U947 ( .A(KEYINPUT118), .B(n852), .ZN(n866) );
  XOR2_X1 U948 ( .A(G164), .B(G2078), .Z(n863) );
  NAND2_X1 U949 ( .A1(G103), .A2(n989), .ZN(n854) );
  NAND2_X1 U950 ( .A1(G139), .A2(n991), .ZN(n853) );
  NAND2_X1 U951 ( .A1(n854), .A2(n853), .ZN(n860) );
  NAND2_X1 U952 ( .A1(G127), .A2(n985), .ZN(n856) );
  NAND2_X1 U953 ( .A1(G115), .A2(n607), .ZN(n855) );
  NAND2_X1 U954 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U955 ( .A(KEYINPUT47), .B(n857), .ZN(n858) );
  XNOR2_X1 U956 ( .A(KEYINPUT113), .B(n858), .ZN(n859) );
  NOR2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U958 ( .A(KEYINPUT114), .B(n861), .Z(n975) );
  XNOR2_X1 U959 ( .A(G2072), .B(n975), .ZN(n862) );
  NOR2_X1 U960 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U961 ( .A(KEYINPUT50), .B(n864), .ZN(n865) );
  NAND2_X1 U962 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U963 ( .A(KEYINPUT52), .B(n867), .ZN(n868) );
  NAND2_X1 U964 ( .A1(n868), .A2(G29), .ZN(n949) );
  XNOR2_X1 U965 ( .A(n869), .B(G25), .ZN(n870) );
  NAND2_X1 U966 ( .A1(n870), .A2(G28), .ZN(n871) );
  XNOR2_X1 U967 ( .A(n871), .B(KEYINPUT119), .ZN(n880) );
  XOR2_X1 U968 ( .A(G32), .B(G1996), .Z(n875) );
  XNOR2_X1 U969 ( .A(G2067), .B(G26), .ZN(n873) );
  XNOR2_X1 U970 ( .A(G2072), .B(G33), .ZN(n872) );
  NOR2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n874) );
  NAND2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n878) );
  XOR2_X1 U973 ( .A(G27), .B(n876), .Z(n877) );
  NOR2_X1 U974 ( .A1(n878), .A2(n877), .ZN(n879) );
  NAND2_X1 U975 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U976 ( .A(n881), .B(KEYINPUT53), .ZN(n884) );
  XOR2_X1 U977 ( .A(G2084), .B(G34), .Z(n882) );
  XNOR2_X1 U978 ( .A(KEYINPUT54), .B(n882), .ZN(n883) );
  NAND2_X1 U979 ( .A1(n884), .A2(n883), .ZN(n886) );
  XNOR2_X1 U980 ( .A(G35), .B(G2090), .ZN(n885) );
  NOR2_X1 U981 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U982 ( .A(n887), .B(KEYINPUT120), .ZN(n888) );
  NOR2_X1 U983 ( .A1(G29), .A2(n888), .ZN(n889) );
  XNOR2_X1 U984 ( .A(KEYINPUT55), .B(n889), .ZN(n890) );
  NAND2_X1 U985 ( .A1(n890), .A2(G11), .ZN(n947) );
  XNOR2_X1 U986 ( .A(G16), .B(KEYINPUT56), .ZN(n916) );
  XNOR2_X1 U987 ( .A(G1341), .B(n1004), .ZN(n891) );
  NOR2_X1 U988 ( .A1(n892), .A2(n891), .ZN(n914) );
  XOR2_X1 U989 ( .A(G1966), .B(G168), .Z(n893) );
  XNOR2_X1 U990 ( .A(KEYINPUT121), .B(n893), .ZN(n895) );
  NAND2_X1 U991 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n896), .B(KEYINPUT57), .ZN(n906) );
  XNOR2_X1 U993 ( .A(n897), .B(G1956), .ZN(n899) );
  XNOR2_X1 U994 ( .A(G166), .B(G1971), .ZN(n898) );
  NAND2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n904) );
  XNOR2_X1 U996 ( .A(KEYINPUT123), .B(n900), .ZN(n902) );
  NAND2_X1 U997 ( .A1(n902), .A2(n901), .ZN(n903) );
  NOR2_X1 U998 ( .A1(n904), .A2(n903), .ZN(n905) );
  NAND2_X1 U999 ( .A1(n906), .A2(n905), .ZN(n912) );
  XOR2_X1 U1000 ( .A(G171), .B(G1961), .Z(n909) );
  XNOR2_X1 U1001 ( .A(n907), .B(G1348), .ZN(n908) );
  NOR2_X1 U1002 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1003 ( .A(KEYINPUT122), .B(n910), .Z(n911) );
  NOR2_X1 U1004 ( .A1(n912), .A2(n911), .ZN(n913) );
  NAND2_X1 U1005 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1006 ( .A1(n916), .A2(n915), .ZN(n945) );
  INV_X1 U1007 ( .A(G16), .ZN(n943) );
  XNOR2_X1 U1008 ( .A(G5), .B(n917), .ZN(n938) );
  XNOR2_X1 U1009 ( .A(G1348), .B(KEYINPUT59), .ZN(n918) );
  XNOR2_X1 U1010 ( .A(n918), .B(G4), .ZN(n922) );
  XNOR2_X1 U1011 ( .A(G1981), .B(G6), .ZN(n920) );
  XNOR2_X1 U1012 ( .A(G1341), .B(G19), .ZN(n919) );
  NOR2_X1 U1013 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1014 ( .A1(n922), .A2(n921), .ZN(n926) );
  XOR2_X1 U1015 ( .A(G20), .B(n923), .Z(n924) );
  XNOR2_X1 U1016 ( .A(KEYINPUT124), .B(n924), .ZN(n925) );
  NOR2_X1 U1017 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1018 ( .A(n927), .B(KEYINPUT125), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(n928), .B(KEYINPUT60), .ZN(n936) );
  XNOR2_X1 U1020 ( .A(G1986), .B(G24), .ZN(n930) );
  XNOR2_X1 U1021 ( .A(G1971), .B(G22), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(n930), .A2(n929), .ZN(n933) );
  XOR2_X1 U1023 ( .A(G1976), .B(KEYINPUT126), .Z(n931) );
  XNOR2_X1 U1024 ( .A(G23), .B(n931), .ZN(n932) );
  NAND2_X1 U1025 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1026 ( .A(KEYINPUT58), .B(n934), .ZN(n935) );
  NOR2_X1 U1027 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1028 ( .A1(n938), .A2(n937), .ZN(n940) );
  XNOR2_X1 U1029 ( .A(G21), .B(G1966), .ZN(n939) );
  NOR2_X1 U1030 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1031 ( .A(KEYINPUT61), .B(n941), .ZN(n942) );
  NAND2_X1 U1032 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1033 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1034 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1035 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1036 ( .A(KEYINPUT62), .B(n950), .Z(G311) );
  XNOR2_X1 U1037 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1038 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1039 ( .A1(n952), .A2(n951), .ZN(G325) );
  INV_X1 U1040 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1041 ( .A(KEYINPUT108), .B(KEYINPUT41), .Z(n954) );
  XNOR2_X1 U1042 ( .A(G1981), .B(G1976), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(n954), .B(n953), .ZN(n955) );
  XOR2_X1 U1044 ( .A(n955), .B(KEYINPUT109), .Z(n957) );
  XNOR2_X1 U1045 ( .A(G1971), .B(G1956), .ZN(n956) );
  XNOR2_X1 U1046 ( .A(n957), .B(n956), .ZN(n961) );
  XOR2_X1 U1047 ( .A(G2474), .B(G1961), .Z(n959) );
  XNOR2_X1 U1048 ( .A(G1986), .B(G1966), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(n959), .B(n958), .ZN(n960) );
  XOR2_X1 U1050 ( .A(n961), .B(n960), .Z(n963) );
  XNOR2_X1 U1051 ( .A(G1996), .B(G1991), .ZN(n962) );
  XNOR2_X1 U1052 ( .A(n963), .B(n962), .ZN(G229) );
  XOR2_X1 U1053 ( .A(G2100), .B(G2096), .Z(n965) );
  XNOR2_X1 U1054 ( .A(G2067), .B(G2090), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(n965), .B(n964), .ZN(n969) );
  XOR2_X1 U1056 ( .A(G2678), .B(KEYINPUT42), .Z(n967) );
  XNOR2_X1 U1057 ( .A(G2072), .B(KEYINPUT43), .ZN(n966) );
  XNOR2_X1 U1058 ( .A(n967), .B(n966), .ZN(n968) );
  XOR2_X1 U1059 ( .A(n969), .B(n968), .Z(n971) );
  XNOR2_X1 U1060 ( .A(G2078), .B(G2084), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(n971), .B(n970), .ZN(G227) );
  INV_X1 U1062 ( .A(n972), .ZN(G319) );
  XOR2_X1 U1063 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n974) );
  XNOR2_X1 U1064 ( .A(G162), .B(KEYINPUT115), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(n974), .B(n973), .ZN(n976) );
  XOR2_X1 U1066 ( .A(n976), .B(n975), .Z(n979) );
  XOR2_X1 U1067 ( .A(G164), .B(n977), .Z(n978) );
  XNOR2_X1 U1068 ( .A(n979), .B(n978), .ZN(n981) );
  XOR2_X1 U1069 ( .A(n981), .B(n980), .Z(n984) );
  XOR2_X1 U1070 ( .A(G160), .B(n982), .Z(n983) );
  XNOR2_X1 U1071 ( .A(n984), .B(n983), .ZN(n1001) );
  NAND2_X1 U1072 ( .A1(n985), .A2(G130), .ZN(n986) );
  XNOR2_X1 U1073 ( .A(n986), .B(KEYINPUT110), .ZN(n988) );
  NAND2_X1 U1074 ( .A1(G118), .A2(n607), .ZN(n987) );
  NAND2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n997) );
  NAND2_X1 U1076 ( .A1(n989), .A2(G106), .ZN(n990) );
  XOR2_X1 U1077 ( .A(KEYINPUT111), .B(n990), .Z(n993) );
  NAND2_X1 U1078 ( .A1(n991), .A2(G142), .ZN(n992) );
  NAND2_X1 U1079 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1080 ( .A(KEYINPUT112), .B(n994), .Z(n995) );
  XNOR2_X1 U1081 ( .A(KEYINPUT45), .B(n995), .ZN(n996) );
  NOR2_X1 U1082 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1083 ( .A(n999), .B(n998), .ZN(n1000) );
  XNOR2_X1 U1084 ( .A(n1001), .B(n1000), .ZN(n1002) );
  NOR2_X1 U1085 ( .A1(G37), .A2(n1002), .ZN(G395) );
  XNOR2_X1 U1086 ( .A(n1004), .B(n1003), .ZN(n1007) );
  XNOR2_X1 U1087 ( .A(G171), .B(n1005), .ZN(n1006) );
  XNOR2_X1 U1088 ( .A(n1007), .B(n1006), .ZN(n1008) );
  XNOR2_X1 U1089 ( .A(G286), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1090 ( .A1(G37), .A2(n1009), .ZN(G397) );
  XNOR2_X1 U1091 ( .A(KEYINPUT49), .B(KEYINPUT116), .ZN(n1011) );
  NOR2_X1 U1092 ( .A1(G229), .A2(G227), .ZN(n1010) );
  XNOR2_X1 U1093 ( .A(n1011), .B(n1010), .ZN(n1022) );
  XOR2_X1 U1094 ( .A(G2446), .B(G2451), .Z(n1013) );
  XNOR2_X1 U1095 ( .A(G1348), .B(G2430), .ZN(n1012) );
  XNOR2_X1 U1096 ( .A(n1013), .B(n1012), .ZN(n1019) );
  XOR2_X1 U1097 ( .A(G2443), .B(G2438), .Z(n1015) );
  XNOR2_X1 U1098 ( .A(G2454), .B(G2435), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(n1015), .B(n1014), .ZN(n1017) );
  XOR2_X1 U1100 ( .A(G1341), .B(G2427), .Z(n1016) );
  XNOR2_X1 U1101 ( .A(n1017), .B(n1016), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(n1019), .B(n1018), .Z(n1020) );
  NAND2_X1 U1103 ( .A1(G14), .A2(n1020), .ZN(n1025) );
  NAND2_X1 U1104 ( .A1(G319), .A2(n1025), .ZN(n1021) );
  NOR2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  NOR2_X1 U1106 ( .A1(G395), .A2(G397), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1024), .A2(n1023), .ZN(G225) );
  INV_X1 U1108 ( .A(G225), .ZN(G308) );
  INV_X1 U1109 ( .A(G108), .ZN(G238) );
  INV_X1 U1110 ( .A(n1025), .ZN(G401) );
endmodule

