//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1294, new_n1295, new_n1297,
    new_n1298, new_n1299, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1373, new_n1374, new_n1375, new_n1376;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0006(.A1(G58), .A2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n212), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n214), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n217), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n222), .B(new_n230), .C1(new_n219), .C2(new_n221), .ZN(G361));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(KEYINPUT66), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n236), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n211), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n212), .A2(G33), .A3(G77), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n254), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n252), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT11), .ZN(new_n257));
  OR2_X1    g0057(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n215), .A2(G13), .A3(G20), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n258), .B(new_n259), .C1(new_n260), .C2(G68), .ZN(new_n261));
  INV_X1    g0061(.A(new_n260), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n203), .ZN(new_n263));
  OAI211_X1 g0063(.A(KEYINPUT72), .B(new_n261), .C1(new_n263), .C2(KEYINPUT12), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n262), .A2(new_n251), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n212), .A2(G1), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(G68), .A3(new_n267), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n264), .B(new_n268), .C1(KEYINPUT72), .C2(new_n261), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n257), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT74), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT74), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(new_n257), .B2(new_n269), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT14), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G1), .A3(G13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n281), .A3(G274), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n215), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n281), .A2(G238), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G226), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n238), .A2(G1698), .ZN(new_n290));
  AND2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR2_X1   g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n289), .B(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G97), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n281), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n276), .B1(new_n286), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n281), .B1(new_n293), .B2(new_n294), .ZN(new_n299));
  INV_X1    g0099(.A(new_n276), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n299), .A2(new_n285), .A3(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n275), .B(G169), .C1(new_n298), .C2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n286), .A2(new_n297), .A3(new_n276), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT13), .B1(new_n299), .B2(new_n285), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(G179), .A3(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT73), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n300), .B1(new_n299), .B2(new_n285), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n275), .B1(new_n309), .B2(G169), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n306), .A2(new_n307), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n302), .A2(new_n305), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT73), .B1(new_n313), .B2(new_n310), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n274), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n303), .A2(G190), .A3(new_n304), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n270), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n298), .A2(new_n301), .ZN(new_n318));
  INV_X1    g0118(.A(G200), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  OR2_X1    g0122(.A1(KEYINPUT3), .A2(G33), .ZN(new_n323));
  NAND2_X1  g0123(.A1(KEYINPUT3), .A2(G33), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n288), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n291), .A2(new_n292), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n325), .A2(G223), .B1(new_n326), .B2(G77), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT3), .B(G33), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n328), .A2(G222), .A3(new_n288), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n296), .ZN(new_n331));
  INV_X1    g0131(.A(new_n282), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n296), .A2(new_n279), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(G226), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G200), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n204), .A2(G20), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n254), .A2(G150), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n212), .A2(G33), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT8), .B(G58), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n337), .B(new_n338), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(new_n251), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n266), .A2(new_n201), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n265), .A2(new_n343), .B1(new_n201), .B2(new_n262), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT9), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n331), .A2(G190), .A3(new_n334), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n342), .A2(KEYINPUT9), .A3(new_n344), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n336), .A2(new_n347), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT10), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n347), .A2(new_n349), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT10), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n352), .A2(new_n353), .A3(new_n348), .A4(new_n336), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n335), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n345), .B1(new_n356), .B2(G169), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n335), .A2(G179), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n332), .B1(G244), .B2(new_n333), .ZN(new_n360));
  OAI211_X1 g0160(.A(G238), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n323), .A2(G107), .A3(new_n324), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(G232), .B(new_n288), .C1(new_n291), .C2(new_n292), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT67), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT67), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n328), .A2(new_n366), .A3(G232), .A4(new_n288), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n296), .B1(new_n368), .B2(KEYINPUT68), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n365), .A2(new_n367), .ZN(new_n370));
  INV_X1    g0170(.A(new_n363), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n370), .A2(KEYINPUT68), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n360), .B1(new_n369), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G200), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n265), .A2(G77), .A3(new_n267), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(G77), .B2(new_n260), .ZN(new_n376));
  INV_X1    g0176(.A(new_n340), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(new_n254), .B1(G20), .B2(G77), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT15), .B(G87), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n378), .B1(new_n339), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n376), .B1(new_n380), .B2(new_n251), .ZN(new_n381));
  INV_X1    g0181(.A(G190), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n374), .B(new_n381), .C1(new_n382), .C2(new_n373), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n355), .A2(new_n359), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n360), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n370), .A2(new_n371), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT68), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n281), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n368), .A2(KEYINPUT68), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(G169), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT69), .B1(new_n391), .B2(new_n381), .ZN(new_n392));
  INV_X1    g0192(.A(G169), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n381), .B1(new_n373), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT69), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G179), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n390), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n392), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n340), .A2(new_n266), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n400), .A2(new_n265), .B1(new_n340), .B2(new_n262), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(KEYINPUT7), .B1(new_n326), .B2(new_n212), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  NOR4_X1   g0204(.A1(new_n291), .A2(new_n292), .A3(new_n404), .A4(G20), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n202), .A2(new_n203), .ZN(new_n407));
  OAI21_X1  g0207(.A(G20), .B1(new_n407), .B2(new_n207), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n254), .A2(G159), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n252), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n406), .A2(KEYINPUT16), .A3(new_n411), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n402), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OR2_X1    g0216(.A1(G223), .A2(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n287), .A2(G1698), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n291), .C2(new_n292), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G87), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n281), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n281), .A2(G232), .A3(new_n283), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n282), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n422), .A2(new_n425), .A3(new_n397), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n393), .B1(new_n421), .B2(new_n424), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT18), .B1(new_n416), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n404), .B1(new_n328), .B2(G20), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n326), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n203), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n413), .B1(new_n432), .B2(new_n410), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(new_n415), .A3(new_n251), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n428), .B1(new_n434), .B2(new_n401), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n422), .A2(new_n425), .A3(new_n382), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n319), .B1(new_n421), .B2(new_n424), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n434), .A2(new_n401), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n434), .A2(new_n440), .A3(KEYINPUT17), .A4(new_n401), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n429), .A2(new_n437), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n322), .A2(new_n384), .A3(new_n399), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT75), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n355), .A2(new_n359), .A3(new_n383), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n445), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT75), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n450), .A2(new_n451), .A3(new_n399), .A4(new_n322), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(G244), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT80), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT80), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n328), .A2(new_n456), .A3(G244), .A4(G1698), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G116), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n328), .A2(G238), .A3(new_n288), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n455), .A2(new_n457), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n296), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n278), .A2(G1), .ZN(new_n462));
  INV_X1    g0262(.A(G274), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G250), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n278), .B2(G1), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n281), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(KEYINPUT83), .B1(new_n468), .B2(new_n382), .ZN(new_n469));
  INV_X1    g0269(.A(new_n467), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n460), .B2(new_n296), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT83), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n471), .A2(new_n472), .A3(G190), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n468), .A2(G200), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT19), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n212), .B1(new_n294), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(G97), .A2(G107), .ZN(new_n478));
  INV_X1    g0278(.A(G87), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n212), .B(G68), .C1(new_n291), .C2(new_n292), .ZN(new_n482));
  INV_X1    g0282(.A(G97), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n476), .B1(new_n339), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n251), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n379), .A2(new_n262), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n215), .A2(G33), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n260), .A2(new_n488), .A3(new_n211), .A4(new_n250), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G87), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n486), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n475), .A2(KEYINPUT82), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT82), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n471), .A2(new_n319), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n485), .A2(new_n251), .B1(new_n379), .B2(new_n262), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n491), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n494), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n474), .A2(new_n493), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n468), .A2(G169), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT81), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n461), .A2(G179), .A3(new_n467), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n471), .A2(new_n393), .ZN(new_n504));
  AOI211_X1 g0304(.A(new_n397), .B(new_n470), .C1(new_n460), .C2(new_n296), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT81), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n379), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n490), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n496), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n503), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  AND2_X1   g0310(.A1(new_n499), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n262), .A2(new_n483), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n489), .B2(new_n483), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(G107), .B1(new_n403), .B2(new_n405), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT6), .ZN(new_n516));
  AND2_X1   g0316(.A1(G97), .A2(G107), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n517), .B2(new_n478), .ZN(new_n518));
  INV_X1    g0318(.A(G107), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n519), .A2(KEYINPUT6), .A3(G97), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(G20), .B1(G77), .B2(new_n254), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n252), .B1(new_n515), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n523), .A2(KEYINPUT76), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT76), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n525), .B(new_n252), .C1(new_n515), .C2(new_n522), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n514), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT78), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n528), .A2(new_n277), .A3(KEYINPUT5), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT5), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G41), .ZN(new_n531));
  AND3_X1   g0331(.A1(new_n529), .A2(new_n462), .A3(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT79), .ZN(new_n533));
  INV_X1    g0333(.A(new_n211), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n463), .B1(new_n534), .B2(new_n280), .ZN(new_n535));
  OAI21_X1  g0335(.A(KEYINPUT78), .B1(new_n530), .B2(G41), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n532), .A2(new_n533), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n536), .A2(new_n529), .A3(new_n462), .A4(new_n531), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n281), .A2(G274), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT79), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n277), .A2(KEYINPUT5), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n462), .A2(new_n541), .A3(new_n531), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n542), .A2(new_n281), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n537), .A2(new_n540), .B1(G257), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G244), .B(new_n288), .C1(new_n291), .C2(new_n292), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G250), .A2(G1698), .ZN(new_n548));
  NAND2_X1  g0348(.A1(KEYINPUT4), .A2(G244), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n548), .B1(new_n549), .B2(G1698), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n328), .A2(new_n550), .B1(G33), .B2(G283), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT77), .B1(new_n552), .B2(new_n296), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT77), .ZN(new_n554));
  AOI211_X1 g0354(.A(new_n554), .B(new_n281), .C1(new_n547), .C2(new_n551), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n397), .B(new_n544), .C1(new_n553), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n552), .A2(new_n296), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n537), .A2(new_n540), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n543), .A2(G257), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n393), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n527), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n544), .B1(new_n553), .B2(new_n555), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G200), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n254), .A2(G77), .ZN(new_n565));
  INV_X1    g0365(.A(new_n520), .ZN(new_n566));
  XNOR2_X1  g0366(.A(G97), .B(G107), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n566), .B1(new_n516), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n565), .B1(new_n568), .B2(new_n212), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n519), .B1(new_n430), .B2(new_n431), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n251), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(new_n525), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n523), .A2(KEYINPUT76), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n544), .A2(G190), .A3(new_n557), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n564), .A2(new_n574), .A3(new_n514), .A4(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(G13), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(G1), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT25), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n578), .A2(new_n579), .A3(G20), .A4(new_n519), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT25), .B1(new_n260), .B2(G107), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n581), .C1(new_n489), .C2(new_n519), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT86), .ZN(new_n583));
  XNOR2_X1  g0383(.A(new_n582), .B(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT23), .B1(new_n212), .B2(G107), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT23), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(new_n519), .A3(G20), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n212), .A2(G33), .A3(G116), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT85), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n585), .A2(new_n587), .A3(new_n588), .A4(KEYINPUT85), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n212), .B(G87), .C1(new_n291), .C2(new_n292), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT22), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT22), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n328), .A2(new_n596), .A3(new_n212), .A4(G87), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT24), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n252), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n591), .A2(new_n592), .B1(new_n595), .B2(new_n597), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT24), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n584), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n215), .B(G45), .C1(new_n277), .C2(KEYINPUT5), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n530), .A2(G41), .ZN(new_n606));
  OAI211_X1 g0406(.A(G264), .B(new_n281), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT87), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n542), .A2(KEYINPUT87), .A3(G264), .A4(new_n281), .ZN(new_n610));
  OAI211_X1 g0410(.A(G257), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n611));
  OAI211_X1 g0411(.A(G250), .B(new_n288), .C1(new_n291), .C2(new_n292), .ZN(new_n612));
  NAND2_X1  g0412(.A1(G33), .A2(G294), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n609), .A2(new_n610), .B1(new_n614), .B2(new_n296), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n615), .A2(G190), .A3(new_n558), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n609), .A2(new_n610), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n296), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n558), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G200), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n604), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n562), .A2(new_n576), .A3(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(G257), .B(new_n288), .C1(new_n291), .C2(new_n292), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n323), .A2(G303), .A3(new_n324), .ZN(new_n624));
  OAI211_X1 g0424(.A(G264), .B(G1698), .C1(new_n291), .C2(new_n292), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(KEYINPUT84), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT84), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n325), .B2(G264), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n296), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n543), .A2(G270), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n558), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G200), .ZN(new_n632));
  NAND2_X1  g0432(.A1(G33), .A2(G283), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n633), .B(new_n212), .C1(G33), .C2(new_n483), .ZN(new_n634));
  INV_X1    g0434(.A(G116), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(G20), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n251), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT20), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n634), .A2(KEYINPUT20), .A3(new_n251), .A4(new_n636), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n260), .A2(G116), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n490), .B2(G116), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n632), .B(new_n644), .C1(new_n382), .C2(new_n631), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n393), .B1(new_n641), .B2(new_n643), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n631), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT21), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT21), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n631), .A2(new_n649), .A3(new_n646), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n582), .B(KEYINPUT86), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n251), .B1(new_n602), .B2(KEYINPUT24), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n599), .A2(new_n600), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n619), .A2(new_n393), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n615), .A2(new_n397), .A3(new_n558), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n644), .A2(new_n397), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n629), .A2(new_n558), .A3(new_n630), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND4_X1   g0461(.A1(new_n645), .A2(new_n651), .A3(new_n658), .A4(new_n661), .ZN(new_n662));
  AND4_X1   g0462(.A1(new_n453), .A2(new_n511), .A3(new_n622), .A4(new_n662), .ZN(G372));
  INV_X1    g0463(.A(new_n359), .ZN(new_n664));
  INV_X1    g0464(.A(new_n274), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n307), .B1(new_n306), .B2(new_n311), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n313), .A2(new_n310), .A3(KEYINPUT73), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n399), .B2(new_n321), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n443), .A2(new_n444), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  AOI211_X1 g0472(.A(KEYINPUT18), .B(new_n428), .C1(new_n434), .C2(new_n401), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n434), .A2(new_n401), .ZN(new_n674));
  INV_X1    g0474(.A(new_n428), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n436), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n664), .B1(new_n678), .B2(new_n355), .ZN(new_n679));
  INV_X1    g0479(.A(new_n453), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT26), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n509), .B1(new_n504), .B2(new_n505), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n492), .B(KEYINPUT88), .C1(new_n471), .C2(new_n319), .ZN(new_n683));
  AND4_X1   g0483(.A1(new_n472), .A2(new_n461), .A3(G190), .A4(new_n467), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n472), .B1(new_n471), .B2(G190), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT88), .B1(new_n475), .B2(new_n492), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n682), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n681), .B1(new_n688), .B2(new_n562), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n513), .B1(new_n572), .B2(new_n573), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n556), .A2(new_n561), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g0492(.A(KEYINPUT89), .B(KEYINPUT26), .Z(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n499), .A2(new_n510), .A3(new_n692), .A4(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n651), .A2(new_n658), .A3(new_n661), .ZN(new_n697));
  INV_X1    g0497(.A(new_n688), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n622), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(new_n699), .A3(new_n682), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n679), .B1(new_n680), .B2(new_n701), .ZN(G369));
  INV_X1    g0502(.A(new_n645), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n631), .A2(new_n649), .A3(new_n646), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n649), .B1(new_n631), .B2(new_n646), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n661), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n578), .A2(new_n212), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT27), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT27), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(G213), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G343), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n644), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n706), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n706), .A2(new_n713), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n703), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n656), .A2(new_n657), .ZN(new_n718));
  INV_X1    g0518(.A(new_n712), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n718), .A2(new_n604), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n621), .B1(new_n604), .B2(new_n712), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n658), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n717), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n706), .A2(new_n712), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT90), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n706), .A2(KEYINPUT90), .A3(new_n712), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n720), .B1(new_n730), .B2(new_n722), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n725), .A2(new_n731), .ZN(G399));
  INV_X1    g0532(.A(new_n218), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G41), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n480), .A2(G116), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(G1), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n209), .B2(new_n735), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT28), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT29), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n700), .A2(new_n740), .A3(new_n712), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n499), .A2(new_n510), .A3(new_n692), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n693), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT88), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n495), .B2(new_n497), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n474), .A2(new_n746), .A3(new_n683), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n747), .A2(new_n692), .A3(KEYINPUT26), .A4(new_n682), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(new_n682), .A3(new_n699), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n740), .B1(new_n750), .B2(new_n712), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n742), .A2(new_n751), .ZN(new_n752));
  AND4_X1   g0552(.A1(KEYINPUT30), .A2(new_n557), .A3(new_n558), .A4(new_n559), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n753), .A2(new_n660), .A3(new_n505), .A4(new_n615), .ZN(new_n754));
  AOI21_X1  g0554(.A(G179), .B1(new_n615), .B2(new_n558), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n563), .A2(new_n468), .A3(new_n631), .A4(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n615), .A2(new_n629), .A3(new_n558), .A4(new_n630), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n757), .A2(new_n502), .A3(new_n560), .ZN(new_n758));
  XNOR2_X1  g0558(.A(KEYINPUT91), .B(KEYINPUT30), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n754), .B(new_n756), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n719), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT31), .B1(new_n760), .B2(new_n719), .ZN(new_n762));
  OAI21_X1  g0562(.A(KEYINPUT92), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n760), .A2(new_n719), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT31), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT92), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n760), .A2(KEYINPUT31), .A3(new_n719), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n511), .A2(new_n622), .A3(new_n662), .A4(new_n712), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n763), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G330), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n752), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n739), .B1(new_n773), .B2(G1), .ZN(G364));
  INV_X1    g0574(.A(new_n717), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n716), .A2(G330), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n577), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n215), .B1(new_n777), .B2(G45), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n734), .A2(new_n779), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n775), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G13), .A2(G33), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(G20), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n716), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n733), .A2(new_n326), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G355), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(G116), .B2(new_n218), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n733), .A2(new_n328), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n278), .B2(new_n210), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n245), .A2(new_n278), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n789), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n211), .B1(G20), .B2(new_n393), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n784), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n780), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(G20), .A2(G179), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G190), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G200), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G322), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n212), .A2(G179), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n805), .A2(new_n382), .A3(G200), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n803), .A2(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n382), .A2(G179), .A3(G200), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n212), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n808), .B1(G294), .B2(new_n811), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n799), .A2(new_n319), .A3(G190), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(KEYINPUT33), .B(G317), .Z(new_n815));
  NOR2_X1   g0615(.A1(G190), .A2(G200), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n800), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n814), .A2(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n805), .A2(new_n816), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n328), .B(new_n819), .C1(G329), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n801), .A2(new_n319), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n805), .A2(G190), .A3(G200), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G326), .A2(new_n823), .B1(new_n825), .B2(G303), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n812), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n806), .A2(new_n519), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n326), .B(new_n828), .C1(G87), .C2(new_n825), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT93), .Z(new_n830));
  INV_X1    g0630(.A(KEYINPUT32), .ZN(new_n831));
  INV_X1    g0631(.A(G159), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n820), .A2(new_n832), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n803), .A2(new_n202), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n823), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n835), .A2(new_n201), .B1(new_n483), .B2(new_n810), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n833), .A2(new_n831), .ZN(new_n838));
  INV_X1    g0638(.A(new_n817), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n839), .A2(G77), .B1(G68), .B2(new_n813), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n827), .B1(new_n830), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n798), .B1(new_n842), .B2(new_n795), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n781), .B1(new_n786), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G396));
  INV_X1    g0645(.A(new_n780), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n795), .A2(new_n782), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT94), .Z(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(G77), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n820), .A2(new_n818), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n326), .B1(new_n817), .B2(new_n635), .ZN(new_n853));
  AOI211_X1 g0653(.A(new_n852), .B(new_n853), .C1(G283), .C2(new_n813), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n802), .A2(G294), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n806), .A2(new_n479), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(G107), .B2(new_n825), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n811), .A2(G97), .B1(new_n823), .B2(G303), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n854), .A2(new_n855), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT95), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n328), .B1(new_n820), .B2(new_n861), .C1(new_n201), .C2(new_n824), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n810), .A2(new_n202), .B1(new_n806), .B2(new_n203), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n839), .A2(G159), .B1(G150), .B2(new_n813), .ZN(new_n864));
  INV_X1    g0664(.A(G143), .ZN(new_n865));
  INV_X1    g0665(.A(G137), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n864), .B1(new_n803), .B2(new_n865), .C1(new_n866), .C2(new_n835), .ZN(new_n867));
  XOR2_X1   g0667(.A(new_n867), .B(KEYINPUT34), .Z(new_n868));
  AOI211_X1 g0668(.A(new_n862), .B(new_n863), .C1(new_n868), .C2(KEYINPUT96), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n868), .A2(KEYINPUT96), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n795), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n381), .A2(new_n712), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n381), .B1(new_n373), .B2(new_n382), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n390), .A2(new_n319), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n398), .B1(new_n394), .B2(new_n395), .ZN(new_n877));
  AOI211_X1 g0677(.A(KEYINPUT69), .B(new_n381), .C1(new_n373), .C2(new_n393), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n392), .A2(new_n396), .A3(new_n398), .A4(new_n873), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n851), .B1(new_n871), .B2(new_n872), .C1(new_n882), .C2(new_n783), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n700), .B2(new_n712), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n879), .A2(new_n880), .A3(new_n712), .ZN(new_n885));
  INV_X1    g0685(.A(new_n682), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n562), .A2(new_n576), .A3(new_n621), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n718), .A2(new_n604), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n706), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n886), .B1(new_n890), .B2(new_n698), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n885), .B1(new_n891), .B2(new_n696), .ZN(new_n892));
  OR2_X1    g0692(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n893), .A2(new_n772), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT97), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(new_n846), .C1(new_n772), .C2(new_n893), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n894), .A2(KEYINPUT97), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n883), .B1(new_n896), .B2(new_n897), .ZN(G384));
  OR2_X1    g0698(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n521), .A2(KEYINPUT35), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n899), .A2(G116), .A3(new_n213), .A4(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(KEYINPUT36), .Z(new_n902));
  OR3_X1    g0702(.A1(new_n209), .A2(new_n850), .A3(new_n407), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n201), .A2(G68), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n215), .B(G13), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n321), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n274), .A2(new_n712), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n668), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n315), .B2(new_n321), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n399), .A2(new_n719), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n912), .B1(new_n892), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT98), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n441), .B1(new_n416), .B2(new_n428), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n416), .A2(new_n710), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT37), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n674), .A2(new_n675), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n674), .A2(new_n711), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT37), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .A4(new_n441), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n445), .A2(new_n917), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT38), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT38), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n915), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT38), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n434), .A2(new_n401), .A3(new_n440), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n929), .A2(new_n435), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n921), .B1(new_n930), .B2(new_n920), .ZN(new_n931));
  AND4_X1   g0731(.A1(new_n921), .A2(new_n919), .A3(new_n920), .A4(new_n441), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n920), .B1(new_n671), .B2(new_n677), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n928), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT38), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(KEYINPUT98), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n914), .B1(new_n927), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n925), .B2(new_n926), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n935), .A2(KEYINPUT39), .A3(new_n936), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n315), .A2(new_n712), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT99), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n943), .B(new_n944), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n942), .A2(new_n945), .B1(new_n677), .B2(new_n711), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n453), .B1(new_n742), .B2(new_n751), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n948), .A2(new_n679), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n947), .B(new_n949), .Z(new_n950));
  AOI21_X1  g0750(.A(new_n881), .B1(new_n910), .B2(new_n911), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n761), .A2(new_n762), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n770), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(new_n927), .B2(new_n937), .ZN(new_n955));
  OAI21_X1  g0755(.A(KEYINPUT40), .B1(new_n925), .B2(new_n926), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n955), .A2(KEYINPUT40), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n453), .A2(new_n953), .ZN(new_n958));
  OAI21_X1  g0758(.A(G330), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n950), .A2(new_n960), .B1(new_n215), .B2(new_n777), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n950), .A2(new_n960), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n906), .B1(new_n961), .B2(new_n962), .ZN(G367));
  OAI21_X1  g0763(.A(new_n698), .B1(new_n492), .B2(new_n712), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n886), .A2(new_n497), .A3(new_n719), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT100), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(KEYINPUT100), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n968), .A2(new_n785), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n236), .A2(new_n790), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n796), .B1(new_n218), .B2(new_n379), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n780), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n824), .A2(new_n635), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n973), .A2(KEYINPUT46), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT107), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n326), .B1(new_n817), .B2(new_n807), .ZN(new_n976));
  INV_X1    g0776(.A(G294), .ZN(new_n977));
  INV_X1    g0777(.A(G317), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n814), .A2(new_n977), .B1(new_n820), .B2(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n976), .B(new_n979), .C1(KEYINPUT46), .C2(new_n973), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n811), .A2(G107), .B1(new_n823), .B2(G311), .ZN(new_n981));
  INV_X1    g0781(.A(new_n806), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G303), .A2(new_n802), .B1(new_n982), .B2(G97), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n975), .A2(new_n980), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n835), .A2(new_n865), .B1(new_n824), .B2(new_n202), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(G150), .B2(new_n802), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n820), .A2(new_n866), .B1(new_n817), .B2(new_n201), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n326), .B(new_n987), .C1(G159), .C2(new_n813), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n806), .A2(new_n850), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G68), .B2(new_n811), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n984), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n972), .B1(new_n993), .B2(new_n795), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n969), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n723), .A2(new_n728), .A3(new_n729), .ZN(new_n996));
  INV_X1    g0796(.A(new_n729), .ZN(new_n997));
  AOI21_X1  g0797(.A(KEYINPUT90), .B1(new_n706), .B2(new_n712), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n722), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AND3_X1   g0799(.A1(new_n996), .A2(new_n775), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n775), .B1(new_n996), .B2(new_n999), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n1002), .A2(new_n752), .A3(new_n772), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n720), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n562), .B(new_n576), .C1(new_n690), .C2(new_n712), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n692), .A2(new_n719), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n999), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT45), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n731), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n999), .A2(new_n1004), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1007), .ZN(new_n1014));
  XOR2_X1   g0814(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n1015));
  NAND3_X1  g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1015), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n731), .B2(new_n1007), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1012), .A2(KEYINPUT104), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT105), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n725), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1022));
  AOI21_X1  g0822(.A(KEYINPUT45), .B1(new_n731), .B2(new_n1007), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1016), .B(new_n1018), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(KEYINPUT104), .B1(new_n724), .B2(KEYINPUT105), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1003), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n773), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n734), .B(KEYINPUT41), .Z(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT106), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1028), .A2(KEYINPUT106), .A3(new_n1030), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n779), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n999), .A2(new_n1014), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT42), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n968), .A2(KEYINPUT101), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n968), .A2(KEYINPUT101), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1038), .A2(new_n1039), .A3(KEYINPUT43), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n576), .A2(new_n888), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n712), .B1(new_n1041), .B2(new_n692), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1037), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT102), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n725), .A2(new_n1014), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1040), .B1(KEYINPUT43), .B2(new_n968), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1037), .A2(new_n1042), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1044), .A2(new_n1045), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1045), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n995), .B1(new_n1035), .B2(new_n1052), .ZN(G387));
  NOR2_X1   g0853(.A1(new_n824), .A2(new_n850), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n810), .A2(new_n379), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1054), .B(new_n1055), .C1(G50), .C2(new_n802), .ZN(new_n1056));
  INV_X1    g0856(.A(G150), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n820), .A2(new_n1057), .B1(new_n817), .B2(new_n203), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n326), .B(new_n1058), .C1(new_n377), .C2(new_n813), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G159), .A2(new_n823), .B1(new_n982), .B2(G97), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1056), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n328), .B1(new_n821), .B2(G326), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n810), .A2(new_n807), .B1(new_n824), .B2(new_n977), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n839), .A2(G303), .B1(G311), .B2(new_n813), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n803), .B2(new_n978), .C1(new_n804), .C2(new_n835), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n1066), .B2(new_n1065), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT49), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1062), .B1(new_n635), .B2(new_n806), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1061), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n795), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n736), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n787), .A2(new_n1074), .B1(new_n519), .B2(new_n733), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n241), .A2(new_n278), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n377), .A2(new_n201), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT50), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n736), .B(new_n278), .C1(new_n203), .C2(new_n850), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n790), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1075), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n846), .B1(new_n1081), .B2(new_n796), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1073), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n723), .B2(new_n784), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1002), .B2(new_n779), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n773), .A2(new_n1002), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n734), .B(KEYINPUT108), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n752), .A2(new_n772), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1087), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1085), .B1(new_n1086), .B2(new_n1090), .ZN(G393));
  NAND3_X1  g0891(.A1(new_n1024), .A2(KEYINPUT109), .A3(new_n724), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n724), .B2(new_n1024), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT109), .B1(new_n1024), .B2(new_n724), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1027), .B(new_n1087), .C1(new_n1095), .C2(new_n1003), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G311), .A2(new_n802), .B1(new_n823), .B2(G317), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT52), .Z(new_n1098));
  NAND2_X1  g0898(.A1(new_n813), .A2(G303), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n810), .B2(new_n635), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n1100), .A2(KEYINPUT110), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(KEYINPUT110), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n326), .B1(new_n817), .B2(new_n977), .C1(new_n804), .C2(new_n820), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n828), .B(new_n1103), .C1(G283), .C2(new_n825), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1098), .A2(new_n1101), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT111), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G150), .A2(new_n823), .B1(new_n802), .B2(G159), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT51), .Z(new_n1109));
  OAI22_X1  g0909(.A1(new_n817), .A2(new_n340), .B1(new_n820), .B2(new_n865), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n326), .B(new_n1110), .C1(G50), .C2(new_n813), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n810), .A2(new_n850), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n856), .B(new_n1112), .C1(G68), .C2(new_n825), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1109), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1107), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n795), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n796), .B1(new_n483), .B2(new_n218), .C1(new_n791), .C2(new_n248), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1117), .A2(new_n780), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n784), .B2(new_n1014), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n1095), .B2(new_n779), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1096), .A2(new_n1121), .ZN(G390));
  NAND2_X1  g0922(.A1(new_n942), .A2(new_n782), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n803), .A2(new_n635), .B1(new_n835), .B2(new_n807), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1112), .B(new_n1124), .C1(G68), .C2(new_n982), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n326), .B1(new_n820), .B2(new_n977), .C1(new_n479), .C2(new_n824), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n814), .A2(new_n519), .B1(new_n817), .B2(new_n483), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(KEYINPUT114), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1125), .B(new_n1128), .C1(KEYINPUT114), .C2(new_n1127), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT54), .B(G143), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n814), .A2(new_n866), .B1(new_n817), .B2(new_n1130), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n326), .B(new_n1131), .C1(G125), .C2(new_n821), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n824), .A2(new_n1057), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT53), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G132), .A2(new_n802), .B1(new_n982), .B2(G50), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n811), .A2(G159), .B1(new_n823), .B2(G128), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n872), .B1(new_n1129), .B2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n846), .B(new_n1138), .C1(new_n340), .C2(new_n849), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1123), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n885), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n913), .B1(new_n700), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n912), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n945), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n942), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n771), .A2(new_n951), .A3(G330), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(KEYINPUT112), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT112), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n771), .A2(new_n951), .A3(new_n1148), .A4(G330), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n935), .A2(new_n936), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1151), .A2(new_n945), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n719), .B1(new_n891), .B2(new_n749), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n913), .B1(new_n1153), .B2(new_n882), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1152), .B1(new_n1154), .B2(new_n1143), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1145), .A2(new_n1150), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT113), .ZN(new_n1157));
  INV_X1    g0957(.A(G330), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n952), .B2(new_n770), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1159), .A2(new_n951), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n914), .A2(new_n945), .B1(new_n940), .B2(new_n941), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1151), .A2(new_n945), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n913), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n697), .A2(new_n562), .A3(new_n576), .A4(new_n621), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n682), .B1(new_n1164), .B2(new_n688), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n688), .A2(new_n562), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1166), .A2(KEYINPUT26), .B1(new_n743), .B2(new_n693), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n712), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1163), .B1(new_n1168), .B2(new_n881), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1162), .B1(new_n1169), .B2(new_n912), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1160), .B1(new_n1161), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT113), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1145), .A2(new_n1150), .A3(new_n1155), .A4(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1157), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1140), .B1(new_n1174), .B2(new_n778), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1087), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1171), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1169), .A2(new_n912), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1178), .A2(new_n1152), .B1(new_n1144), .B2(new_n942), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1172), .B1(new_n1179), .B2(new_n1150), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1177), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n453), .A2(new_n1159), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n948), .A2(new_n1182), .A3(new_n679), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n771), .A2(G330), .A3(new_n882), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1184), .A2(new_n1143), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n1185), .A2(new_n1160), .B1(new_n892), .B2(new_n913), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n912), .B1(new_n1159), .B2(new_n882), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1169), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1150), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1183), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1176), .B1(new_n1181), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1190), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1174), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1175), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(G378));
  INV_X1    g0995(.A(KEYINPUT120), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n927), .A2(new_n937), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n953), .A2(new_n882), .A3(new_n912), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT40), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(G330), .B1(new_n954), .B2(new_n956), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1196), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT40), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n935), .B2(new_n936), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1158), .B1(new_n1198), .B2(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1204), .B(KEYINPUT120), .C1(new_n955), .C2(KEYINPUT40), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n355), .A2(new_n359), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n345), .A2(new_n711), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1206), .B(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1208), .B(new_n1209), .Z(new_n1210));
  NAND3_X1  g1010(.A1(new_n1201), .A2(new_n1205), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1210), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1212), .B(new_n1196), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1211), .A2(new_n947), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n947), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n779), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n846), .B1(new_n201), .B2(new_n847), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT118), .Z(new_n1219));
  NOR2_X1   g1019(.A1(G33), .A2(G41), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT115), .Z(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n201), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n277), .B2(new_n326), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n803), .A2(new_n519), .B1(new_n806), .B2(new_n202), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G116), .B2(new_n823), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G41), .B(new_n328), .C1(G97), .C2(new_n813), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(G283), .A2(new_n821), .B1(new_n839), .B2(new_n507), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1054), .B1(G68), .B2(new_n811), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT58), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1223), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  XNOR2_X1  g1031(.A(KEYINPUT117), .B(G124), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1221), .B1(new_n821), .B2(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n839), .A2(G137), .B1(G132), .B2(new_n813), .ZN(new_n1234));
  INV_X1    g1034(.A(G128), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1234), .B1(new_n1235), .B2(new_n803), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n811), .A2(G150), .B1(new_n823), .B2(G125), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT116), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1130), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1236), .B(new_n1238), .C1(new_n825), .C2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT59), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1233), .B1(new_n832), .B2(new_n806), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1231), .B1(new_n1230), .B2(new_n1229), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1219), .B1(new_n1244), .B2(new_n795), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1245), .B1(new_n1212), .B2(new_n783), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT119), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1217), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n947), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1211), .A2(new_n947), .A3(new_n1213), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(KEYINPUT57), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1186), .A2(new_n1189), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1183), .B1(new_n1181), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT121), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT121), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1190), .A2(new_n1157), .A3(new_n1171), .A4(new_n1173), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1183), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1216), .A2(new_n1258), .A3(KEYINPUT57), .A4(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1257), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1253), .A3(new_n1252), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT57), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1176), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1249), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(G375));
  NAND2_X1  g1068(.A1(new_n1143), .A2(new_n782), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n780), .B1(new_n848), .B2(G68), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n839), .A2(G107), .B1(G116), .B2(new_n813), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1271), .B(KEYINPUT123), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n328), .B(new_n989), .C1(G303), .C2(new_n821), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1055), .B1(G283), .B2(new_n802), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(G294), .A2(new_n823), .B1(new_n825), .B2(G97), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT124), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n803), .A2(new_n866), .B1(new_n201), .B2(new_n810), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(G159), .B2(new_n825), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n820), .A2(new_n1235), .B1(new_n817), .B2(new_n1057), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n326), .B(new_n1281), .C1(new_n813), .C2(new_n1239), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(G132), .A2(new_n823), .B1(new_n982), .B2(G58), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1280), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1278), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1270), .B1(new_n1286), .B2(new_n795), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1255), .A2(new_n779), .B1(new_n1269), .B2(new_n1287), .ZN(new_n1288));
  XOR2_X1   g1088(.A(new_n1029), .B(KEYINPUT122), .Z(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1192), .A2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1255), .A2(new_n1260), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1288), .B1(new_n1291), .B2(new_n1292), .ZN(G381));
  OR2_X1    g1093(.A1(G393), .A2(G396), .ZN(new_n1294));
  OR4_X1    g1094(.A1(G384), .A2(G381), .A3(G390), .A4(new_n1294), .ZN(new_n1295));
  OR4_X1    g1095(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1295), .ZN(G407));
  INV_X1    g1096(.A(G213), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(G343), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1267), .A2(new_n1194), .A3(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(G407), .A2(G213), .A3(new_n1299), .ZN(G409));
  NAND2_X1  g1100(.A1(G387), .A2(KEYINPUT127), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT106), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1302));
  AOI211_X1 g1102(.A(new_n1032), .B(new_n1029), .C1(new_n1027), .C2(new_n773), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n778), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1051), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT127), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1305), .A2(new_n1306), .A3(new_n995), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(G393), .A2(G396), .ZN(new_n1308));
  AND3_X1   g1108(.A1(G390), .A2(new_n1294), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G390), .B1(new_n1294), .B2(new_n1308), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1301), .A2(new_n1307), .A3(new_n1311), .ZN(new_n1312));
  OR2_X1    g1112(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1306), .B1(new_n1305), .B2(new_n995), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n995), .ZN(new_n1315));
  AOI211_X1 g1115(.A(KEYINPUT127), .B(new_n1315), .C1(new_n1304), .C2(new_n1051), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1313), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1312), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT61), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1214), .A2(new_n1215), .A3(new_n1265), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1258), .B1(new_n1320), .B2(new_n1261), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1254), .A2(new_n1256), .A3(KEYINPUT121), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1266), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1249), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1323), .A2(G378), .A3(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1261), .A2(new_n1253), .A3(new_n1252), .A4(new_n1290), .ZN(new_n1326));
  AND2_X1   g1126(.A1(new_n1326), .A2(new_n1246), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1216), .A2(KEYINPUT125), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT125), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1329), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1328), .A2(new_n779), .A3(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1327), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1332), .A2(new_n1194), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1298), .B1(new_n1325), .B2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1292), .A2(KEYINPUT60), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT60), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1336), .B1(new_n1255), .B2(new_n1260), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1335), .A2(new_n1087), .A3(new_n1192), .A4(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1338), .A2(G384), .A3(new_n1288), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(G384), .B1(new_n1338), .B2(new_n1288), .ZN(new_n1341));
  OAI211_X1 g1141(.A(G2897), .B(new_n1298), .C1(new_n1340), .C2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1341), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1298), .A2(G2897), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(new_n1339), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1342), .A2(new_n1345), .ZN(new_n1346));
  OAI211_X1 g1146(.A(new_n1318), .B(new_n1319), .C1(new_n1334), .C2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT126), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1350), .ZN(new_n1351));
  AOI211_X1 g1151(.A(new_n1298), .B(new_n1351), .C1(new_n1325), .C2(new_n1333), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1349), .B1(new_n1352), .B2(KEYINPUT63), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1352), .A2(KEYINPUT63), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1298), .ZN(new_n1355));
  AOI211_X1 g1155(.A(new_n1194), .B(new_n1249), .C1(new_n1263), .C2(new_n1266), .ZN(new_n1356));
  AOI21_X1  g1156(.A(G378), .B1(new_n1327), .B2(new_n1331), .ZN(new_n1357));
  OAI211_X1 g1157(.A(new_n1355), .B(new_n1350), .C1(new_n1356), .C2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT63), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1358), .A2(KEYINPUT126), .A3(new_n1359), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1348), .A2(new_n1353), .A3(new_n1354), .A4(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1358), .A2(KEYINPUT62), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1325), .A2(new_n1333), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT62), .ZN(new_n1364));
  NAND4_X1  g1164(.A1(new_n1363), .A2(new_n1364), .A3(new_n1355), .A4(new_n1350), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1346), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1357), .B1(new_n1267), .B2(G378), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1366), .B1(new_n1367), .B2(new_n1298), .ZN(new_n1368));
  NAND4_X1  g1168(.A1(new_n1362), .A2(new_n1319), .A3(new_n1365), .A4(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1318), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1369), .A2(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1361), .A2(new_n1371), .ZN(G405));
  NOR2_X1   g1172(.A1(new_n1267), .A2(G378), .ZN(new_n1373));
  OR3_X1    g1173(.A1(new_n1373), .A2(new_n1356), .A3(new_n1350), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1350), .B1(new_n1373), .B2(new_n1356), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1374), .A2(new_n1375), .ZN(new_n1376));
  XNOR2_X1  g1176(.A(new_n1376), .B(new_n1370), .ZN(G402));
endmodule


