//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT22), .ZN(new_n192));
  INV_X1    g006(.A(G137), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G110), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n206), .B1(new_n210), .B2(new_n204), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(G146), .B(new_n206), .C1(new_n210), .C2(new_n204), .ZN(new_n214));
  XNOR2_X1  g028(.A(G119), .B(G128), .ZN(new_n215));
  AND2_X1   g029(.A1(KEYINPUT24), .A2(G110), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT24), .A2(G110), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT76), .B1(new_n218), .B2(new_n215), .ZN(new_n220));
  INV_X1    g034(.A(G110), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n198), .A2(new_n201), .A3(new_n221), .A4(new_n200), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n200), .A2(new_n196), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT24), .B(G110), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT76), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n220), .A2(new_n222), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT77), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n210), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G125), .B(G140), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT77), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n231), .A3(new_n212), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n214), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT78), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT78), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n227), .A2(new_n235), .A3(new_n214), .A4(new_n232), .ZN(new_n236));
  AOI221_X4 g050(.A(new_n194), .B1(new_n203), .B2(new_n219), .C1(new_n234), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n194), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n236), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n219), .A2(new_n203), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT25), .B1(new_n242), .B2(new_n188), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n232), .A2(new_n214), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n235), .B1(new_n244), .B2(new_n227), .ZN(new_n245));
  INV_X1    g059(.A(new_n236), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n240), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n194), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n239), .A2(new_n240), .A3(new_n238), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n248), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n189), .B1(new_n243), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n242), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n189), .A2(G902), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(KEYINPUT79), .B1(new_n252), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n189), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n248), .A2(new_n188), .A3(new_n249), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT25), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n259), .B1(new_n262), .B2(new_n250), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT79), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n263), .A2(new_n264), .A3(new_n256), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT11), .ZN(new_n267));
  INV_X1    g081(.A(G134), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(G137), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(G137), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n193), .A2(KEYINPUT11), .A3(G134), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G131), .ZN(new_n273));
  INV_X1    g087(.A(G131), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n269), .A2(new_n271), .A3(new_n274), .A4(new_n270), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n212), .A2(G143), .ZN(new_n277));
  INV_X1    g091(.A(G143), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G146), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n281));
  NAND2_X1  g095(.A1(KEYINPUT0), .A2(G128), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR3_X1   g097(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(G143), .B(G146), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n282), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n276), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(KEYINPUT2), .A2(G113), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT68), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n294));
  INV_X1    g108(.A(G113), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n292), .A2(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(G116), .B(G119), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n292), .A2(new_n293), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n294), .A2(new_n295), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n299), .A2(new_n300), .A3(new_n297), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n303));
  AND4_X1   g117(.A1(new_n303), .A2(new_n277), .A3(new_n279), .A4(G128), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT1), .B1(new_n278), .B2(G146), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT67), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT67), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n277), .A2(new_n307), .A3(KEYINPUT1), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n306), .A2(G128), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n304), .B1(new_n309), .B2(new_n280), .ZN(new_n310));
  XNOR2_X1  g124(.A(G134), .B(G137), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT66), .B1(new_n311), .B2(new_n274), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT66), .ZN(new_n313));
  INV_X1    g127(.A(new_n270), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n268), .A2(G137), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n313), .B(G131), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n312), .A2(new_n316), .A3(new_n275), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n289), .B(new_n302), .C1(new_n310), .C2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT26), .ZN(new_n319));
  AND2_X1   g133(.A1(KEYINPUT69), .A2(G237), .ZN(new_n320));
  NOR2_X1   g134(.A1(KEYINPUT69), .A2(G237), .ZN(new_n321));
  OAI211_X1 g135(.A(G210), .B(new_n190), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT27), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT69), .B(G237), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G210), .A4(new_n190), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n319), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n326), .A3(new_n319), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(G101), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(G101), .ZN(new_n331));
  INV_X1    g145(.A(new_n329), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(new_n327), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n318), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT70), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n318), .A2(new_n333), .A3(new_n330), .A4(KEYINPUT70), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n298), .A2(new_n301), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n273), .A2(new_n275), .B1(new_n285), .B2(new_n287), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n309), .A2(new_n280), .ZN(new_n341));
  INV_X1    g155(.A(new_n304), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n317), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT64), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT30), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n289), .B1(new_n310), .B2(new_n317), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT30), .B1(new_n349), .B2(KEYINPUT64), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n339), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n338), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT31), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT71), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT28), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n354), .B1(new_n318), .B2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n310), .A2(new_n317), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n339), .B1(new_n357), .B2(new_n340), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n358), .A2(new_n318), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n359), .B2(new_n355), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n333), .A2(new_n330), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n358), .A2(new_n318), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n354), .A3(KEYINPUT28), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT31), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n338), .A2(new_n351), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n353), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(G472), .A2(G902), .ZN(new_n368));
  AND3_X1   g182(.A1(new_n367), .A2(KEYINPUT32), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT73), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n358), .A2(new_n370), .A3(new_n318), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n349), .A2(KEYINPUT73), .A3(new_n339), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(KEYINPUT28), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT74), .ZN(new_n374));
  INV_X1    g188(.A(new_n318), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n374), .B1(new_n375), .B2(KEYINPUT28), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT29), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n361), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n371), .A2(new_n374), .A3(KEYINPUT28), .A4(new_n372), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n188), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT75), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n347), .B1(new_n345), .B2(new_n346), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n349), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n375), .B1(new_n387), .B2(new_n339), .ZN(new_n388));
  INV_X1    g202(.A(new_n361), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n378), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n361), .B1(new_n360), .B2(new_n363), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n381), .A2(KEYINPUT75), .A3(new_n188), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n384), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n369), .B1(new_n394), .B2(G472), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT32), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT72), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n367), .A2(new_n397), .A3(new_n368), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n397), .B1(new_n367), .B2(new_n368), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n266), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G475), .ZN(new_n402));
  OAI211_X1 g216(.A(G214), .B(new_n190), .C1(new_n320), .C2(new_n321), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n278), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n324), .A2(G143), .A3(G214), .A4(new_n190), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G131), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT89), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT89), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n410), .A3(G131), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n404), .A2(new_n405), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n274), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n408), .A2(new_n409), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n213), .A2(new_n214), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n410), .B1(new_n406), .B2(G131), .ZN(new_n416));
  AOI211_X1 g230(.A(KEYINPUT89), .B(new_n274), .C1(new_n404), .C2(new_n405), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT17), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n412), .B1(new_n420), .B2(new_n274), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n232), .B1(new_n212), .B2(new_n230), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n406), .A2(KEYINPUT18), .A3(G131), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G113), .B(G122), .ZN(new_n426));
  INV_X1    g240(.A(G104), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n419), .A2(new_n428), .A3(new_n424), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n402), .B1(new_n432), .B2(new_n188), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT90), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n229), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT19), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n228), .B1(new_n436), .B2(KEYINPUT90), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n435), .A2(new_n436), .B1(new_n230), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n214), .B1(new_n438), .B2(G146), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n416), .A2(new_n417), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n439), .B1(new_n440), .B2(new_n413), .ZN(new_n441));
  INV_X1    g255(.A(new_n424), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n429), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n431), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(G475), .A2(G902), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n444), .A2(KEYINPUT20), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT20), .B1(new_n444), .B2(new_n445), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n433), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G952), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(G953), .ZN(new_n450));
  NAND2_X1  g264(.A1(G234), .A2(G237), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT21), .B(G898), .Z(new_n453));
  NAND3_X1  g267(.A1(new_n451), .A2(G902), .A3(G953), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G116), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(G122), .ZN(new_n457));
  INV_X1    g271(.A(G122), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G116), .ZN(new_n459));
  OAI21_X1  g273(.A(G107), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(G116), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n456), .A2(G122), .ZN(new_n462));
  INV_X1    g276(.A(G107), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT13), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n195), .B2(G143), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n195), .A2(G143), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n278), .A2(KEYINPUT13), .A3(G128), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G134), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n278), .A2(G128), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n468), .A3(new_n268), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n465), .A2(new_n471), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT14), .B1(new_n456), .B2(G122), .ZN(new_n475));
  OAI211_X1 g289(.A(G107), .B(new_n475), .C1(new_n457), .C2(new_n459), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n461), .B(new_n462), .C1(KEYINPUT14), .C2(new_n463), .ZN(new_n477));
  INV_X1    g291(.A(new_n473), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n268), .B1(new_n472), .B2(new_n468), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n476), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(KEYINPUT9), .B(G234), .Z(new_n481));
  INV_X1    g295(.A(KEYINPUT91), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n481), .A2(new_n482), .A3(G217), .A4(new_n190), .ZN(new_n483));
  OR2_X1    g297(.A1(KEYINPUT9), .A2(G234), .ZN(new_n484));
  NAND2_X1  g298(.A1(KEYINPUT9), .A2(G234), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n484), .A2(G217), .A3(new_n190), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT91), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n474), .A2(new_n480), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n488), .B1(new_n474), .B2(new_n480), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n188), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G478), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n492), .B(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n448), .A2(new_n455), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G469), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT3), .B1(new_n427), .B2(G107), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT3), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n463), .A3(G104), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n427), .A2(G107), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n498), .A2(new_n500), .A3(new_n331), .A4(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n463), .A2(G104), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n427), .A2(G107), .ZN(new_n504));
  OAI21_X1  g318(.A(G101), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT83), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n502), .B2(new_n505), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n343), .A2(new_n508), .A3(KEYINPUT10), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(KEYINPUT81), .A3(G101), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n512), .A2(KEYINPUT81), .A3(KEYINPUT4), .A4(G101), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n288), .ZN(new_n518));
  INV_X1    g332(.A(new_n276), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT82), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n195), .B1(new_n305), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n277), .A2(KEYINPUT82), .A3(KEYINPUT1), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n286), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n506), .B1(new_n523), .B2(new_n304), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT10), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n511), .A2(new_n518), .A3(new_n519), .A4(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G110), .B(G140), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n190), .A2(G227), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n524), .B1(new_n343), .B2(new_n506), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT12), .B1(new_n276), .B2(KEYINPUT84), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n276), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n502), .A2(new_n505), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n341), .A2(new_n342), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n521), .A2(new_n522), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n280), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n539), .B2(new_n342), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n276), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(new_n533), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n531), .B1(new_n535), .B2(new_n542), .ZN(new_n543));
  AOI22_X1  g357(.A1(new_n517), .A2(new_n288), .B1(new_n524), .B2(new_n525), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n511), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n276), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n530), .B1(new_n546), .B2(new_n527), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n497), .B(new_n188), .C1(new_n543), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(G469), .A2(G902), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n532), .A2(new_n276), .A3(new_n534), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n534), .B1(new_n532), .B2(new_n276), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n527), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n530), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n546), .A2(new_n527), .A3(new_n530), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(G469), .A3(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n548), .A2(new_n549), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n481), .A2(new_n188), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G221), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n559), .B(KEYINPUT80), .Z(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  XOR2_X1   g376(.A(G110), .B(G122), .Z(new_n563));
  AOI21_X1  g377(.A(new_n302), .B1(new_n515), .B2(new_n516), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n536), .A2(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n199), .A2(G116), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n456), .A2(G119), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT5), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n568), .B(G113), .C1(KEYINPUT5), .C2(new_n566), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n296), .A2(new_n297), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n565), .A2(new_n571), .A3(new_n509), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n563), .B1(new_n564), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n517), .A2(new_n339), .ZN(new_n574));
  INV_X1    g388(.A(new_n571), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(new_n510), .A3(new_n508), .ZN(new_n576));
  INV_X1    g390(.A(new_n563), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n573), .A2(KEYINPUT6), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT6), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n580), .B(new_n563), .C1(new_n564), .C2(new_n572), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n310), .A2(new_n208), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n285), .A2(G125), .A3(new_n287), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n190), .A2(G224), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n585), .B(KEYINPUT85), .Z(new_n586));
  XNOR2_X1  g400(.A(new_n584), .B(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n579), .A2(new_n581), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT87), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n582), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n310), .A2(KEYINPUT87), .A3(new_n208), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n583), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n585), .A2(KEYINPUT7), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n536), .A2(KEYINPUT86), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n575), .B(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n563), .B(KEYINPUT8), .Z(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n585), .A2(KEYINPUT88), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n582), .A2(new_n583), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT7), .B1(new_n585), .B2(KEYINPUT88), .ZN(new_n601));
  OR2_X1    g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n594), .A2(new_n598), .A3(new_n578), .A4(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n588), .A2(new_n188), .A3(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(G210), .B1(G237), .B2(G902), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n588), .A2(new_n603), .A3(new_n188), .A4(new_n605), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(G214), .B1(G237), .B2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n496), .A2(new_n562), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n401), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  NAND2_X1  g428(.A1(new_n367), .A2(new_n188), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n615), .A2(G472), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n398), .B2(new_n399), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n617), .A2(new_n266), .A3(new_n562), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT92), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT94), .B1(new_n489), .B2(new_n490), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n474), .A2(new_n488), .A3(new_n480), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT94), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n620), .A2(KEYINPUT33), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT95), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n491), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT95), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n620), .A2(new_n628), .A3(KEYINPUT33), .A4(new_n623), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n625), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n630), .A2(KEYINPUT96), .A3(G478), .A4(new_n188), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n625), .A2(G478), .A3(new_n627), .A4(new_n629), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(G902), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT97), .B(G478), .Z(new_n636));
  NAND2_X1  g450(.A1(new_n492), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n431), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n428), .B1(new_n419), .B2(new_n424), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n188), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(G475), .ZN(new_n642));
  INV_X1    g456(.A(new_n447), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n444), .A2(KEYINPUT20), .A3(new_n445), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n638), .A2(KEYINPUT98), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n631), .A2(new_n634), .B1(new_n492), .B2(new_n636), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n647), .B1(new_n648), .B2(new_n448), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT93), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n607), .A2(new_n650), .A3(new_n608), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n604), .A2(KEYINPUT93), .A3(new_n606), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n651), .A2(new_n455), .A3(new_n610), .A4(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  AND3_X1   g468(.A1(new_n646), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n619), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT34), .B(G104), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  INV_X1    g473(.A(new_n495), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n448), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n619), .A2(new_n653), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT35), .B(G107), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NOR2_X1   g478(.A1(new_n194), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n247), .B(new_n665), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n263), .B1(new_n254), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n668), .B(new_n616), .C1(new_n399), .C2(new_n398), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n612), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(KEYINPUT37), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n221), .ZN(G12));
  NAND2_X1  g487(.A1(new_n395), .A2(new_n400), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n452), .B1(G900), .B2(new_n454), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n448), .A2(new_n660), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n651), .A2(new_n610), .A3(new_n652), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n562), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n674), .A2(new_n676), .A3(new_n668), .A4(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT99), .B(G128), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G30));
  INV_X1    g495(.A(KEYINPUT101), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n367), .A2(KEYINPUT32), .A3(new_n368), .ZN(new_n683));
  INV_X1    g497(.A(new_n352), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n371), .A2(new_n361), .A3(new_n372), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n188), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(G472), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n400), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n688), .A2(new_n667), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n557), .A2(new_n561), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n675), .B(KEYINPUT39), .Z(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n693), .A2(KEYINPUT100), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(KEYINPUT100), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT40), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(KEYINPUT40), .B1(new_n694), .B2(new_n695), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n689), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n609), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n701), .A2(KEYINPUT38), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n448), .A2(new_n495), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(KEYINPUT38), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n702), .A2(new_n703), .A3(new_n610), .A4(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n682), .B1(new_n700), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n696), .B(new_n697), .ZN(new_n707));
  INV_X1    g521(.A(new_n705), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n707), .A2(KEYINPUT101), .A3(new_n708), .A4(new_n689), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n278), .ZN(G45));
  NAND3_X1  g525(.A1(new_n638), .A2(new_n645), .A3(new_n675), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n674), .A2(new_n668), .A3(new_n678), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G146), .ZN(G48));
  INV_X1    g529(.A(new_n547), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n542), .A2(new_n535), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n527), .A3(new_n530), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n497), .B1(new_n719), .B2(new_n188), .ZN(new_n720));
  INV_X1    g534(.A(new_n548), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n720), .A2(new_n721), .A3(new_n560), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n655), .A2(new_n401), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  NOR2_X1   g539(.A1(new_n661), .A2(new_n653), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n401), .A2(new_n726), .A3(new_n722), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT102), .B(G116), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G18));
  AOI21_X1  g543(.A(new_n667), .B1(new_n395), .B2(new_n400), .ZN(new_n730));
  INV_X1    g544(.A(new_n496), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n720), .A2(new_n721), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n561), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n677), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n730), .A2(new_n731), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n338), .A2(new_n351), .A3(new_n365), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n365), .B1(new_n338), .B2(new_n351), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n377), .A2(new_n380), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n361), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n368), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n263), .A2(new_n256), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n616), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(KEYINPUT103), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT103), .ZN(new_n748));
  INV_X1    g562(.A(G472), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n749), .B1(new_n367), .B2(new_n188), .ZN(new_n750));
  INV_X1    g564(.A(new_n368), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n751), .B1(new_n740), .B2(new_n742), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n748), .B1(new_n753), .B2(new_n745), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n722), .B1(new_n747), .B2(new_n754), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n448), .A2(KEYINPUT104), .A3(new_n495), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n757), .B1(new_n645), .B2(new_n660), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n756), .A2(new_n758), .A3(new_n653), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n737), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n746), .A2(KEYINPUT103), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n753), .A2(new_n748), .A3(new_n745), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n733), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(KEYINPUT105), .A3(new_n759), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  NOR3_X1   g581(.A1(new_n667), .A2(new_n750), .A3(new_n752), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n734), .A2(new_n713), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G125), .ZN(G27));
  OR2_X1    g584(.A1(new_n258), .A2(new_n265), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n381), .A2(KEYINPUT75), .A3(new_n188), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT75), .B1(new_n381), .B2(new_n188), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n390), .A2(new_n391), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n683), .B1(new_n775), .B2(new_n749), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n367), .A2(new_n368), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT72), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n367), .A2(new_n397), .A3(new_n368), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT32), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n771), .B1(new_n776), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n607), .A2(new_n610), .A3(new_n608), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT106), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n607), .A2(KEYINPUT106), .A3(new_n610), .A4(new_n608), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n648), .A2(new_n448), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n690), .A3(new_n787), .A4(new_n675), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT107), .B1(new_n781), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT42), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n690), .A2(new_n784), .A3(new_n785), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n712), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT107), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n401), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n777), .A2(new_n396), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n683), .B(new_n796), .C1(new_n775), .C2(new_n749), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n797), .A2(KEYINPUT108), .A3(new_n745), .ZN(new_n798));
  AOI21_X1  g612(.A(KEYINPUT108), .B1(new_n797), .B2(new_n745), .ZN(new_n799));
  OAI211_X1 g613(.A(KEYINPUT42), .B(new_n792), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G131), .ZN(G33));
  INV_X1    g616(.A(new_n791), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n401), .A2(new_n676), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G134), .ZN(G36));
  NAND2_X1  g619(.A1(new_n784), .A2(new_n785), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n638), .B(new_n448), .C1(KEYINPUT109), .C2(KEYINPUT43), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT109), .A4(new_n644), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT43), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n808), .B(new_n809), .C1(new_n648), .C2(new_n645), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT110), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n667), .ZN(new_n814));
  INV_X1    g628(.A(new_n617), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n815), .B1(new_n811), .B2(new_n812), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n806), .B1(new_n817), .B2(KEYINPUT44), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT45), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n530), .B1(new_n717), .B2(new_n527), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n519), .B1(new_n544), .B2(new_n511), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n531), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n819), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n554), .A2(KEYINPUT45), .A3(new_n555), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n823), .A2(new_n824), .A3(G469), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n549), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT46), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n825), .A2(KEYINPUT46), .A3(new_n549), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n548), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n561), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n691), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n814), .A2(new_n816), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT44), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n818), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(G137), .ZN(G39));
  NOR2_X1   g652(.A1(new_n674), .A2(new_n712), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n266), .A3(new_n786), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n840), .A2(KEYINPUT111), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n825), .A2(KEYINPUT46), .A3(new_n549), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT46), .B1(new_n825), .B2(new_n549), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n842), .A2(new_n843), .A3(new_n721), .ZN(new_n844));
  OAI21_X1  g658(.A(KEYINPUT47), .B1(new_n844), .B2(new_n560), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT47), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n830), .A2(new_n846), .A3(new_n561), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n840), .A2(KEYINPUT111), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n841), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(G140), .ZN(G42));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  INV_X1    g668(.A(new_n804), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n795), .B2(new_n800), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n612), .B1(new_n401), .B2(new_n670), .ZN(new_n857));
  INV_X1    g671(.A(new_n611), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n661), .B1(new_n448), .B2(new_n648), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n618), .A2(new_n455), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n761), .B2(new_n765), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n768), .A2(new_n787), .A3(new_n675), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT112), .B1(new_n863), .B2(new_n791), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT112), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n803), .A2(new_n713), .A3(new_n865), .A4(new_n768), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n448), .A2(new_n495), .A3(new_n675), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n667), .B(new_n867), .C1(new_n395), .C2(new_n400), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n864), .A2(new_n866), .B1(new_n868), .B2(new_n803), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n723), .A2(new_n727), .A3(new_n735), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n856), .A2(new_n862), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n756), .A2(new_n758), .A3(new_n677), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n667), .A3(new_n675), .A4(new_n688), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n562), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n679), .A2(new_n714), .A3(new_n769), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT52), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n689), .A2(new_n690), .A3(new_n675), .A4(new_n872), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n730), .B(new_n678), .C1(new_n676), .C2(new_n713), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n769), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n854), .B1(new_n871), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT113), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n876), .A2(new_n880), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n857), .A2(new_n860), .ZN(new_n885));
  AND4_X1   g699(.A1(new_n766), .A2(new_n870), .A3(new_n869), .A4(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT53), .A4(new_n856), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n882), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n871), .A2(new_n881), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n889), .A2(KEYINPUT113), .A3(KEYINPUT53), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n888), .A2(KEYINPUT54), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n882), .A2(new_n892), .A3(new_n887), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n786), .A2(new_n451), .A3(new_n450), .A4(new_n722), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n895), .A2(new_n688), .A3(new_n266), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(KEYINPUT114), .A3(new_n448), .A4(new_n648), .ZN(new_n897));
  AND4_X1   g711(.A1(new_n771), .A2(new_n400), .A3(new_n683), .A4(new_n687), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n733), .A2(new_n806), .A3(new_n452), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(new_n448), .A3(new_n648), .A4(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT114), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n452), .B1(new_n807), .B2(new_n810), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n610), .B1(new_n702), .B2(new_n704), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n764), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT50), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n764), .A2(KEYINPUT50), .A3(new_n904), .A4(new_n905), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n732), .A2(new_n560), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n830), .A2(new_n846), .A3(new_n561), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n846), .B1(new_n830), .B2(new_n561), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n762), .A2(new_n763), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n904), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n914), .A2(new_n916), .A3(new_n786), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n811), .A2(new_n895), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n768), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n903), .A2(new_n910), .A3(new_n917), .A4(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT51), .B1(new_n917), .B2(KEYINPUT115), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n806), .B1(new_n848), .B2(new_n911), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n902), .A2(new_n897), .B1(new_n924), .B2(new_n916), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n925), .A2(new_n921), .A3(new_n919), .A4(new_n910), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  OR4_X1    g741(.A1(new_n452), .A2(new_n755), .A3(new_n677), .A4(new_n811), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT48), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n798), .A2(new_n799), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(new_n918), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n918), .B(new_n929), .C1(new_n798), .C2(new_n799), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n450), .B(new_n928), .C1(new_n931), .C2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n896), .A2(new_n649), .A3(new_n646), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n927), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT116), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n934), .B1(new_n923), .B2(new_n926), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(KEYINPUT116), .A3(new_n936), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n853), .B1(new_n894), .B2(new_n942), .ZN(new_n943));
  AND4_X1   g757(.A1(KEYINPUT116), .A2(new_n927), .A3(new_n935), .A4(new_n936), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT116), .B1(new_n940), .B2(new_n936), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n946), .A2(KEYINPUT117), .A3(new_n891), .A4(new_n893), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n449), .A2(new_n190), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n943), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n702), .A2(new_n704), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n648), .A2(new_n645), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n950), .A2(new_n561), .A3(new_n610), .A4(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n732), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(KEYINPUT49), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT49), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n745), .B1(new_n732), .B2(new_n955), .ZN(new_n956));
  OR4_X1    g770(.A1(new_n688), .A2(new_n952), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n949), .A2(new_n957), .ZN(G75));
  NOR2_X1   g772(.A1(new_n190), .A2(G952), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT120), .Z(new_n960));
  AOI21_X1  g774(.A(new_n188), .B1(new_n882), .B2(new_n887), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(G210), .ZN(new_n962));
  NAND2_X1  g776(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n962), .A2(KEYINPUT119), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n579), .A2(new_n581), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(new_n587), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT55), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT119), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT56), .B1(new_n970), .B2(KEYINPUT118), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n962), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n960), .B1(new_n968), .B2(new_n972), .ZN(G51));
  XNOR2_X1  g787(.A(new_n719), .B(KEYINPUT121), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n882), .A2(new_n887), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(KEYINPUT54), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n893), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n549), .B(KEYINPUT57), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n974), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n825), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n961), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n959), .B1(new_n980), .B2(new_n982), .ZN(G54));
  INV_X1    g797(.A(new_n959), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n961), .A2(KEYINPUT58), .A3(G475), .ZN(new_n985));
  INV_X1    g799(.A(new_n444), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT122), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n985), .A2(new_n988), .A3(new_n986), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n988), .B1(new_n985), .B2(new_n986), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n984), .B(new_n987), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(G60));
  INV_X1    g806(.A(KEYINPUT123), .ZN(new_n993));
  NAND2_X1  g807(.A1(G478), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT59), .Z(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n630), .B1(new_n894), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n630), .A2(new_n996), .ZN(new_n998));
  INV_X1    g812(.A(new_n893), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n892), .B1(new_n882), .B2(new_n887), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n960), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n993), .B1(new_n997), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n960), .B1(new_n977), .B2(new_n998), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n995), .B1(new_n891), .B2(new_n893), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1005), .B(KEYINPUT123), .C1(new_n630), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1004), .A2(new_n1007), .ZN(G63));
  INV_X1    g822(.A(KEYINPUT61), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G217), .A2(G902), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1010), .B(KEYINPUT60), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1011), .B1(new_n882), .B2(new_n887), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1002), .B1(new_n1012), .B2(new_n242), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT124), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1009), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT125), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1011), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n975), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n960), .B1(new_n1018), .B2(new_n253), .ZN(new_n1019));
  INV_X1    g833(.A(new_n666), .ZN(new_n1020));
  AOI211_X1 g834(.A(new_n1020), .B(new_n1011), .C1(new_n882), .C2(new_n887), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1016), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n1013), .A2(KEYINPUT125), .A3(new_n1021), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1015), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(KEYINPUT61), .B1(new_n1019), .B2(KEYINPUT124), .ZN(new_n1026));
  OAI21_X1  g840(.A(KEYINPUT125), .B1(new_n1013), .B2(new_n1021), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1019), .A2(new_n1016), .A3(new_n1022), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1025), .A2(new_n1029), .ZN(G66));
  AOI21_X1  g844(.A(new_n190), .B1(new_n453), .B2(G224), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n862), .A2(new_n870), .ZN(new_n1032));
  INV_X1    g846(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1031), .B1(new_n1033), .B2(new_n190), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n965), .B1(G898), .B2(new_n190), .ZN(new_n1035));
  XOR2_X1   g849(.A(new_n1034), .B(new_n1035), .Z(G69));
  XOR2_X1   g850(.A(new_n387), .B(new_n438), .Z(new_n1037));
  NAND2_X1  g851(.A1(G900), .A2(G953), .ZN(new_n1038));
  AND3_X1   g852(.A1(new_n841), .A2(new_n849), .A3(new_n850), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1039), .B1(new_n818), .B2(new_n836), .ZN(new_n1040));
  INV_X1    g854(.A(new_n875), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n930), .A2(new_n832), .A3(new_n872), .ZN(new_n1042));
  XNOR2_X1  g856(.A(new_n1042), .B(KEYINPUT127), .ZN(new_n1043));
  NAND4_X1  g857(.A1(new_n1040), .A2(new_n856), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1044));
  OAI211_X1 g858(.A(new_n1037), .B(new_n1038), .C1(new_n1044), .C2(G953), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n832), .B1(new_n817), .B2(KEYINPUT44), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n786), .B1(new_n834), .B2(new_n835), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n851), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n706), .A2(new_n709), .A3(new_n1041), .ZN(new_n1049));
  INV_X1    g863(.A(KEYINPUT62), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g865(.A1(new_n706), .A2(new_n709), .A3(KEYINPUT62), .A4(new_n1041), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1048), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g867(.A1(new_n696), .A2(new_n806), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n1054), .A2(new_n401), .A3(new_n859), .ZN(new_n1055));
  AOI21_X1  g869(.A(G953), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1045), .B1(new_n1056), .B2(new_n1037), .ZN(new_n1057));
  AOI21_X1  g871(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n1058), .B1(new_n1045), .B2(KEYINPUT126), .ZN(new_n1059));
  AND2_X1   g873(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g874(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1061));
  NOR2_X1   g875(.A1(new_n1060), .A2(new_n1061), .ZN(G72));
  NAND3_X1  g876(.A1(new_n1053), .A2(new_n1032), .A3(new_n1055), .ZN(new_n1063));
  NAND2_X1  g877(.A1(G472), .A2(G902), .ZN(new_n1064));
  XOR2_X1   g878(.A(new_n1064), .B(KEYINPUT63), .Z(new_n1065));
  AOI211_X1 g879(.A(new_n361), .B(new_n388), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g880(.A(new_n1065), .B1(new_n1044), .B2(new_n1033), .ZN(new_n1067));
  AND3_X1   g881(.A1(new_n1067), .A2(new_n361), .A3(new_n388), .ZN(new_n1068));
  OAI21_X1  g882(.A(new_n352), .B1(new_n389), .B2(new_n388), .ZN(new_n1069));
  AND4_X1   g883(.A1(new_n890), .A2(new_n888), .A3(new_n1065), .A4(new_n1069), .ZN(new_n1070));
  NOR4_X1   g884(.A1(new_n1066), .A2(new_n1068), .A3(new_n959), .A4(new_n1070), .ZN(G57));
endmodule


