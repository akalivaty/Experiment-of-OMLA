//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  OR3_X1    g0009(.A1(new_n209), .A2(KEYINPUT64), .A3(G13), .ZN(new_n210));
  OAI21_X1  g0010(.A(KEYINPUT64), .B1(new_n209), .B2(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n202), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G107), .ZN(new_n223));
  INV_X1    g0023(.A(G264), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT1), .Z(new_n227));
  NAND2_X1  g0027(.A1(new_n203), .A2(G50), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT66), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT65), .B(G20), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n214), .A2(new_n227), .A3(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT67), .Z(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n202), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n246), .B(new_n252), .Z(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n231), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n257), .A3(new_n231), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G150), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT8), .A2(G58), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT69), .B(G58), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT8), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n230), .A2(G33), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n261), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT70), .ZN(new_n269));
  AND2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(new_n268), .B2(new_n269), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n259), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n207), .A2(G1), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(new_n247), .ZN(new_n275));
  INV_X1    g0075(.A(G13), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G1), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G20), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n256), .A2(new_n275), .A3(new_n258), .A4(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n279), .B1(G50), .B2(new_n278), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT71), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n273), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  OAI211_X1 g0085(.A(G1), .B(G13), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  AOI21_X1  g0087(.A(G1), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(G274), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G226), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n289), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT3), .B(G33), .ZN(new_n294));
  INV_X1    g0094(.A(G1698), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(G222), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G223), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n296), .B1(new_n221), .B2(new_n294), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n293), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n303), .A2(KEYINPUT72), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n303), .A2(KEYINPUT72), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n283), .B1(G169), .B2(new_n301), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n301), .A2(G190), .ZN(new_n308));
  XNOR2_X1  g0108(.A(KEYINPUT74), .B(G200), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(new_n301), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT9), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(new_n283), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n273), .A2(new_n282), .A3(KEYINPUT9), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n307), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n283), .A2(new_n311), .ZN(new_n315));
  INV_X1    g0115(.A(new_n310), .ZN(new_n316));
  AND4_X1   g0116(.A1(new_n307), .A2(new_n315), .A3(new_n316), .A4(new_n313), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n306), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n289), .ZN(new_n319));
  INV_X1    g0119(.A(G232), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT81), .B1(new_n291), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT81), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n286), .A2(new_n322), .A3(G232), .A4(new_n290), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n319), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n284), .A2(KEYINPUT3), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n327), .B2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(G223), .A2(G1698), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n292), .B2(G1698), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n328), .A2(new_n330), .B1(G33), .B2(G87), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n324), .B1(new_n286), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G169), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n302), .B2(new_n332), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n206), .A2(G13), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(new_n207), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n259), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n266), .A2(new_n274), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n338), .A2(new_n339), .B1(new_n337), .B2(new_n266), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT80), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT7), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n230), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(G68), .B1(new_n328), .B2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT3), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT79), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT79), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT3), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n349), .A3(G33), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n325), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n343), .B1(new_n351), .B2(new_n207), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n342), .B1(new_n345), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT7), .B1(new_n328), .B2(G20), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n207), .A2(KEYINPUT65), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT65), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G20), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(KEYINPUT7), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n202), .B1(new_n351), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(new_n360), .A3(KEYINPUT80), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n353), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n203), .B1(new_n264), .B2(new_n202), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT16), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n254), .A2(new_n231), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n346), .A2(G33), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n325), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT7), .B1(new_n370), .B2(new_n207), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n369), .B1(new_n327), .B2(G33), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n358), .A2(new_n343), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n364), .B1(new_n374), .B2(new_n202), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n368), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n341), .B1(new_n367), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT18), .B1(new_n335), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G200), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n321), .A2(new_n323), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n289), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n331), .A2(new_n286), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n380), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n324), .B(new_n385), .C1(new_n286), .C2(new_n331), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n375), .A2(new_n376), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n255), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n365), .B1(new_n353), .B2(new_n361), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n387), .B(new_n340), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT17), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n340), .B1(new_n389), .B2(new_n390), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT18), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n395), .A3(new_n334), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n378), .A2(KEYINPUT17), .A3(new_n387), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n379), .A2(new_n393), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n337), .A2(new_n255), .ZN(new_n399));
  INV_X1    g0199(.A(new_n274), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n399), .A2(G77), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(G77), .B2(new_n278), .ZN(new_n402));
  XOR2_X1   g0202(.A(KEYINPUT8), .B(G58), .Z(new_n403));
  AOI22_X1  g0203(.A1(new_n403), .A2(new_n260), .B1(new_n358), .B2(G77), .ZN(new_n404));
  XNOR2_X1  g0204(.A(KEYINPUT15), .B(G87), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n404), .B1(new_n267), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n402), .B1(new_n406), .B2(new_n255), .ZN(new_n407));
  INV_X1    g0207(.A(G169), .ZN(new_n408));
  OAI22_X1  g0208(.A1(new_n297), .A2(new_n216), .B1(new_n223), .B2(new_n294), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n370), .A2(new_n320), .A3(G1698), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n300), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n291), .A2(new_n222), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n319), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n407), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n414), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(new_n302), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(G190), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n419), .B(KEYINPUT73), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n407), .B1(new_n416), .B2(new_n309), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR3_X1   g0222(.A1(new_n318), .A2(new_n398), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n259), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n230), .A2(G33), .A3(G77), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n260), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n427), .A2(KEYINPUT11), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n337), .A2(new_n202), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT12), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(KEYINPUT11), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n399), .A2(G68), .A3(new_n400), .ZN(new_n432));
  XNOR2_X1  g0232(.A(new_n432), .B(KEYINPUT77), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n428), .A2(new_n430), .A3(new_n431), .A4(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n292), .A2(G1698), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT75), .B1(new_n294), .B2(new_n435), .ZN(new_n436));
  AND4_X1   g0236(.A1(KEYINPUT75), .A2(new_n435), .A3(new_n325), .A4(new_n369), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n325), .A2(new_n369), .A3(G232), .A4(G1698), .ZN(new_n439));
  NAND2_X1  g0239(.A1(G33), .A2(G97), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n286), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n289), .B1(new_n291), .B2(new_n216), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT13), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n435), .A2(new_n325), .A3(new_n369), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT75), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n435), .A2(new_n325), .A3(new_n369), .A4(KEYINPUT75), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n447), .A2(new_n440), .A3(new_n439), .A4(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n443), .B1(new_n449), .B2(new_n300), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT13), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(new_n385), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n434), .B1(new_n444), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT76), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n450), .B2(new_n451), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n444), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n455), .B(KEYINPUT13), .C1(new_n442), .C2(new_n443), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(G200), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT78), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(G169), .A3(new_n458), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT14), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n457), .A2(KEYINPUT14), .A3(new_n458), .A4(G169), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n444), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n467), .A2(new_n302), .A3(new_n452), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n461), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  AOI211_X1 g0270(.A(KEYINPUT78), .B(new_n468), .C1(new_n464), .C2(new_n465), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n434), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n423), .A2(new_n460), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT83), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n222), .A2(G1698), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n351), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT4), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n350), .A2(KEYINPUT83), .A3(new_n325), .A4(new_n475), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n294), .A2(KEYINPUT4), .A3(new_n475), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n294), .A2(G250), .A3(G1698), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n286), .B1(new_n480), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n287), .A2(G1), .ZN(new_n486));
  XNOR2_X1  g0286(.A(KEYINPUT5), .B(G41), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n300), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G257), .ZN(new_n489));
  INV_X1    g0289(.A(G274), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n300), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(new_n486), .A3(new_n487), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n408), .B1(new_n485), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT83), .B1(new_n328), .B2(new_n475), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n479), .A2(new_n478), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n484), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n493), .B1(new_n497), .B2(new_n300), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n302), .ZN(new_n499));
  AOI21_X1  g0299(.A(G33), .B1(new_n347), .B2(new_n349), .ZN(new_n500));
  INV_X1    g0300(.A(new_n369), .ZN(new_n501));
  OAI211_X1 g0301(.A(KEYINPUT7), .B(new_n230), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n343), .B1(new_n294), .B2(G20), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n223), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n221), .A2(G20), .A3(G33), .ZN(new_n505));
  XNOR2_X1  g0305(.A(new_n505), .B(KEYINPUT82), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT6), .ZN(new_n507));
  INV_X1    g0307(.A(G97), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n507), .A2(new_n508), .A3(G107), .ZN(new_n509));
  XNOR2_X1  g0309(.A(G97), .B(G107), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n509), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n506), .B1(new_n230), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n255), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n278), .A2(G97), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n206), .A2(G33), .ZN(new_n515));
  AND4_X1   g0315(.A1(new_n256), .A2(new_n258), .A3(new_n278), .A4(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(G97), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n494), .A2(new_n499), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(G200), .B1(new_n485), .B2(new_n493), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n513), .A2(new_n517), .ZN(new_n521));
  INV_X1    g0321(.A(new_n493), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n482), .A2(new_n481), .A3(new_n483), .ZN(new_n523));
  INV_X1    g0323(.A(new_n496), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n477), .ZN(new_n525));
  OAI211_X1 g0325(.A(G190), .B(new_n522), .C1(new_n525), .C2(new_n286), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n520), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT84), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n520), .A2(new_n521), .A3(new_n526), .A4(KEYINPUT84), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n519), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(G257), .A2(G1698), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n532), .B1(new_n224), .B2(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n328), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n370), .A2(G303), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n286), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n488), .A2(G270), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n492), .ZN(new_n538));
  OAI21_X1  g0338(.A(G200), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(G116), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n206), .B2(G33), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n207), .A2(G116), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n399), .A2(new_n541), .B1(new_n277), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n368), .A2(new_n542), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n284), .A2(G97), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n230), .A2(new_n483), .A3(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n544), .A2(KEYINPUT20), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT20), .B1(new_n544), .B2(new_n546), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n487), .A2(new_n486), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n488), .A2(G270), .B1(new_n551), .B2(new_n491), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n328), .A2(new_n533), .B1(G303), .B2(new_n370), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n286), .B2(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n539), .B(new_n550), .C1(new_n385), .C2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n549), .A3(G169), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT21), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n554), .A2(new_n549), .A3(KEYINPUT21), .A4(G169), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n536), .A2(new_n538), .A3(new_n302), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n549), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n555), .A2(new_n558), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n278), .A2(G107), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n563), .B(KEYINPUT25), .ZN(new_n564));
  INV_X1    g0364(.A(new_n516), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(new_n223), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT22), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n567), .A2(new_n217), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n328), .A2(new_n230), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n358), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n284), .A2(new_n540), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n223), .A2(G20), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n572), .A2(new_n207), .B1(new_n573), .B2(KEYINPUT23), .ZN(new_n574));
  AND2_X1   g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n567), .B1(new_n370), .B2(new_n217), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n569), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT86), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n578), .A2(KEYINPUT24), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n368), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  XNOR2_X1  g0380(.A(KEYINPUT86), .B(KEYINPUT24), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n569), .A2(new_n575), .A3(new_n576), .A4(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n566), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n488), .A2(G264), .ZN(new_n584));
  NAND2_X1  g0384(.A1(G257), .A2(G1698), .ZN(new_n585));
  INV_X1    g0385(.A(G294), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n351), .A2(new_n585), .B1(new_n284), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT87), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n218), .A2(G1698), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n328), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n350), .A2(new_n325), .A3(new_n589), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT87), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n587), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n492), .B(new_n584), .C1(new_n593), .C2(new_n286), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n583), .B1(new_n408), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n594), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n302), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n562), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n594), .A2(G200), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n590), .A2(new_n592), .ZN(new_n600));
  INV_X1    g0400(.A(new_n585), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n328), .A2(new_n601), .B1(G33), .B2(G294), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n300), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n604), .A2(G190), .A3(new_n492), .A4(new_n584), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n599), .A2(new_n583), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n486), .A2(new_n218), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n491), .A2(new_n486), .B1(new_n286), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(G238), .A2(G1698), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n222), .B2(G1698), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n572), .B1(new_n328), .B2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n608), .B1(new_n611), .B2(new_n286), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n309), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(G190), .B2(new_n612), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n355), .A2(new_n357), .A3(G33), .A4(G97), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT19), .ZN(new_n616));
  NAND3_X1  g0416(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n355), .A2(new_n357), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n217), .A2(new_n508), .A3(new_n223), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n615), .A2(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n350), .A2(G68), .A3(new_n230), .A4(new_n325), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n368), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n405), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n623), .A2(new_n278), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT85), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n618), .A2(new_n619), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n615), .A2(new_n616), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n621), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n255), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT85), .ZN(new_n630));
  INV_X1    g0430(.A(new_n624), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n565), .A2(new_n217), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n614), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n516), .A2(new_n623), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n612), .A2(new_n408), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n302), .B(new_n608), .C1(new_n611), .C2(new_n286), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n606), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n473), .A2(new_n531), .A3(new_n598), .A4(new_n643), .ZN(G372));
  NAND2_X1  g0444(.A1(new_n393), .A2(new_n397), .ZN(new_n645));
  INV_X1    g0445(.A(new_n418), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n460), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n472), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n379), .A2(new_n396), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n648), .A2(new_n649), .B1(new_n314), .B2(new_n317), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(new_n306), .ZN(new_n651));
  INV_X1    g0451(.A(new_n473), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n639), .A2(KEYINPUT88), .ZN(new_n653));
  INV_X1    g0453(.A(new_n612), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n639), .A2(KEYINPUT88), .B1(new_n654), .B2(new_n302), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n638), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n519), .A2(new_n636), .A3(new_n642), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n657), .B2(KEYINPUT26), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT89), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n633), .B2(new_n635), .ZN(new_n660));
  AOI211_X1 g0460(.A(KEYINPUT89), .B(new_n634), .C1(new_n625), .C2(new_n632), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n614), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n638), .A2(new_n653), .A3(new_n655), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n662), .A2(new_n663), .A3(new_n519), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n595), .A2(new_n597), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n633), .A2(new_n635), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(KEYINPUT89), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n633), .A2(new_n659), .A3(new_n635), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n656), .B1(new_n675), .B2(new_n614), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(new_n531), .A3(new_n606), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT90), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n671), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n676), .A2(new_n531), .A3(KEYINPUT90), .A4(new_n606), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n666), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n651), .B1(new_n652), .B2(new_n681), .ZN(G369));
  NOR3_X1   g0482(.A1(new_n358), .A2(KEYINPUT27), .A3(new_n336), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT91), .Z(new_n684));
  INV_X1    g0484(.A(G213), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT27), .B1(new_n358), .B2(new_n336), .ZN(new_n687));
  XNOR2_X1  g0487(.A(new_n687), .B(KEYINPUT92), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G343), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n669), .B(new_n555), .C1(new_n691), .C2(new_n550), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n690), .A2(G343), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(new_n549), .A3(new_n668), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT93), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n667), .A2(new_n693), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n606), .B1(new_n691), .B2(new_n583), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n667), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n693), .A2(new_n669), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n698), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n212), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n619), .A2(G116), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT94), .Z(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n228), .B2(new_n707), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n664), .B1(new_n657), .B2(KEYINPUT26), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n676), .A2(new_n519), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(KEYINPUT26), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n676), .A2(new_n531), .A3(new_n670), .A4(new_n606), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .A3(new_n691), .ZN(new_n718));
  INV_X1    g0518(.A(new_n519), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n518), .B1(G190), .B2(new_n498), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT84), .B1(new_n720), .B2(new_n520), .ZN(new_n721));
  INV_X1    g0521(.A(new_n530), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n662), .A2(new_n606), .A3(new_n664), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n678), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n680), .A3(new_n670), .ZN(new_n726));
  INV_X1    g0526(.A(new_n666), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n693), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n718), .B1(new_n728), .B2(KEYINPUT29), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT95), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n554), .A2(new_n302), .A3(new_n612), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n522), .B1(new_n525), .B2(new_n286), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n730), .B1(new_n733), .B2(new_n596), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n554), .A2(new_n612), .A3(new_n302), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n603), .A2(new_n300), .B1(G264), .B2(new_n488), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n735), .A2(new_n498), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT30), .A4(new_n498), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n731), .A2(new_n732), .A3(new_n594), .A4(KEYINPUT95), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n734), .A2(new_n739), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n693), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT31), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n691), .A2(new_n744), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n739), .B(new_n740), .C1(new_n596), .C2(new_n733), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n743), .A2(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n531), .A2(new_n598), .A3(new_n643), .A4(new_n691), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G330), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n729), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n712), .B1(new_n752), .B2(G1), .ZN(G364));
  NOR2_X1   g0553(.A1(new_n358), .A2(new_n276), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G45), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G1), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n706), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n697), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n758), .B1(G330), .B2(new_n696), .ZN(new_n759));
  INV_X1    g0559(.A(new_n757), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n705), .A2(new_n370), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n761), .A2(G355), .B1(new_n540), .B2(new_n705), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n328), .B(new_n705), .C1(new_n287), .C2(new_n229), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n764), .A2(KEYINPUT96), .B1(new_n252), .B2(new_n287), .ZN(new_n765));
  AND2_X1   g0565(.A1(new_n764), .A2(KEYINPUT96), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n231), .B1(G20), .B2(new_n408), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n767), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n309), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G20), .A3(G190), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT100), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n230), .A2(G190), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT97), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n302), .A2(G200), .ZN(new_n783));
  AND3_X1   g0583(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n782), .B1(new_n781), .B2(new_n783), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n780), .A2(G303), .B1(G311), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G179), .A2(G200), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT99), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n781), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT103), .B(G326), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n302), .A2(new_n380), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n358), .A2(G190), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n792), .A2(G329), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n781), .A2(new_n794), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT33), .B(G317), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n358), .A2(G190), .A3(new_n783), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n799), .A2(new_n800), .B1(G322), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n781), .A2(new_n774), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n370), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OR2_X1    g0606(.A1(new_n790), .A2(new_n230), .ZN(new_n807));
  INV_X1    g0607(.A(new_n781), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n806), .B1(new_n810), .B2(G294), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n788), .A2(new_n797), .A3(new_n803), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n780), .A2(G87), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n813), .B(new_n294), .C1(new_n223), .C2(new_n804), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(KEYINPUT101), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n786), .A2(new_n221), .B1(new_n264), .B2(new_n801), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT98), .Z(new_n817));
  INV_X1    g0617(.A(G159), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n791), .A2(KEYINPUT32), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(KEYINPUT32), .B1(new_n791), .B2(new_n818), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n247), .B2(new_n795), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n809), .A2(new_n508), .B1(new_n202), .B2(new_n798), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n819), .B(new_n821), .C1(new_n822), .C2(KEYINPUT102), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n817), .B(new_n823), .C1(KEYINPUT102), .C2(new_n822), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n812), .B1(new_n815), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n760), .B(new_n773), .C1(new_n771), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n770), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n826), .B1(new_n695), .B2(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n759), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G396));
  NOR2_X1   g0630(.A1(new_n420), .A2(new_n421), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n691), .A2(new_n407), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n418), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n646), .A2(new_n691), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n422), .A2(new_n693), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n728), .A2(new_n836), .B1(new_n681), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n750), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n760), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n838), .A2(new_n750), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n771), .A2(new_n768), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n760), .B1(new_n221), .B2(new_n842), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G137), .A2(new_n796), .B1(new_n802), .B2(G143), .ZN(new_n844));
  INV_X1    g0644(.A(G150), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n844), .B1(new_n845), .B2(new_n798), .C1(new_n786), .C2(new_n818), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT34), .ZN(new_n847));
  INV_X1    g0647(.A(new_n804), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n351), .B1(new_n848), .B2(G68), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n849), .B1(new_n850), .B2(new_n791), .C1(new_n264), .C2(new_n809), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(G50), .B2(new_n780), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n370), .B1(new_n586), .B2(new_n801), .C1(new_n809), .C2(new_n508), .ZN(new_n853));
  INV_X1    g0653(.A(G311), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n791), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n804), .A2(new_n217), .ZN(new_n856));
  INV_X1    g0656(.A(G303), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n798), .A2(new_n805), .B1(new_n857), .B2(new_n795), .ZN(new_n858));
  NOR4_X1   g0658(.A1(new_n853), .A2(new_n855), .A3(new_n856), .A4(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n780), .A2(G107), .B1(G116), .B2(new_n787), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n847), .A2(new_n852), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT104), .Z(new_n862));
  INV_X1    g0662(.A(new_n771), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n843), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n836), .A2(new_n769), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n840), .A2(new_n841), .B1(new_n864), .B2(new_n865), .ZN(G384));
  NOR2_X1   g0666(.A1(new_n754), .A2(new_n206), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT40), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT107), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n743), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n742), .A2(KEYINPUT107), .A3(new_n693), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n744), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n742), .A2(new_n745), .ZN(new_n873));
  AND2_X1   g0673(.A1(new_n748), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n693), .A2(new_n434), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n472), .A2(new_n460), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n876), .B1(new_n472), .B2(new_n460), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n836), .B(new_n875), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n367), .A2(new_n259), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT16), .B1(new_n362), .B2(new_n364), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n340), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n690), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n398), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT105), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n345), .A2(new_n352), .A3(new_n342), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT80), .B1(new_n354), .B2(new_n360), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n364), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n376), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n390), .A2(new_n424), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n341), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n391), .B1(new_n892), .B2(new_n689), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n335), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n886), .B(KEYINPUT37), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n394), .A2(new_n334), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n394), .A2(new_n690), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n896), .A2(new_n897), .A3(new_n898), .A4(new_n391), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n882), .A2(new_n334), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n883), .A3(new_n391), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n886), .B1(new_n902), .B2(KEYINPUT37), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n885), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT38), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n893), .B2(new_n894), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(KEYINPUT105), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(new_n899), .A3(new_n895), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n905), .B1(new_n398), .B2(new_n884), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n904), .A2(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n868), .B1(new_n879), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n909), .B1(new_n900), .B2(new_n903), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n391), .B1(new_n335), .B2(new_n378), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n378), .A2(new_n689), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT37), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n899), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n398), .A2(new_n914), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n905), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n868), .B1(new_n912), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n466), .A2(new_n469), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT78), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n466), .A2(new_n461), .A3(new_n469), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n460), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n434), .B(new_n693), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n472), .A2(new_n460), .A3(new_n876), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n920), .A2(new_n928), .A3(new_n836), .A4(new_n875), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n911), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g0730(.A1(new_n473), .A2(new_n875), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(G330), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n934), .A2(KEYINPUT108), .B1(new_n930), .B2(new_n931), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(KEYINPUT108), .B2(new_n934), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n908), .B2(new_n885), .ZN(new_n937));
  INV_X1    g0737(.A(new_n912), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT39), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n912), .A2(new_n919), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT106), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT106), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n912), .A2(new_n919), .A3(new_n943), .A4(new_n940), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n939), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n924), .A2(new_n434), .A3(new_n691), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n834), .B1(new_n681), .B2(new_n837), .ZN(new_n949));
  INV_X1    g0749(.A(new_n910), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(new_n950), .A3(new_n928), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n649), .A2(new_n689), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n948), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n718), .B(new_n473), .C1(KEYINPUT29), .C2(new_n728), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n651), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n953), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n867), .B1(new_n936), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n956), .B2(new_n936), .ZN(new_n958));
  INV_X1    g0758(.A(new_n511), .ZN(new_n959));
  OR2_X1    g0759(.A1(new_n959), .A2(KEYINPUT35), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(KEYINPUT35), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n960), .A2(G116), .A3(new_n232), .A4(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT36), .ZN(new_n963));
  INV_X1    g0763(.A(new_n228), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n964), .B(G77), .C1(new_n202), .C2(new_n264), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n248), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(G1), .A3(new_n276), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n958), .A2(new_n963), .A3(new_n967), .ZN(G367));
  OAI21_X1  g0768(.A(new_n531), .B1(new_n521), .B2(new_n691), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n693), .A2(new_n519), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OR3_X1    g0772(.A1(new_n701), .A2(KEYINPUT112), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT112), .B1(new_n701), .B2(new_n972), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n675), .A2(new_n691), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n664), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n676), .B2(new_n976), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT109), .Z(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n667), .B1(new_n529), .B2(new_n530), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n691), .B1(new_n981), .B2(new_n519), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT110), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n700), .A2(new_n702), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n983), .B1(new_n972), .B2(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n971), .A2(new_n700), .A3(KEYINPUT110), .A4(new_n702), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT42), .ZN(new_n988));
  OAI211_X1 g0788(.A(KEYINPUT111), .B(new_n982), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT111), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n988), .B1(new_n985), .B2(new_n986), .ZN(new_n991));
  INV_X1    g0791(.A(new_n982), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n987), .A2(new_n988), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n989), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n975), .A2(new_n980), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n975), .B1(new_n980), .B2(new_n995), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n997), .A2(new_n998), .B1(KEYINPUT43), .B2(new_n979), .ZN(new_n999));
  INV_X1    g0799(.A(new_n756), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT45), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n698), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n984), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1001), .B1(new_n1003), .B2(new_n972), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n703), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1003), .A2(KEYINPUT44), .A3(new_n972), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT44), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n703), .B2(new_n971), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n1006), .A2(new_n701), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n701), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n700), .B(new_n702), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n697), .B(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n751), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n706), .B(KEYINPUT41), .Z(new_n1017));
  OAI21_X1  g0817(.A(new_n1000), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n975), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n995), .A2(new_n980), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1021), .A2(new_n1022), .A3(new_n996), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n999), .A2(new_n1018), .A3(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n705), .A2(new_n328), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n242), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n772), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n705), .B2(new_n623), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n760), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(G143), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n294), .B1(new_n1030), .B2(new_n795), .C1(new_n809), .C2(new_n202), .ZN(new_n1031));
  INV_X1    g0831(.A(G137), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n791), .A2(new_n1032), .B1(new_n845), .B2(new_n801), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n804), .A2(new_n221), .B1(new_n798), .B2(new_n818), .ZN(new_n1034));
  NOR3_X1   g0834(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n247), .B2(new_n786), .C1(new_n264), .C2(new_n779), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n351), .B1(new_n586), .B2(new_n798), .C1(new_n809), .C2(new_n223), .ZN(new_n1037));
  INV_X1    g0837(.A(G317), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n791), .A2(new_n1038), .B1(new_n854), .B2(new_n795), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n804), .A2(new_n508), .B1(new_n857), .B2(new_n801), .ZN(new_n1040));
  NOR3_X1   g0840(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n805), .B2(new_n786), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n779), .A2(new_n540), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT46), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1036), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  XOR2_X1   g0845(.A(new_n1045), .B(KEYINPUT47), .Z(new_n1046));
  OAI221_X1 g0846(.A(new_n1029), .B1(new_n863), .B2(new_n1046), .C1(new_n979), .C2(new_n827), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT113), .Z(new_n1048));
  NAND2_X1  g0848(.A1(new_n1024), .A2(new_n1048), .ZN(G387));
  OAI21_X1  g0849(.A(new_n1025), .B1(new_n239), .B2(new_n287), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n761), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1050), .B1(new_n709), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n287), .B1(new_n202), .B2(new_n221), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n403), .A2(new_n247), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1053), .B1(new_n1054), .B2(KEYINPUT50), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n709), .B(new_n1055), .C1(KEYINPUT50), .C2(new_n1054), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1052), .A2(new_n1056), .B1(new_n223), .B2(new_n705), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n757), .B1(new_n1057), .B2(new_n1027), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT114), .Z(new_n1059));
  NOR2_X1   g0859(.A1(new_n809), .A2(new_n405), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n791), .A2(new_n845), .B1(new_n247), .B2(new_n801), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n798), .A2(new_n266), .B1(new_n818), .B2(new_n795), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n328), .B1(new_n804), .B2(new_n508), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n202), .B2(new_n786), .C1(new_n221), .C2(new_n779), .ZN(new_n1065));
  INV_X1    g0865(.A(G322), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n798), .A2(new_n854), .B1(new_n1066), .B2(new_n795), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT116), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n857), .B2(new_n786), .C1(new_n1038), .C2(new_n801), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n779), .A2(new_n586), .B1(new_n809), .B2(new_n805), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT115), .Z(new_n1074));
  NAND3_X1  g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(KEYINPUT117), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n351), .B1(new_n804), .B2(new_n540), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n792), .B2(new_n793), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1076), .A2(KEYINPUT117), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1065), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1059), .B1(new_n1082), .B2(new_n771), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT118), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n700), .A2(new_n827), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1085), .A2(new_n1087), .B1(new_n756), .B2(new_n1015), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n752), .A2(new_n1015), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n706), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n752), .A2(new_n1015), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(G393));
  OAI21_X1  g0892(.A(new_n772), .B1(new_n212), .B2(new_n508), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1025), .B2(new_n246), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n760), .A2(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n779), .A2(new_n805), .B1(new_n586), .B2(new_n786), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G322), .A2(new_n792), .B1(new_n799), .B2(G303), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n370), .C1(new_n223), .C2(new_n804), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n854), .A2(new_n801), .B1(new_n795), .B2(new_n1038), .ZN(new_n1099));
  XOR2_X1   g0899(.A(new_n1099), .B(KEYINPUT52), .Z(new_n1100));
  NOR2_X1   g0900(.A1(new_n809), .A2(new_n540), .ZN(new_n1101));
  NOR4_X1   g0901(.A1(new_n1096), .A2(new_n1098), .A3(new_n1100), .A4(new_n1101), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1102), .A2(KEYINPUT119), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(KEYINPUT119), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n809), .A2(new_n221), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n791), .A2(new_n1030), .B1(new_n798), .B2(new_n247), .ZN(new_n1106));
  NOR4_X1   g0906(.A1(new_n1105), .A2(new_n351), .A3(new_n856), .A4(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n845), .A2(new_n795), .B1(new_n801), .B2(new_n818), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT51), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n780), .A2(G68), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n787), .A2(new_n403), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1103), .A2(new_n1104), .A3(new_n1112), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1095), .B1(new_n827), .B2(new_n971), .C1(new_n1113), .C2(new_n863), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1013), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n706), .B1(new_n1115), .B2(new_n1089), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1013), .B1(new_n752), .B2(new_n1015), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n1114), .B1(new_n1000), .B2(new_n1115), .C1(new_n1116), .C2(new_n1117), .ZN(G390));
  AOI21_X1  g0918(.A(new_n947), .B1(new_n912), .B2(new_n919), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n834), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n693), .B1(new_n715), .B2(new_n716), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n833), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n877), .A2(new_n878), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1119), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n947), .B1(new_n949), .B2(new_n928), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n945), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n933), .B1(new_n872), .B2(new_n874), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n928), .A2(new_n836), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n928), .A2(G330), .A3(new_n749), .A4(new_n836), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n1124), .B(new_n1131), .C1(new_n945), .C2(new_n1125), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n756), .A3(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n294), .B(new_n1105), .C1(G68), .C2(new_n848), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n791), .A2(new_n586), .B1(new_n798), .B2(new_n223), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n540), .A2(new_n801), .B1(new_n795), .B2(new_n805), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n787), .A2(G97), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1134), .A2(new_n813), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n809), .A2(new_n818), .B1(new_n1032), .B2(new_n798), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(KEYINPUT54), .B(G143), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1140), .B1(new_n787), .B2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT120), .ZN(new_n1144));
  XOR2_X1   g0944(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1145));
  OR3_X1    g0945(.A1(new_n779), .A2(new_n845), .A3(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n779), .B2(new_n845), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n294), .B1(new_n804), .B2(new_n247), .ZN(new_n1148));
  INV_X1    g0948(.A(G125), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n791), .A2(new_n1149), .B1(new_n850), .B2(new_n801), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1148), .B(new_n1150), .C1(G128), .C2(new_n796), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1146), .A2(new_n1147), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1139), .B1(new_n1144), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n771), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n760), .B1(new_n266), .B2(new_n842), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n945), .C2(new_n769), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1133), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n473), .A2(new_n1127), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n954), .A2(new_n306), .A3(new_n650), .A4(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n927), .B(new_n926), .C1(new_n750), .C2(new_n835), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1128), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n949), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1127), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1123), .B1(new_n1164), .B2(new_n835), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n1122), .A3(new_n1131), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1160), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n707), .B1(new_n1158), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1130), .A2(new_n1132), .A3(new_n1167), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1157), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(G378));
  AOI221_X4 g0972(.A(new_n835), .B1(new_n872), .B2(new_n874), .C1(new_n926), .C2(new_n927), .ZN(new_n1173));
  AOI21_X1  g0973(.A(KEYINPUT40), .B1(new_n1173), .B2(new_n950), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n929), .A2(G330), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n690), .A2(new_n283), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n318), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n318), .A2(new_n1177), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  OR3_X1    g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1174), .A2(new_n1175), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n933), .B1(new_n1173), .B2(new_n920), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1184), .B1(new_n1187), .B2(new_n911), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n953), .B1(new_n1186), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1185), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n837), .B1(new_n726), .B2(new_n727), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n1191), .A2(new_n1120), .B1(new_n877), .B2(new_n878), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n952), .B1(new_n1192), .B2(new_n910), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n947), .B2(new_n945), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1187), .A2(new_n911), .A3(new_n1184), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1190), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1189), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n756), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1185), .A2(new_n768), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n842), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n757), .B1(G50), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n351), .A2(new_n285), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n804), .A2(new_n264), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(G283), .C2(new_n792), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n221), .B2(new_n779), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT122), .Z(new_n1206));
  AOI22_X1  g1006(.A1(new_n799), .A2(G97), .B1(G116), .B2(new_n796), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n223), .B2(new_n801), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G68), .B2(new_n810), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1206), .B(new_n1209), .C1(new_n405), .C2(new_n786), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT58), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1202), .B(new_n247), .C1(G33), .C2(G41), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n780), .A2(new_n1142), .B1(G137), .B2(new_n787), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n798), .A2(new_n850), .B1(new_n1149), .B2(new_n795), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(G128), .B2(new_n802), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1215), .B(new_n1217), .C1(new_n845), .C2(new_n809), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n848), .A2(G159), .ZN(new_n1221));
  AOI211_X1 g1021(.A(G33), .B(G41), .C1(new_n792), .C2(G124), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1201), .B1(new_n1224), .B2(new_n771), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1199), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1198), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1160), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1170), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n1197), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT57), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n706), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1230), .A2(new_n1197), .A3(KEYINPUT57), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1228), .B1(new_n1234), .B2(new_n1236), .ZN(G375));
  OAI21_X1  g1037(.A(new_n757), .B1(G68), .B2(new_n1200), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n780), .A2(G159), .B1(G150), .B2(new_n787), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n351), .B(new_n1203), .C1(new_n810), .C2(G50), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n799), .A2(new_n1142), .B1(G132), .B2(new_n796), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n792), .A2(G128), .B1(G137), .B2(new_n802), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n294), .B(new_n1060), .C1(G77), .C2(new_n848), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n799), .A2(G116), .B1(G294), .B2(new_n796), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n792), .A2(G303), .B1(G283), .B2(new_n802), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n779), .A2(new_n508), .B1(new_n223), .B2(new_n786), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1243), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1238), .B1(new_n1249), .B2(new_n771), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n928), .B2(new_n769), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1253), .B2(new_n1000), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1167), .A2(new_n1017), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1160), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1254), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(G381));
  NOR4_X1   g1058(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n1257), .ZN(new_n1260));
  OR4_X1    g1060(.A1(G387), .A2(new_n1260), .A3(G375), .A4(G378), .ZN(G407));
  NOR2_X1   g1061(.A1(new_n685), .A2(G343), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  OR3_X1    g1063(.A1(G375), .A2(G378), .A3(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(G407), .A2(new_n1264), .A3(G213), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1265), .B(KEYINPUT123), .ZN(G409));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1256), .B1(new_n1267), .B2(new_n1167), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1252), .A2(new_n1267), .A3(new_n1229), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(new_n707), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1254), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  OR2_X1    g1071(.A1(new_n1271), .A2(G384), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(G384), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1231), .A2(new_n1017), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT124), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1190), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1194), .B1(new_n1190), .B2(new_n1195), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1189), .A2(KEYINPUT124), .A3(new_n1196), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n756), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n1226), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1275), .B1(new_n1282), .B2(KEYINPUT125), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT125), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1281), .A2(new_n1284), .A3(new_n1226), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G378), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n707), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1171), .B(new_n1227), .C1(new_n1287), .C2(new_n1235), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1263), .B(new_n1274), .C1(new_n1286), .C2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(KEYINPUT62), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G378), .B(new_n1228), .C1(new_n1234), .C2(new_n1236), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1281), .A2(new_n1284), .A3(new_n1226), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1284), .B1(new_n1281), .B2(new_n1226), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n1292), .A2(new_n1293), .A3(new_n1275), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1291), .B1(new_n1294), .B2(G378), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT62), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1295), .A2(new_n1296), .A3(new_n1263), .A4(new_n1274), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1262), .A2(G2897), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1298), .B(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1282), .A2(KEYINPUT125), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1275), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1301), .A2(new_n1285), .A3(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1288), .B1(new_n1303), .B2(new_n1171), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1300), .B1(new_n1304), .B2(new_n1262), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1290), .A2(new_n1297), .A3(new_n1305), .A4(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT126), .ZN(new_n1308));
  INV_X1    g1108(.A(G390), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G387), .A2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1024), .A2(G390), .A3(new_n1048), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(G393), .B(G396), .ZN(new_n1312));
  AND4_X1   g1112(.A1(new_n1308), .A2(new_n1310), .A3(new_n1311), .A4(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(KEYINPUT126), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n1314), .A2(new_n1312), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1313), .A2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1307), .A2(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(KEYINPUT61), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT63), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1289), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1295), .A2(KEYINPUT63), .A3(new_n1263), .A4(new_n1274), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1318), .A2(new_n1320), .A3(new_n1305), .A4(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1317), .A2(new_n1322), .ZN(G405));
  NAND2_X1  g1123(.A1(G375), .A2(new_n1171), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1291), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1316), .A2(new_n1325), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1291), .B(new_n1324), .C1(new_n1313), .C2(new_n1315), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1326), .A2(new_n1274), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1274), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(G402));
endmodule


