//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1017, new_n1018, new_n1019, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT86), .Z(new_n190));
  INV_X1    g004(.A(KEYINPUT78), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G104), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT78), .A3(G107), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n192), .A2(KEYINPUT3), .A3(G104), .ZN(new_n196));
  AOI21_X1  g010(.A(KEYINPUT3), .B1(new_n192), .B2(G104), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n193), .B(new_n195), .C1(new_n196), .C2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT4), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n198), .A2(new_n199), .A3(G101), .ZN(new_n200));
  INV_X1    g014(.A(G116), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G119), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n201), .A2(KEYINPUT67), .A3(G119), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT67), .B1(new_n201), .B2(G119), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT68), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G116), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n201), .A2(KEYINPUT67), .A3(G119), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n202), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n215));
  INV_X1    g029(.A(G113), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT66), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(KEYINPUT2), .B2(G113), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n215), .B2(new_n216), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n207), .A2(new_n214), .A3(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n212), .B(new_n220), .C1(new_n215), .C2(new_n216), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n200), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n194), .B2(G107), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n192), .A2(KEYINPUT3), .A3(G104), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT79), .B(G101), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n228), .A2(new_n229), .A3(new_n193), .A4(new_n195), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT80), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n193), .A2(new_n195), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n233), .A2(KEYINPUT80), .A3(new_n229), .A4(new_n228), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n199), .B1(new_n198), .B2(G101), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n224), .A2(new_n237), .ZN(new_n238));
  AOI211_X1 g052(.A(KEYINPUT68), .B(new_n202), .C1(new_n210), .C2(new_n211), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n210), .A2(new_n211), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n213), .B1(new_n240), .B2(new_n203), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT5), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT5), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n216), .B1(new_n202), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n194), .A2(G107), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n192), .A2(G104), .ZN(new_n247));
  OAI21_X1  g061(.A(G101), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n249), .B1(new_n232), .B2(new_n234), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n245), .A2(new_n223), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n238), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G110), .B(G122), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n238), .A2(new_n251), .A3(new_n253), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n255), .A2(KEYINPUT6), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT6), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n252), .A2(new_n258), .A3(new_n254), .ZN(new_n259));
  INV_X1    g073(.A(G143), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT1), .B1(new_n260), .B2(G146), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(G146), .ZN(new_n262));
  INV_X1    g076(.A(G146), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(G143), .ZN(new_n264));
  OAI211_X1 g078(.A(G128), .B(new_n261), .C1(new_n262), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(G143), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(G146), .ZN(new_n267));
  INV_X1    g081(.A(G128), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n266), .B(new_n267), .C1(KEYINPUT1), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G125), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n266), .A2(new_n267), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G143), .B(G146), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT0), .B(G128), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G125), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G224), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(G953), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n279), .B(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n257), .A2(new_n259), .A3(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n244), .B1(new_n206), .B2(new_n243), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n223), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n250), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n253), .B(KEYINPUT8), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n243), .B1(new_n207), .B2(new_n214), .ZN(new_n289));
  INV_X1    g103(.A(new_n244), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n223), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n287), .B(new_n288), .C1(new_n291), .C2(new_n250), .ZN(new_n292));
  INV_X1    g106(.A(new_n278), .ZN(new_n293));
  AOI21_X1  g107(.A(G125), .B1(new_n265), .B2(new_n269), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n281), .B2(KEYINPUT84), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(KEYINPUT84), .B2(new_n281), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n293), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n272), .A2(KEYINPUT83), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT83), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n294), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n278), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT7), .B1(new_n280), .B2(G953), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n298), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n292), .A2(new_n304), .A3(KEYINPUT85), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n256), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT85), .B1(new_n292), .B2(new_n304), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n284), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n190), .B1(new_n283), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n257), .A2(new_n259), .A3(new_n282), .ZN(new_n310));
  INV_X1    g124(.A(new_n307), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n256), .A3(new_n305), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n310), .A2(new_n312), .A3(new_n284), .A4(new_n189), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n188), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G113), .B(G122), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n194), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(G104), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(G237), .A2(G953), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n321), .A2(G143), .A3(G214), .ZN(new_n322));
  AOI21_X1  g136(.A(G143), .B1(new_n321), .B2(G214), .ZN(new_n323));
  OAI21_X1  g137(.A(G131), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT17), .ZN(new_n325));
  INV_X1    g139(.A(G237), .ZN(new_n326));
  INV_X1    g140(.A(G953), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(G214), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n260), .ZN(new_n329));
  INV_X1    g143(.A(G131), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n321), .A2(G143), .A3(G214), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n324), .A2(new_n325), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT16), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(new_n335), .A3(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n271), .A2(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n336), .B1(new_n339), .B2(new_n334), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n263), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n330), .B1(new_n329), .B2(new_n331), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(KEYINPUT17), .ZN(new_n343));
  OAI211_X1 g157(.A(G146), .B(new_n336), .C1(new_n339), .C2(new_n334), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n333), .A2(new_n341), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n337), .A2(new_n338), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n263), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(G146), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT87), .A2(KEYINPUT18), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n329), .B(new_n331), .C1(new_n330), .C2(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n349), .B(new_n351), .C1(new_n324), .C2(new_n350), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n320), .B1(new_n345), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n319), .A2(KEYINPUT90), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT90), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n317), .A2(new_n356), .A3(new_n318), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(new_n345), .A3(new_n352), .ZN(new_n359));
  AOI21_X1  g173(.A(G902), .B1(new_n354), .B2(new_n359), .ZN(new_n360));
  XOR2_X1   g174(.A(KEYINPUT92), .B(G475), .Z(new_n361));
  NOR2_X1   g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(G475), .A2(G902), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT19), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT19), .B1(new_n337), .B2(new_n338), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n263), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT89), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n344), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n346), .A2(KEYINPUT16), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(KEYINPUT76), .A3(G146), .A4(new_n336), .ZN(new_n374));
  OAI211_X1 g188(.A(KEYINPUT89), .B(new_n263), .C1(new_n366), .C2(new_n367), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n370), .A2(new_n372), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n322), .A2(new_n323), .A3(G131), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT88), .B1(new_n377), .B2(new_n342), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT88), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n324), .A2(new_n379), .A3(new_n332), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n352), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n319), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n365), .B1(new_n383), .B2(new_n359), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT91), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n324), .A2(new_n379), .A3(new_n332), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n379), .B1(new_n324), .B2(new_n332), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT19), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n339), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT19), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT89), .B1(new_n392), .B2(new_n263), .ZN(new_n393));
  INV_X1    g207(.A(new_n375), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n374), .A2(new_n372), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n388), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n320), .B1(new_n397), .B2(new_n352), .ZN(new_n398));
  INV_X1    g212(.A(new_n359), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n385), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT20), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n384), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n345), .A2(new_n352), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n319), .A2(new_n382), .B1(new_n403), .B2(new_n358), .ZN(new_n404));
  NOR4_X1   g218(.A1(new_n404), .A2(new_n385), .A3(KEYINPUT20), .A4(new_n365), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n363), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G478), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(KEYINPUT15), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n260), .A2(G128), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n268), .A2(G143), .ZN(new_n411));
  INV_X1    g225(.A(G134), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT95), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT13), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT94), .B1(new_n410), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n410), .A2(new_n415), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT94), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n418), .A2(new_n260), .A3(KEYINPUT13), .A4(G128), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n416), .A2(new_n417), .A3(new_n411), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G134), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT93), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n201), .B2(G122), .ZN(new_n423));
  INV_X1    g237(.A(G122), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(KEYINPUT93), .A3(G116), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n201), .A2(G122), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n192), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n192), .B1(new_n426), .B2(new_n427), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n414), .B(new_n421), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n427), .B(KEYINPUT14), .ZN(new_n432));
  INV_X1    g246(.A(new_n426), .ZN(new_n433));
  OAI21_X1  g247(.A(G107), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n410), .A2(new_n411), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G134), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n413), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n428), .A3(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT9), .B(G234), .ZN(new_n439));
  INV_X1    g253(.A(G217), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n439), .A2(new_n440), .A3(G953), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n431), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT96), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT96), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n431), .A2(new_n444), .A3(new_n438), .A4(new_n441), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n431), .A2(new_n438), .ZN(new_n446));
  INV_X1    g260(.A(new_n441), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n409), .B1(new_n449), .B2(new_n284), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n284), .A3(new_n409), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G952), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(G953), .ZN(new_n455));
  INV_X1    g269(.A(G234), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n455), .B1(new_n456), .B2(new_n326), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(G902), .B(G953), .C1(new_n456), .C2(new_n326), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT97), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT21), .B(G898), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n406), .A2(new_n453), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n314), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT32), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n321), .A2(G210), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT27), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT26), .B(G101), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT11), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(new_n412), .B2(G137), .ZN(new_n471));
  INV_X1    g285(.A(G137), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(KEYINPUT11), .A3(G134), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n412), .A2(G137), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(KEYINPUT64), .A2(G131), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n471), .A2(new_n473), .A3(new_n476), .A4(new_n474), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT65), .ZN(new_n481));
  XNOR2_X1  g295(.A(G134), .B(G137), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n481), .B1(new_n482), .B2(new_n330), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n471), .A2(new_n473), .A3(new_n330), .A4(new_n474), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n412), .A2(G137), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n472), .A2(G134), .ZN(new_n486));
  OAI211_X1 g300(.A(KEYINPUT65), .B(G131), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  OAI22_X1  g302(.A1(new_n480), .A2(new_n277), .B1(new_n488), .B2(new_n270), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n222), .A2(new_n223), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n265), .A2(new_n269), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(new_n484), .A3(new_n483), .A4(new_n487), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n478), .A2(new_n479), .ZN(new_n494));
  INV_X1    g308(.A(new_n277), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n493), .A2(new_n496), .B1(new_n222), .B2(new_n223), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT28), .B1(new_n491), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n488), .A2(new_n270), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n277), .B1(new_n478), .B2(new_n479), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n222), .A2(new_n223), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT28), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n469), .B1(new_n498), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n493), .B2(new_n496), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT30), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n490), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n503), .A3(new_n469), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT31), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT30), .B1(new_n499), .B2(new_n500), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n496), .B(new_n507), .C1(new_n270), .C2(new_n488), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n491), .B1(new_n516), .B2(new_n490), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(KEYINPUT31), .A3(new_n469), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n506), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(G472), .A2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n465), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT69), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n469), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n489), .A2(new_n490), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n504), .B1(new_n503), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n491), .A2(KEYINPUT28), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT31), .B1(new_n517), .B2(new_n469), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n502), .B1(new_n514), .B2(new_n515), .ZN(new_n531));
  NOR4_X1   g345(.A1(new_n531), .A2(new_n512), .A3(new_n491), .A4(new_n525), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n529), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n520), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(KEYINPUT69), .A3(new_n465), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(KEYINPUT32), .A3(new_n520), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT29), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n525), .B1(new_n498), .B2(new_n505), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n531), .A2(new_n491), .A3(new_n469), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT70), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n505), .A2(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n527), .A2(new_n528), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n543), .B2(new_n541), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n469), .A2(KEYINPUT29), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n540), .B(new_n284), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(G472), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n524), .A2(new_n535), .A3(new_n536), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n341), .A2(new_n344), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n209), .A2(G128), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n268), .A2(G119), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT24), .B(G110), .ZN(new_n553));
  OR3_X1    g367(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT71), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT71), .B1(new_n552), .B2(new_n553), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G110), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n550), .A2(KEYINPUT23), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(KEYINPUT72), .A3(new_n551), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n209), .A2(G128), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT72), .ZN(new_n561));
  OAI211_X1 g375(.A(KEYINPUT23), .B(new_n550), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n549), .B(new_n556), .C1(new_n557), .C2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT22), .B(G137), .ZN(new_n565));
  INV_X1    g379(.A(G221), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n566), .A2(new_n456), .A3(G953), .ZN(new_n567));
  XOR2_X1   g381(.A(new_n565), .B(new_n567), .Z(new_n568));
  XOR2_X1   g382(.A(KEYINPUT73), .B(G110), .Z(new_n569));
  NAND3_X1  g383(.A1(new_n559), .A2(new_n562), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT74), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(new_n552), .B2(new_n553), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n552), .A2(new_n553), .A3(new_n571), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(KEYINPUT75), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT75), .ZN(new_n577));
  INV_X1    g391(.A(new_n574), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n572), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n577), .B1(new_n579), .B2(new_n570), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n374), .A2(new_n372), .A3(new_n347), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n564), .B(new_n568), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n568), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n575), .A2(KEYINPUT75), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n579), .A2(new_n577), .A3(new_n570), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n582), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n564), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n583), .A2(new_n589), .A3(new_n284), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT25), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT25), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n583), .A2(new_n589), .A3(new_n592), .A4(new_n284), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n440), .B1(G234), .B2(new_n284), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n594), .A2(G902), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n583), .A2(new_n589), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(KEYINPUT77), .ZN(new_n598));
  OR2_X1    g412(.A1(new_n597), .A2(KEYINPUT77), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n439), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n566), .B1(new_n602), .B2(new_n284), .ZN(new_n603));
  INV_X1    g417(.A(G469), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(new_n284), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n265), .A2(new_n269), .A3(new_n248), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n235), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT81), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n606), .B1(new_n232), .B2(new_n234), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT81), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n610), .A2(new_n611), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n200), .A2(new_n277), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n237), .A2(new_n615), .B1(new_n612), .B2(KEYINPUT10), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n480), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n235), .A2(new_n248), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n270), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n610), .A2(new_n619), .A3(new_n613), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT82), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT12), .B1(new_n494), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n620), .A2(new_n494), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n620), .B2(new_n494), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n617), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(G110), .B(G140), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n327), .A2(G227), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n617), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n612), .A2(KEYINPUT81), .ZN(new_n633));
  AOI211_X1 g447(.A(new_n609), .B(new_n606), .C1(new_n232), .C2(new_n234), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n633), .A2(new_n634), .A3(KEYINPUT10), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n237), .A2(new_n615), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n612), .A2(KEYINPUT10), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n494), .B1(new_n635), .B2(new_n638), .ZN(new_n639));
  AOI22_X1  g453(.A1(new_n626), .A2(new_n629), .B1(new_n632), .B2(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n605), .B1(new_n640), .B2(G469), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n620), .A2(new_n494), .A3(new_n623), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n250), .A2(new_n492), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n643), .A2(new_n633), .A3(new_n634), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n622), .B1(new_n644), .B2(new_n480), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n631), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n630), .B1(new_n639), .B2(new_n617), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n604), .B(new_n284), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n603), .B1(new_n641), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n464), .A2(new_n548), .A3(new_n601), .A4(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(new_n229), .Z(G3));
  INV_X1    g465(.A(new_n189), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n652), .B1(new_n283), .B2(new_n308), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n188), .B1(new_n653), .B2(new_n313), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT91), .B1(new_n383), .B2(new_n359), .ZN(new_n655));
  OAI22_X1  g469(.A1(new_n655), .A2(KEYINPUT20), .B1(new_n404), .B2(new_n365), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n383), .A2(new_n359), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n657), .A2(KEYINPUT91), .A3(new_n401), .A4(new_n364), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n362), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT33), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n446), .B2(new_n447), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n449), .A2(new_n660), .B1(new_n442), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n407), .A2(G902), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n449), .A2(new_n284), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n662), .A2(new_n663), .B1(new_n407), .B2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n659), .A2(new_n462), .A3(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n654), .A2(KEYINPUT98), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT98), .B1(new_n654), .B2(new_n666), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n519), .B2(G902), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n601), .A2(new_n534), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n649), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT34), .B(G104), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G6));
  XNOR2_X1  g489(.A(new_n384), .B(new_n401), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT99), .B1(new_n360), .B2(new_n361), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n284), .B1(new_n399), .B2(new_n353), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT99), .ZN(new_n679));
  INV_X1    g493(.A(new_n361), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n462), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n676), .A2(new_n682), .A3(new_n453), .A4(new_n683), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n684), .A2(KEYINPUT100), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(KEYINPUT100), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n654), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n685), .A2(new_n686), .A3(new_n654), .A4(KEYINPUT101), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n672), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT35), .B(G107), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G9));
  NOR2_X1   g507(.A1(new_n587), .A2(new_n588), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n584), .A2(KEYINPUT36), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n596), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n595), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n670), .A2(new_n698), .A3(new_n534), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT102), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n670), .A2(new_n698), .A3(KEYINPUT102), .A4(new_n534), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n464), .A2(new_n649), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT37), .B(G110), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G12));
  INV_X1    g519(.A(G900), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n460), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n457), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n676), .A2(new_n682), .A3(new_n453), .A4(new_n708), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n595), .A2(new_n697), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n649), .A2(new_n548), .A3(new_n654), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G128), .ZN(G30));
  NOR2_X1   g527(.A1(new_n491), .A2(new_n497), .ZN(new_n714));
  AOI21_X1  g528(.A(G902), .B1(new_n714), .B2(new_n525), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n469), .B1(new_n531), .B2(new_n491), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G472), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n536), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n524), .A3(new_n535), .ZN(new_n720));
  INV_X1    g534(.A(new_n452), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n450), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n659), .A2(new_n722), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n187), .A2(new_n720), .A3(new_n710), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n708), .B(KEYINPUT39), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n649), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT40), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT40), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n649), .A2(new_n728), .A3(new_n725), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n309), .A2(new_n313), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n730), .A2(KEYINPUT38), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(KEYINPUT38), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n724), .A2(new_n727), .A3(new_n729), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G143), .ZN(G45));
  INV_X1    g549(.A(new_n665), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n406), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n708), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n737), .A2(new_n710), .A3(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n649), .A2(new_n739), .A3(new_n548), .A4(new_n654), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G146), .ZN(G48));
  NAND2_X1  g555(.A1(new_n645), .A2(new_n642), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n647), .B1(new_n742), .B2(new_n632), .ZN(new_n743));
  OAI21_X1  g557(.A(G469), .B1(new_n743), .B2(G902), .ZN(new_n744));
  INV_X1    g558(.A(new_n603), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n745), .A3(new_n648), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n548), .A3(new_n601), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n669), .A2(new_n748), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT41), .B(G113), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G15));
  AOI21_X1  g565(.A(new_n748), .B1(new_n689), .B2(new_n690), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n201), .ZN(G18));
  NOR4_X1   g567(.A1(new_n710), .A2(new_n406), .A3(new_n462), .A4(new_n453), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n747), .A2(new_n754), .A3(new_n548), .A4(new_n654), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G119), .ZN(G21));
  NAND2_X1  g570(.A1(new_n653), .A2(new_n313), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n187), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n746), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n544), .A2(new_n525), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n513), .A2(new_n518), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n521), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT103), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n670), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(KEYINPUT103), .B(G472), .C1(new_n519), .C2(G902), .ZN(new_n765));
  AOI211_X1 g579(.A(new_n600), .B(new_n762), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n406), .A2(KEYINPUT104), .A3(new_n453), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT104), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n659), .B2(new_n722), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n770), .A2(new_n462), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n759), .A2(new_n766), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G122), .ZN(G24));
  AOI211_X1 g587(.A(new_n762), .B(new_n710), .C1(new_n764), .C2(new_n765), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n737), .A2(new_n738), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n759), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(KEYINPUT105), .B(G125), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(G27));
  INV_X1    g592(.A(KEYINPUT106), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n639), .A2(new_n630), .A3(new_n617), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n635), .A2(new_n494), .A3(new_n638), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n642), .B2(new_n645), .ZN(new_n782));
  OAI211_X1 g596(.A(G469), .B(new_n780), .C1(new_n782), .C2(new_n630), .ZN(new_n783));
  INV_X1    g597(.A(new_n605), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n630), .B(new_n617), .C1(new_n624), .C2(new_n625), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n480), .B1(new_n614), .B2(new_n616), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n629), .B1(new_n781), .B2(new_n787), .ZN(new_n788));
  AOI211_X1 g602(.A(G469), .B(G902), .C1(new_n786), .C2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n779), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n648), .A2(KEYINPUT106), .A3(new_n783), .A4(new_n784), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n547), .A2(new_n536), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT69), .B1(new_n534), .B2(new_n465), .ZN(new_n794));
  AOI211_X1 g608(.A(new_n523), .B(KEYINPUT32), .C1(new_n533), .C2(new_n520), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n600), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n730), .A2(new_n603), .A3(new_n188), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n737), .A2(KEYINPUT42), .A3(new_n738), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n792), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n790), .A3(new_n791), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n547), .A2(new_n536), .ZN(new_n802));
  INV_X1    g616(.A(new_n522), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n775), .B(new_n601), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT42), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n800), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n330), .ZN(G33));
  INV_X1    g621(.A(new_n709), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n792), .A2(new_n797), .A3(new_n808), .A4(new_n798), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G134), .ZN(G36));
  OAI21_X1  g624(.A(new_n780), .B1(new_n782), .B2(new_n630), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT45), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n604), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n640), .A2(KEYINPUT45), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n605), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT46), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n648), .B1(new_n815), .B2(KEYINPUT46), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n745), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n725), .ZN(new_n821));
  INV_X1    g635(.A(new_n730), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n187), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT110), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT43), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n406), .B2(new_n665), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT107), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n406), .A2(KEYINPUT108), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT108), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n659), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n829), .A2(new_n831), .A3(KEYINPUT43), .A4(new_n736), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n827), .A2(KEYINPUT107), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n828), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n834), .A2(KEYINPUT109), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n710), .B1(new_n534), .B2(new_n670), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n834), .B2(KEYINPUT109), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT44), .ZN(new_n838));
  OR3_X1    g652(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n838), .B1(new_n835), .B2(new_n837), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n825), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G137), .ZN(G39));
  XNOR2_X1  g656(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n843));
  INV_X1    g657(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n819), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n813), .A2(new_n814), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n784), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT46), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n648), .A3(new_n816), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n843), .B1(new_n850), .B2(new_n745), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n845), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n823), .ZN(new_n853));
  INV_X1    g667(.A(new_n548), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n600), .A4(new_n775), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT112), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(G140), .ZN(G42));
  NAND2_X1  g672(.A1(new_n744), .A2(new_n648), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(KEYINPUT49), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT113), .Z(new_n861));
  NAND3_X1  g675(.A1(new_n829), .A2(new_n736), .A3(new_n831), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n603), .A2(new_n188), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n601), .A2(new_n863), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n862), .B(new_n864), .C1(KEYINPUT49), .C2(new_n859), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n733), .A2(new_n720), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n861), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n822), .A2(new_n863), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n744), .A2(new_n648), .A3(new_n458), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n600), .B1(new_n793), .B2(new_n522), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n834), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XOR2_X1   g686(.A(KEYINPUT120), .B(KEYINPUT48), .Z(new_n873));
  XNOR2_X1  g687(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n764), .A2(new_n765), .ZN(new_n875));
  INV_X1    g689(.A(new_n762), .ZN(new_n876));
  AND4_X1   g690(.A1(new_n601), .A2(new_n875), .A3(new_n458), .A4(new_n876), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n877), .A2(new_n834), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n759), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n720), .A2(new_n600), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n870), .A2(new_n880), .A3(new_n406), .A4(new_n736), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n874), .A2(new_n455), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n747), .A2(new_n731), .A3(new_n188), .A4(new_n732), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT50), .B1(new_n878), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n877), .A2(new_n834), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT50), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n886), .A2(new_n887), .A3(new_n883), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n870), .A2(new_n880), .A3(new_n659), .A4(new_n665), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n834), .A2(new_n870), .A3(new_n774), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(KEYINPUT51), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n889), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n744), .A2(new_n603), .A3(new_n648), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n845), .B2(new_n851), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n824), .A2(new_n886), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n882), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n892), .B(new_n891), .C1(new_n885), .C2(new_n888), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT118), .B1(new_n845), .B2(new_n851), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n819), .A2(new_n844), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n850), .A2(new_n745), .A3(new_n843), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n903), .A2(new_n907), .A3(new_n897), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n902), .B1(new_n908), .B2(new_n899), .ZN(new_n909));
  XOR2_X1   g723(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n910));
  OAI21_X1  g724(.A(new_n901), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n901), .B(KEYINPUT121), .C1(new_n909), .C2(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n648), .A2(new_n784), .A3(new_n783), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n916), .A2(new_n314), .A3(new_n745), .A4(new_n463), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n548), .A2(new_n601), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n701), .A2(new_n702), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n667), .A2(new_n668), .ZN(new_n921));
  INV_X1    g735(.A(new_n748), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n659), .A2(new_n453), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n462), .B1(new_n737), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n671), .A2(new_n649), .A3(new_n314), .A4(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n772), .A2(new_n755), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n689), .A2(new_n690), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n922), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n923), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n875), .A2(new_n775), .A3(new_n698), .A4(new_n876), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n790), .A2(new_n791), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT114), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n404), .A2(KEYINPUT20), .A3(new_n365), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n401), .B1(new_n657), .B2(new_n364), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n677), .B(new_n681), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n451), .A2(new_n452), .A3(new_n708), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n721), .A2(new_n450), .A3(new_n738), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(KEYINPUT114), .A3(new_n682), .A4(new_n676), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n941), .A2(new_n916), .A3(new_n698), .ZN(new_n942));
  OAI22_X1  g756(.A1(new_n931), .A2(new_n932), .B1(new_n854), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n798), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(new_n805), .A3(new_n800), .A4(new_n809), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n930), .A2(new_n945), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n916), .A2(new_n654), .A3(new_n745), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n947), .B(new_n548), .C1(new_n711), .C2(new_n739), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n710), .A2(new_n745), .A3(new_n708), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n949), .B1(new_n796), .B2(new_n719), .ZN(new_n950));
  AND4_X1   g764(.A1(new_n187), .A2(new_n757), .A3(new_n767), .A4(new_n769), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n950), .A2(new_n790), .A3(new_n791), .A4(new_n951), .ZN(new_n952));
  AND4_X1   g766(.A1(KEYINPUT52), .A2(new_n948), .A3(new_n952), .A4(new_n776), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT52), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n747), .A2(new_n654), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n740), .B(new_n712), .C1(new_n955), .C2(new_n931), .ZN(new_n956));
  INV_X1    g770(.A(new_n951), .ZN(new_n957));
  INV_X1    g771(.A(new_n949), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n720), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n957), .A2(new_n959), .A3(new_n932), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n954), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n953), .B1(KEYINPUT115), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n956), .ZN(new_n963));
  AND4_X1   g777(.A1(KEYINPUT115), .A2(new_n963), .A3(KEYINPUT52), .A4(new_n952), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n946), .B(KEYINPUT53), .C1(new_n962), .C2(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n948), .A2(new_n952), .A3(new_n776), .A4(KEYINPUT52), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n961), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n800), .A2(new_n809), .A3(new_n805), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n792), .A2(new_n775), .A3(new_n774), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n854), .A2(new_n942), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n868), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n703), .B(new_n650), .C1(new_n669), .C2(new_n748), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n772), .A2(new_n755), .A3(new_n926), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n973), .A2(new_n752), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n967), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT53), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT54), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n965), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n976), .A2(new_n977), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n946), .B1(new_n962), .B2(new_n964), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(KEYINPUT116), .B(new_n980), .C1(new_n983), .C2(new_n979), .ZN(new_n984));
  OR3_X1    g798(.A1(new_n983), .A2(KEYINPUT116), .A3(new_n979), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n915), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g800(.A1(G952), .A2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n867), .B1(new_n986), .B2(new_n987), .ZN(G75));
  NAND2_X1  g802(.A1(new_n454), .A2(G953), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT122), .Z(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n257), .A2(new_n259), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(new_n282), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT55), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n284), .B1(new_n965), .B2(new_n978), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(G210), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT56), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n190), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n994), .A2(new_n997), .ZN(new_n1000));
  AOI211_X1 g814(.A(new_n991), .B(new_n998), .C1(new_n999), .C2(new_n1000), .ZN(G51));
  INV_X1    g815(.A(KEYINPUT123), .ZN(new_n1002));
  AOI211_X1 g816(.A(new_n284), .B(new_n846), .C1(new_n965), .C2(new_n978), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n605), .B(KEYINPUT57), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n965), .A2(new_n978), .A3(new_n979), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n979), .B1(new_n965), .B2(new_n978), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n743), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1003), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1002), .B1(new_n1009), .B2(new_n991), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n965), .A2(new_n978), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(KEYINPUT54), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n980), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n743), .B1(new_n1013), .B2(new_n1004), .ZN(new_n1014));
  OAI211_X1 g828(.A(KEYINPUT123), .B(new_n990), .C1(new_n1014), .C2(new_n1003), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1010), .A2(new_n1015), .ZN(G54));
  NAND3_X1  g830(.A1(new_n995), .A2(KEYINPUT58), .A3(G475), .ZN(new_n1017));
  OR2_X1    g831(.A1(new_n1017), .A2(new_n657), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n657), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n991), .B1(new_n1018), .B2(new_n1019), .ZN(G60));
  NAND2_X1  g834(.A1(G478), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT59), .Z(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1013), .A2(new_n662), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n990), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n985), .A2(new_n984), .A3(new_n1023), .ZN(new_n1026));
  INV_X1    g840(.A(new_n662), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(G63));
  NAND2_X1  g842(.A1(G217), .A2(G902), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT60), .Z(new_n1030));
  NAND2_X1  g844(.A1(new_n1011), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n583), .A2(new_n589), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(new_n696), .ZN(new_n1034));
  OAI211_X1 g848(.A(new_n1033), .B(new_n990), .C1(new_n1034), .C2(new_n1031), .ZN(new_n1035));
  INV_X1    g849(.A(KEYINPUT61), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1035), .B(new_n1036), .ZN(G66));
  OAI21_X1  g851(.A(G953), .B1(new_n461), .B2(new_n280), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1038), .B1(new_n975), .B2(G953), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n992), .B1(G898), .B2(new_n327), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1039), .B(new_n1040), .ZN(G69));
  NAND2_X1  g855(.A1(new_n737), .A2(new_n924), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n853), .A2(new_n1042), .ZN(new_n1043));
  NOR3_X1   g857(.A1(new_n1043), .A2(new_n918), .A3(new_n726), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n963), .A2(new_n734), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT62), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n963), .A2(KEYINPUT62), .A3(new_n734), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g864(.A1(new_n841), .A2(new_n857), .A3(new_n1045), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1051), .A2(new_n327), .ZN(new_n1052));
  XOR2_X1   g866(.A(new_n516), .B(new_n392), .Z(new_n1053));
  AOI21_X1  g867(.A(KEYINPUT124), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g868(.A(KEYINPUT124), .ZN(new_n1055));
  INV_X1    g869(.A(new_n1053), .ZN(new_n1056));
  AOI211_X1 g870(.A(new_n1055), .B(new_n1056), .C1(new_n1051), .C2(new_n327), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(KEYINPUT125), .ZN(new_n1059));
  AOI22_X1  g873(.A1(new_n852), .A2(new_n856), .B1(new_n1059), .B2(new_n968), .ZN(new_n1060));
  NAND4_X1  g874(.A1(new_n820), .A2(new_n725), .A3(new_n871), .A4(new_n951), .ZN(new_n1061));
  AND2_X1   g875(.A1(new_n1061), .A2(new_n963), .ZN(new_n1062));
  OR2_X1    g876(.A1(new_n968), .A2(new_n1059), .ZN(new_n1063));
  AND4_X1   g877(.A1(new_n841), .A2(new_n1060), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n1064), .A2(new_n327), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n1053), .B1(G900), .B2(G953), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n327), .B1(G227), .B2(G900), .ZN(new_n1068));
  INV_X1    g882(.A(new_n1068), .ZN(new_n1069));
  OAI211_X1 g883(.A(new_n1058), .B(new_n1067), .C1(KEYINPUT126), .C2(new_n1069), .ZN(new_n1070));
  AND2_X1   g884(.A1(new_n1050), .A2(new_n857), .ZN(new_n1071));
  AND2_X1   g885(.A1(new_n839), .A2(new_n840), .ZN(new_n1072));
  AOI21_X1  g886(.A(new_n1044), .B1(new_n1072), .B2(new_n825), .ZN(new_n1073));
  AOI21_X1  g887(.A(G953), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g888(.A(new_n1055), .B1(new_n1074), .B2(new_n1056), .ZN(new_n1075));
  NAND3_X1  g889(.A1(new_n1052), .A2(KEYINPUT124), .A3(new_n1053), .ZN(new_n1076));
  NAND3_X1  g890(.A1(new_n1075), .A2(new_n1067), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g891(.A1(new_n1075), .A2(KEYINPUT126), .A3(new_n1076), .ZN(new_n1078));
  NAND3_X1  g892(.A1(new_n1077), .A2(new_n1078), .A3(new_n1068), .ZN(new_n1079));
  NAND2_X1  g893(.A1(new_n1070), .A2(new_n1079), .ZN(G72));
  NAND2_X1  g894(.A1(G472), .A2(G902), .ZN(new_n1081));
  XOR2_X1   g895(.A(new_n1081), .B(KEYINPUT63), .Z(new_n1082));
  OAI21_X1  g896(.A(new_n1082), .B1(new_n1051), .B2(new_n930), .ZN(new_n1083));
  INV_X1    g897(.A(new_n716), .ZN(new_n1084));
  NAND2_X1  g898(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g899(.A(new_n539), .ZN(new_n1086));
  NAND3_X1  g900(.A1(new_n1086), .A2(new_n716), .A3(new_n1082), .ZN(new_n1087));
  OAI21_X1  g901(.A(new_n1085), .B1(new_n983), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g902(.A(KEYINPUT127), .ZN(new_n1089));
  NAND2_X1  g903(.A1(new_n1064), .A2(new_n975), .ZN(new_n1090));
  AND2_X1   g904(.A1(new_n1090), .A2(new_n1082), .ZN(new_n1091));
  OAI211_X1 g905(.A(new_n1089), .B(new_n990), .C1(new_n1091), .C2(new_n1086), .ZN(new_n1092));
  AOI21_X1  g906(.A(new_n1086), .B1(new_n1090), .B2(new_n1082), .ZN(new_n1093));
  OAI21_X1  g907(.A(KEYINPUT127), .B1(new_n1093), .B2(new_n991), .ZN(new_n1094));
  AOI21_X1  g908(.A(new_n1088), .B1(new_n1092), .B2(new_n1094), .ZN(G57));
endmodule


