//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n791, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908;
  XNOR2_X1  g000(.A(KEYINPUT80), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(G78gat), .B(G106gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT31), .B(G50gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G211gat), .B(G218gat), .Z(new_n208));
  OR2_X1    g007(.A1(G197gat), .A2(G204gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G197gat), .A2(G204gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n208), .A2(KEYINPUT71), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT69), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(G211gat), .ZN(new_n213));
  INV_X1    g012(.A(G211gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(KEYINPUT69), .ZN(new_n215));
  OAI21_X1  g014(.A(G218gat), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT70), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G218gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(KEYINPUT69), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n212), .A2(G211gat), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT70), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT22), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n211), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n208), .A2(KEYINPUT71), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI221_X1 g026(.A(new_n211), .B1(KEYINPUT71), .B2(new_n208), .C1(new_n218), .C2(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(G155gat), .A2(G162gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G141gat), .B(G148gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT2), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(G155gat), .B2(G162gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n232), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G141gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G148gat), .ZN(new_n238));
  INV_X1    g037(.A(G148gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G141gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G155gat), .B(G162gat), .ZN(new_n242));
  INV_X1    g041(.A(G155gat), .ZN(new_n243));
  INV_X1    g042(.A(G162gat), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT2), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n241), .A2(new_n242), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n236), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(KEYINPUT74), .B(KEYINPUT3), .Z(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n229), .B1(KEYINPUT29), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(G228gat), .A3(G233gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT29), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n227), .A2(new_n228), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT78), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n227), .A2(new_n228), .A3(new_n254), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT3), .B1(new_n258), .B2(KEYINPUT78), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n248), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n253), .B1(new_n260), .B2(KEYINPUT79), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(new_n255), .B2(new_n256), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n258), .A2(KEYINPUT78), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n247), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT79), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n249), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n247), .B1(new_n255), .B2(new_n269), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n270), .A2(new_n252), .B1(G228gat), .B2(G233gat), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n207), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  AOI211_X1 g072(.A(new_n271), .B(new_n206), .C1(new_n261), .C2(new_n267), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n203), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT27), .B(G183gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n276), .B(KEYINPUT64), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT28), .B1(new_n277), .B2(G190gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT28), .ZN(new_n279));
  INV_X1    g078(.A(G190gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n276), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT65), .ZN(new_n285));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NOR3_X1   g086(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n284), .A2(KEYINPUT65), .A3(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n278), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n283), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n293), .A2(new_n294), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n286), .ZN(new_n297));
  NAND3_X1  g096(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n295), .A2(new_n299), .A3(KEYINPUT25), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n291), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G134gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G127gat), .ZN(new_n307));
  INV_X1    g106(.A(G127gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G134gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT1), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G120gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G113gat), .ZN(new_n313));
  INV_X1    g112(.A(G113gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT67), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G113gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n317), .A3(G120gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n311), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(G120gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT1), .B1(new_n321), .B2(KEYINPUT66), .ZN(new_n322));
  XNOR2_X1  g121(.A(G113gat), .B(G120gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT66), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n307), .A2(new_n309), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n319), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n305), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G227gat), .ZN(new_n330));
  INV_X1    g129(.A(G233gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n278), .A2(new_n290), .B1(new_n302), .B2(new_n303), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n310), .B1(new_n323), .B2(new_n324), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n313), .A2(new_n320), .A3(new_n324), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n327), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n313), .ZN(new_n337));
  INV_X1    g136(.A(new_n327), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n310), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n329), .A2(new_n332), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT32), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT68), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT68), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n345), .A3(KEYINPUT32), .ZN(new_n346));
  XNOR2_X1  g145(.A(G15gat), .B(G43gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(G71gat), .B(G99gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT33), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n349), .B1(new_n342), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n344), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n342), .B(KEYINPUT32), .C1(new_n350), .C2(new_n349), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n332), .B1(new_n329), .B2(new_n341), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT34), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n352), .B2(new_n353), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(KEYINPUT79), .B(new_n247), .C1(new_n263), .C2(new_n264), .ZN(new_n360));
  INV_X1    g159(.A(new_n253), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n260), .A2(KEYINPUT79), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n272), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(new_n206), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n268), .A2(new_n272), .A3(new_n207), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n202), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n275), .A2(new_n359), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369));
  XNOR2_X1  g168(.A(G1gat), .B(G29gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT0), .ZN(new_n371));
  XNOR2_X1  g170(.A(G57gat), .B(G85gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n371), .B(new_n372), .Z(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n247), .A2(KEYINPUT3), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n250), .A2(new_n340), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n378), .B1(new_n328), .B2(new_n248), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n338), .B1(new_n322), .B2(new_n325), .ZN(new_n380));
  NOR4_X1   g179(.A1(new_n380), .A2(new_n247), .A3(new_n319), .A4(KEYINPUT4), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n375), .B(new_n377), .C1(new_n379), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT75), .ZN(new_n383));
  INV_X1    g182(.A(new_n375), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n380), .A2(new_n247), .A3(new_n319), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n336), .A2(new_n339), .B1(new_n236), .B2(new_n246), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT5), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n383), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n388), .A2(new_n382), .A3(KEYINPUT75), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n374), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT76), .B1(new_n392), .B2(KEYINPUT6), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n388), .A2(new_n382), .A3(KEYINPUT75), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n388), .B1(KEYINPUT75), .B2(new_n382), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n373), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n390), .A2(new_n391), .A3(new_n374), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n393), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n398), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n229), .ZN(new_n405));
  INV_X1    g204(.A(G226gat), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(new_n331), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n408), .B1(new_n333), .B2(KEYINPUT29), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT73), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n305), .B2(new_n407), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n333), .A2(KEYINPUT73), .A3(new_n408), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n405), .B(new_n409), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT72), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n305), .A2(new_n414), .A3(new_n407), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n407), .B1(new_n305), .B2(new_n254), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT72), .B1(new_n333), .B2(new_n408), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n229), .B(new_n415), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G8gat), .B(G36gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420));
  XOR2_X1   g219(.A(new_n419), .B(new_n420), .Z(new_n421));
  NAND3_X1  g220(.A1(new_n413), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT30), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n413), .A2(new_n418), .ZN(new_n425));
  INV_X1    g224(.A(new_n421), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n413), .A2(new_n418), .A3(KEYINPUT30), .A4(new_n421), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n369), .B1(new_n404), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n431));
  AOI211_X1 g230(.A(KEYINPUT77), .B(new_n431), .C1(new_n401), .C2(new_n403), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n368), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT35), .ZN(new_n434));
  OAI21_X1  g233(.A(KEYINPUT85), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT85), .ZN(new_n436));
  INV_X1    g235(.A(new_n400), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n396), .A2(new_n398), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n437), .B1(new_n438), .B2(KEYINPUT76), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n402), .B1(new_n439), .B2(new_n399), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT77), .B1(new_n440), .B2(new_n431), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n404), .A2(new_n369), .A3(new_n429), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n436), .B(KEYINPUT35), .C1(new_n443), .C2(new_n368), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n403), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n434), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n368), .A2(new_n431), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n435), .A2(new_n444), .A3(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n359), .B(KEYINPUT36), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n377), .B1(new_n379), .B2(new_n381), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n384), .ZN(new_n453));
  OR2_X1    g252(.A1(new_n385), .A2(new_n386), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n453), .B(KEYINPUT39), .C1(new_n384), .C2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(KEYINPUT81), .B(KEYINPUT39), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n452), .A2(new_n384), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n457), .A2(new_n458), .A3(new_n373), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n457), .B2(new_n373), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n455), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(KEYINPUT40), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n400), .A3(new_n431), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT37), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n427), .B1(new_n464), .B2(new_n421), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT73), .B1(new_n333), .B2(new_n408), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n305), .A2(new_n410), .A3(new_n407), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n416), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT83), .B1(new_n468), .B2(new_n405), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n229), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(new_n405), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n469), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n465), .B1(new_n475), .B2(new_n464), .ZN(new_n476));
  XOR2_X1   g275(.A(KEYINPUT84), .B(KEYINPUT38), .Z(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(new_n425), .B2(KEYINPUT37), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n476), .A2(new_n477), .B1(new_n465), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n403), .A2(new_n445), .A3(new_n422), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n463), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n275), .A2(new_n367), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n451), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n275), .A2(new_n367), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n441), .B2(new_n442), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n450), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G29gat), .A2(G36gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n488), .B(KEYINPUT88), .Z(new_n489));
  NOR2_X1   g288(.A1(G29gat), .A2(G36gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(KEYINPUT14), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G43gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(G50gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT90), .B(G50gat), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(new_n493), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT89), .B(KEYINPUT15), .Z(new_n497));
  OAI21_X1  g296(.A(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n494), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n493), .A2(G50gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(KEYINPUT15), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  OR3_X1    g301(.A1(new_n489), .A2(new_n491), .A3(new_n501), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT17), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(KEYINPUT92), .A3(KEYINPUT17), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT16), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(G1gat), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(G1gat), .B2(new_n510), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(G8gat), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT91), .B1(new_n504), .B2(KEYINPUT17), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT17), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n502), .A2(new_n516), .A3(new_n517), .A4(new_n503), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n514), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n509), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n504), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n514), .ZN(new_n522));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT18), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT87), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(G113gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(new_n237), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n529), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT12), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n520), .A2(KEYINPUT18), .A3(new_n522), .A4(new_n523), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n504), .B(new_n514), .Z(new_n536));
  XOR2_X1   g335(.A(new_n523), .B(KEYINPUT13), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(KEYINPUT93), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n535), .A2(new_n543), .A3(new_n538), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n526), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT94), .ZN(new_n546));
  INV_X1    g345(.A(new_n533), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n541), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT95), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n554), .B2(new_n553), .ZN(new_n556));
  XNOR2_X1  g355(.A(G71gat), .B(G78gat), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(new_n552), .ZN(new_n559));
  INV_X1    g358(.A(G57gat), .ZN(new_n560));
  INV_X1    g359(.A(G64gat), .ZN(new_n561));
  OR3_X1    g360(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT96), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n560), .B2(KEYINPUT96), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g363(.A1(new_n556), .A2(new_n558), .B1(new_n559), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n565), .A2(KEYINPUT21), .ZN(new_n566));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G127gat), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n514), .B1(new_n565), .B2(KEYINPUT21), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n569), .A2(new_n570), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(new_n243), .ZN(new_n575));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  OR2_X1    g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n571), .A2(new_n572), .A3(new_n577), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n515), .A2(new_n518), .ZN(new_n581));
  XOR2_X1   g380(.A(G99gat), .B(G106gat), .Z(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT98), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n584));
  NAND2_X1  g383(.A1(G85gat), .A2(G92gat), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n585), .ZN(new_n587));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  AOI22_X1  g389(.A1(KEYINPUT8), .A2(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(new_n587), .A3(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n583), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n583), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n509), .A2(new_n581), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n595), .ZN(new_n597));
  AND2_X1   g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n521), .A2(new_n597), .B1(KEYINPUT41), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G190gat), .B(G218gat), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n600), .B(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n604));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n603), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n580), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n592), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n609), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(new_n583), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT100), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(new_n565), .A3(new_n593), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n597), .A2(new_n565), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT101), .Z(new_n620));
  XOR2_X1   g419(.A(G120gat), .B(G148gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT102), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(KEYINPUT103), .ZN(new_n623));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT10), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n614), .A2(new_n627), .A3(new_n615), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n565), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n617), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n620), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n619), .B(KEYINPUT101), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n618), .B1(new_n628), .B2(new_n629), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n625), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n608), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n487), .A2(new_n551), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n404), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g439(.A1(new_n638), .A2(new_n429), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT16), .B(G8gat), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT104), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT42), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n642), .A2(G8gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT105), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(G1325gat));
  OAI21_X1  g447(.A(G15gat), .B1(new_n638), .B2(new_n451), .ZN(new_n649));
  INV_X1    g448(.A(new_n359), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n650), .A2(G15gat), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n649), .B1(new_n638), .B2(new_n651), .ZN(G1326gat));
  NOR2_X1   g451(.A1(new_n638), .A2(new_n484), .ZN(new_n653));
  XOR2_X1   g452(.A(KEYINPUT43), .B(G22gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(G1327gat));
  AOI21_X1  g454(.A(new_n607), .B1(new_n450), .B2(new_n486), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n545), .A2(new_n547), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT94), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n540), .B1(new_n658), .B2(new_n548), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n659), .A2(new_n580), .A3(new_n636), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n662), .A2(G29gat), .A3(new_n404), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n483), .A2(new_n485), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT35), .B1(new_n443), .B2(new_n368), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n448), .B1(new_n668), .B2(KEYINPUT85), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n667), .B1(new_n669), .B2(new_n444), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n666), .B1(new_n670), .B2(new_n607), .ZN(new_n671));
  INV_X1    g470(.A(new_n607), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n487), .A2(KEYINPUT44), .A3(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n674), .A2(new_n660), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G29gat), .B1(new_n676), .B2(new_n404), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n665), .A2(new_n677), .ZN(G1328gat));
  NOR3_X1   g477(.A1(new_n662), .A2(G36gat), .A3(new_n429), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT46), .ZN(new_n680));
  OAI21_X1  g479(.A(G36gat), .B1(new_n676), .B2(new_n429), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(G1329gat));
  OAI21_X1  g481(.A(new_n493), .B1(new_n662), .B2(new_n650), .ZN(new_n683));
  INV_X1    g482(.A(new_n451), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(G43gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n676), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g486(.A(new_n495), .B1(new_n661), .B2(new_n482), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n689), .B2(KEYINPUT48), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n482), .A2(new_n495), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n676), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n689), .A2(KEYINPUT48), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n692), .B(new_n693), .Z(G1331gat));
  INV_X1    g493(.A(new_n636), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n551), .A2(new_n695), .A3(new_n608), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n487), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n404), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(new_n560), .ZN(G1332gat));
  NOR2_X1   g498(.A1(new_n697), .A2(new_n429), .ZN(new_n700));
  NOR2_X1   g499(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n701));
  AND2_X1   g500(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n700), .B2(new_n701), .ZN(G1333gat));
  NOR3_X1   g503(.A1(new_n697), .A2(G71gat), .A3(new_n650), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n487), .A2(new_n684), .A3(new_n696), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(G71gat), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1334gat));
  NOR2_X1   g508(.A1(new_n697), .A2(new_n484), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT109), .B(G78gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1335gat));
  NOR3_X1   g511(.A1(new_n551), .A2(new_n580), .A3(new_n695), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n674), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G85gat), .B1(new_n714), .B2(new_n404), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n551), .A2(new_n580), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n656), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT51), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n636), .A2(new_n589), .A3(new_n440), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n715), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT110), .ZN(G1336gat));
  OAI21_X1  g520(.A(G92gat), .B1(new_n714), .B2(new_n429), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT112), .B(KEYINPUT52), .Z(new_n723));
  NOR3_X1   g522(.A1(new_n695), .A2(G92gat), .A3(new_n429), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n722), .B(new_n723), .C1(new_n718), .C2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT111), .ZN(new_n728));
  AND4_X1   g527(.A1(new_n487), .A2(new_n672), .A3(new_n716), .A4(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n656), .B2(new_n716), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n724), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n722), .A2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n726), .B1(new_n732), .B2(new_n733), .ZN(G1337gat));
  OAI21_X1  g533(.A(G99gat), .B1(new_n714), .B2(new_n451), .ZN(new_n735));
  OR3_X1    g534(.A1(new_n695), .A2(G99gat), .A3(new_n650), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n718), .B2(new_n736), .ZN(G1338gat));
  NAND4_X1  g536(.A1(new_n671), .A2(new_n673), .A3(new_n482), .A4(new_n713), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G106gat), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT113), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n695), .A2(G106gat), .A3(new_n484), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n729), .B2(new_n730), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n738), .A2(new_n745), .A3(G106gat), .ZN(new_n746));
  OAI211_X1 g545(.A(KEYINPUT114), .B(new_n741), .C1(new_n729), .C2(new_n730), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n740), .A2(new_n744), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT53), .ZN(new_n749));
  XOR2_X1   g548(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n750));
  INV_X1    g549(.A(new_n741), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n739), .B(new_n750), .C1(new_n718), .C2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n749), .A2(KEYINPUT116), .A3(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1339gat));
  NAND2_X1  g556(.A1(new_n637), .A2(new_n659), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n628), .A2(new_n618), .A3(new_n629), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n631), .A2(KEYINPUT54), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n626), .B1(new_n634), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(KEYINPUT55), .A3(new_n763), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n632), .A3(new_n767), .ZN(new_n768));
  AND2_X1   g567(.A1(new_n520), .A2(new_n522), .ZN(new_n769));
  OAI22_X1  g568(.A1(new_n769), .A2(new_n523), .B1(new_n536), .B2(new_n537), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n532), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n541), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n768), .A2(new_n607), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n772), .B1(new_n635), .B2(new_n632), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n766), .A2(new_n632), .A3(new_n767), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n551), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n774), .B1(new_n777), .B2(new_n672), .ZN(new_n778));
  INV_X1    g577(.A(new_n580), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n759), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(new_n482), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n781), .A2(new_n440), .A3(new_n429), .A4(new_n359), .ZN(new_n782));
  OAI21_X1  g581(.A(G113gat), .B1(new_n782), .B2(new_n659), .ZN(new_n783));
  NOR4_X1   g582(.A1(new_n780), .A2(new_n404), .A3(new_n431), .A4(new_n368), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n784), .A2(new_n315), .A3(new_n317), .A4(new_n551), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(KEYINPUT117), .Z(G1340gat));
  NOR3_X1   g586(.A1(new_n782), .A2(new_n312), .A3(new_n695), .ZN(new_n788));
  AOI21_X1  g587(.A(G120gat), .B1(new_n784), .B2(new_n636), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(G1341gat));
  OAI21_X1  g589(.A(G127gat), .B1(new_n782), .B2(new_n779), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n784), .A2(new_n308), .A3(new_n580), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(G1342gat));
  NAND3_X1  g592(.A1(new_n784), .A2(new_n306), .A3(new_n672), .ZN(new_n794));
  OR2_X1    g593(.A1(new_n794), .A2(KEYINPUT56), .ZN(new_n795));
  OAI21_X1  g594(.A(G134gat), .B1(new_n782), .B2(new_n607), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(KEYINPUT56), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(G1343gat));
  NOR2_X1   g597(.A1(new_n780), .A2(new_n404), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n451), .A2(new_n482), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n431), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n802), .A2(G141gat), .A3(new_n659), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(KEYINPUT58), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT57), .B1(new_n780), .B2(new_n484), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n659), .A2(new_n768), .B1(new_n695), .B2(new_n772), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n773), .B1(new_n806), .B2(new_n607), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n758), .B1(new_n807), .B2(new_n580), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n808), .A2(new_n809), .A3(new_n482), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n684), .A2(new_n404), .A3(new_n431), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n805), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G141gat), .B1(new_n812), .B2(new_n659), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n804), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(KEYINPUT118), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n805), .A2(new_n810), .A3(new_n816), .A4(new_n811), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n551), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n803), .B1(new_n819), .B2(G141gat), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n814), .B1(new_n820), .B2(new_n821), .ZN(G1344gat));
  NAND3_X1  g621(.A1(new_n815), .A2(new_n636), .A3(new_n817), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n239), .A2(KEYINPUT59), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n823), .A2(KEYINPUT119), .A3(new_n824), .ZN(new_n828));
  OAI21_X1  g627(.A(G148gat), .B1(new_n812), .B2(new_n695), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT59), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n802), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n832), .A2(new_n239), .A3(new_n636), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(G1345gat));
  AOI21_X1  g633(.A(G155gat), .B1(new_n832), .B2(new_n580), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n580), .A2(G155gat), .ZN(new_n836));
  XOR2_X1   g635(.A(new_n836), .B(KEYINPUT120), .Z(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n818), .B2(new_n837), .ZN(G1346gat));
  AOI21_X1  g637(.A(G162gat), .B1(new_n832), .B2(new_n672), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n607), .A2(new_n244), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n818), .B2(new_n840), .ZN(G1347gat));
  NOR4_X1   g640(.A1(new_n780), .A2(new_n440), .A3(new_n429), .A4(new_n368), .ZN(new_n842));
  INV_X1    g641(.A(G169gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(new_n551), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n440), .A2(new_n429), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n781), .A2(new_n359), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(G169gat), .B1(new_n846), .B2(new_n659), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n844), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g652(.A(KEYINPUT122), .B(new_n844), .C1(new_n849), .C2(new_n850), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1348gat));
  OAI21_X1  g654(.A(G176gat), .B1(new_n846), .B2(new_n695), .ZN(new_n856));
  INV_X1    g655(.A(G176gat), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n857), .A3(new_n636), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(G1349gat));
  OAI21_X1  g658(.A(G183gat), .B1(new_n846), .B2(new_n779), .ZN(new_n860));
  INV_X1    g659(.A(new_n277), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n842), .A2(new_n861), .A3(new_n580), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g663(.A(G190gat), .B1(new_n846), .B2(new_n607), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT61), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n842), .A2(new_n280), .A3(new_n672), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1351gat));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n869));
  INV_X1    g668(.A(new_n810), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n809), .B1(new_n808), .B2(new_n482), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n805), .A2(new_n810), .A3(KEYINPUT124), .ZN(new_n873));
  INV_X1    g672(.A(new_n845), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n684), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n872), .A2(new_n551), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(G197gat), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n780), .A2(new_n440), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n800), .A2(new_n429), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n659), .A2(G197gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT123), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT125), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n877), .A2(new_n885), .A3(new_n882), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1352gat));
  NAND2_X1  g686(.A1(new_n878), .A2(new_n879), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n888), .A2(G204gat), .A3(new_n695), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT62), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n872), .A2(new_n636), .A3(new_n873), .A4(new_n875), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G204gat), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1353gat));
  NOR2_X1   g692(.A1(new_n870), .A2(new_n871), .ZN(new_n894));
  INV_X1    g693(.A(new_n875), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n779), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT126), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n214), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n894), .A2(KEYINPUT126), .A3(new_n896), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n899), .A2(KEYINPUT63), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT63), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n580), .A2(new_n220), .A3(new_n221), .ZN(new_n903));
  OAI22_X1  g702(.A1(new_n901), .A2(new_n902), .B1(new_n888), .B2(new_n903), .ZN(G1354gat));
  NOR3_X1   g703(.A1(new_n895), .A2(new_n219), .A3(new_n607), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n872), .A2(new_n873), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n219), .B1(new_n888), .B2(new_n607), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT127), .Z(G1355gat));
endmodule


