//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT64), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT64), .A2(G143), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n192), .B1(G143), .B2(new_n190), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n196));
  OAI21_X1  g010(.A(G128), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n193), .A2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT64), .A2(G143), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT64), .A2(G143), .ZN(new_n200));
  OAI21_X1  g014(.A(G146), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n195), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n201), .A2(new_n196), .A3(G128), .A4(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G137), .ZN(new_n209));
  INV_X1    g023(.A(G134), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(G134), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n205), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT11), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(new_n210), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n208), .A2(G137), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n206), .A2(KEYINPUT66), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n210), .A2(G137), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(KEYINPUT65), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT11), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n212), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n219), .A2(new_n205), .A3(new_n220), .A4(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n225), .A2(new_n226), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n204), .B(new_n214), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n219), .A2(new_n220), .A3(new_n224), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G131), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(new_n227), .B2(new_n228), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n189), .A2(new_n191), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n195), .B1(new_n234), .B2(G146), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT0), .A3(G128), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT0), .B(G128), .Z(new_n237));
  NAND2_X1  g051(.A1(new_n193), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n230), .B1(new_n233), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n207), .A2(new_n209), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n242), .A2(new_n216), .B1(new_n243), .B2(new_n212), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n244), .A2(KEYINPUT67), .A3(new_n205), .A4(new_n220), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n225), .A2(new_n226), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n245), .A2(new_n246), .B1(G131), .B2(new_n231), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n247), .A2(KEYINPUT70), .A3(new_n239), .ZN(new_n248));
  OAI211_X1 g062(.A(KEYINPUT30), .B(new_n229), .C1(new_n241), .C2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G119), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G116), .ZN(new_n251));
  INV_X1    g065(.A(G116), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G119), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT2), .B(G113), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(KEYINPUT69), .ZN(new_n257));
  XNOR2_X1  g071(.A(G116), .B(G119), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n256), .B1(new_n261), .B2(new_n255), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n213), .B1(new_n245), .B2(new_n246), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n233), .A2(new_n240), .B1(new_n264), .B2(new_n204), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n265), .A2(KEYINPUT68), .A3(KEYINPUT30), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n229), .B1(new_n239), .B2(new_n247), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT30), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n249), .B(new_n263), .C1(new_n266), .C2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT68), .B1(new_n265), .B2(KEYINPUT30), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n268), .A2(new_n267), .A3(new_n269), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n276), .A2(KEYINPUT71), .A3(new_n263), .A4(new_n249), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT31), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n233), .A2(new_n230), .A3(new_n240), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT70), .B1(new_n247), .B2(new_n239), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n283), .A2(new_n262), .A3(new_n229), .ZN(new_n284));
  INV_X1    g098(.A(G237), .ZN(new_n285));
  INV_X1    g099(.A(G953), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(G210), .ZN(new_n287));
  INV_X1    g101(.A(G101), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n287), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n289), .B(new_n290), .Z(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n280), .B1(new_n284), .B2(new_n292), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n281), .A2(new_n282), .B1(new_n204), .B2(new_n264), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n262), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(KEYINPUT72), .A3(new_n291), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n278), .A2(new_n279), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n294), .A2(KEYINPUT28), .A3(new_n262), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n268), .A2(new_n263), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT28), .B1(new_n265), .B2(new_n262), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n299), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n292), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n298), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(KEYINPUT73), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n273), .A2(new_n277), .B1(new_n293), .B2(new_n296), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(new_n279), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n187), .B(new_n188), .C1(new_n308), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT32), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n310), .A2(new_n279), .B1(new_n305), .B2(new_n306), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n278), .A2(new_n297), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT31), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n309), .A3(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n318), .A2(KEYINPUT32), .A3(new_n187), .A4(new_n188), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n299), .A2(new_n291), .A3(new_n300), .A4(new_n302), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT29), .B1(new_n320), .B2(new_n321), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n284), .B1(new_n273), .B2(new_n277), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n322), .B(new_n323), .C1(new_n324), .C2(new_n291), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT28), .ZN(new_n326));
  OR2_X1    g140(.A1(new_n294), .A2(new_n262), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(new_n295), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(new_n301), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n291), .A2(KEYINPUT29), .ZN(new_n330));
  AOI21_X1  g144(.A(G902), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT75), .B1(new_n332), .B2(G472), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n334));
  AOI211_X1 g148(.A(new_n334), .B(new_n187), .C1(new_n325), .C2(new_n331), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n314), .B(new_n319), .C1(new_n333), .C2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G140), .ZN(new_n337));
  INV_X1    g151(.A(G227), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(G953), .ZN(new_n339));
  XOR2_X1   g153(.A(new_n337), .B(new_n339), .Z(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G104), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G107), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n342), .A2(G107), .ZN(new_n345));
  OAI21_X1  g159(.A(G101), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT3), .B1(new_n342), .B2(G107), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n348));
  INV_X1    g162(.A(G107), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(G104), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n347), .A2(new_n350), .A3(new_n288), .A4(new_n343), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n204), .A2(KEYINPUT10), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n347), .A2(new_n350), .A3(new_n343), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G101), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT4), .A3(new_n351), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n357), .A3(G101), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n353), .B1(new_n359), .B2(new_n239), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n361));
  INV_X1    g175(.A(G128), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n203), .B1(new_n363), .B2(new_n235), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n364), .A2(KEYINPUT85), .A3(new_n352), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT85), .B1(new_n364), .B2(new_n352), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n361), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT86), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT86), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n369), .B(new_n361), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n360), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(new_n247), .ZN(new_n372));
  AOI211_X1 g186(.A(new_n233), .B(new_n360), .C1(new_n368), .C2(new_n370), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n341), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT87), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI22_X1  g190(.A1(new_n365), .A2(new_n366), .B1(new_n352), .B2(new_n204), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n233), .ZN(new_n378));
  XOR2_X1   g192(.A(new_n378), .B(KEYINPUT12), .Z(new_n379));
  INV_X1    g193(.A(new_n373), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(new_n340), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT87), .B(new_n341), .C1(new_n372), .C2(new_n373), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n376), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G469), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n188), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n384), .A2(new_n188), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n340), .B1(new_n379), .B2(new_n380), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n372), .A2(new_n373), .A3(new_n341), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n386), .B1(new_n389), .B2(G469), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT9), .B(G234), .Z(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G221), .B1(new_n393), .B2(G902), .ZN(new_n394));
  XOR2_X1   g208(.A(new_n394), .B(KEYINPUT83), .Z(new_n395));
  XOR2_X1   g209(.A(new_n395), .B(KEYINPUT84), .Z(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n391), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n263), .A2(KEYINPUT88), .A3(new_n358), .A4(new_n356), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT88), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n359), .B2(new_n262), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n257), .A2(new_n260), .A3(KEYINPUT5), .ZN(new_n403));
  OAI21_X1  g217(.A(G113), .B1(new_n251), .B2(KEYINPUT5), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n256), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(new_n352), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT89), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n256), .B1(new_n403), .B2(new_n405), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT89), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(new_n411), .A3(new_n352), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n402), .A2(new_n413), .ZN(new_n414));
  XOR2_X1   g228(.A(G110), .B(G122), .Z(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n415), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n402), .A2(new_n413), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(KEYINPUT6), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n414), .A2(new_n420), .A3(new_n415), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n239), .A2(G125), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(G125), .B2(new_n204), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT90), .B(G224), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n286), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT91), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n423), .B(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n419), .A2(new_n421), .A3(new_n427), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n410), .A2(new_n352), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n429), .A2(KEYINPUT94), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(KEYINPUT94), .ZN(new_n431));
  INV_X1    g245(.A(new_n352), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n258), .A2(KEYINPUT5), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n407), .B1(new_n433), .B2(new_n404), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT93), .ZN(new_n435));
  OAI22_X1  g249(.A1(new_n430), .A2(new_n431), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(KEYINPUT92), .B(KEYINPUT8), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n415), .B(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT7), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n426), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n423), .B(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n442), .A3(new_n418), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n428), .A2(new_n188), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G210), .B1(G237), .B2(G902), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n428), .A2(new_n443), .A3(new_n188), .A4(new_n445), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G214), .B1(G237), .B2(G902), .ZN(new_n450));
  INV_X1    g264(.A(G952), .ZN(new_n451));
  AOI211_X1 g265(.A(G953), .B(new_n451), .C1(G234), .C2(G237), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT21), .B(G898), .Z(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI211_X1 g268(.A(new_n188), .B(new_n286), .C1(G234), .C2(G237), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n452), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n449), .A2(new_n450), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n398), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT78), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n362), .A2(G119), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT23), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n362), .A2(G119), .ZN(new_n464));
  OAI211_X1 g278(.A(KEYINPUT78), .B(KEYINPUT23), .C1(new_n362), .C2(G119), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n362), .A2(KEYINPUT23), .A3(G119), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT77), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G110), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n466), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT79), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT79), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n466), .A2(new_n469), .A3(new_n473), .A4(new_n470), .ZN(new_n474));
  INV_X1    g288(.A(new_n464), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(new_n461), .ZN(new_n476));
  XOR2_X1   g290(.A(KEYINPUT24), .B(G110), .Z(new_n477));
  OAI211_X1 g291(.A(new_n472), .B(new_n474), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(G125), .B(G140), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT16), .ZN(new_n480));
  INV_X1    g294(.A(G125), .ZN(new_n481));
  OR3_X1    g295(.A1(new_n481), .A2(KEYINPUT16), .A3(G140), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(G146), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(KEYINPUT80), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n479), .A2(new_n190), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n478), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT81), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n480), .A2(new_n482), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n190), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n483), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n476), .A2(new_n477), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n466), .A2(new_n469), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n490), .B(new_n491), .C1(new_n470), .C2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n486), .A2(new_n487), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT22), .B(G137), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n286), .A2(G221), .A3(G234), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n495), .B(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n487), .B1(new_n486), .B2(new_n493), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n494), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n500), .B1(new_n503), .B2(new_n497), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT82), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT25), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n504), .A2(new_n188), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G234), .ZN(new_n511));
  OAI21_X1  g325(.A(G217), .B1(new_n511), .B2(G902), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT76), .ZN(new_n513));
  INV_X1    g327(.A(new_n494), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n497), .B1(new_n514), .B2(new_n501), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n515), .A2(new_n188), .A3(new_n509), .A4(new_n499), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n507), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n510), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n512), .A2(new_n188), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n504), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n234), .A2(G128), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT13), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n194), .A2(G128), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n234), .B2(G128), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n525), .B(KEYINPUT97), .C1(new_n524), .C2(new_n527), .ZN(new_n528));
  OR3_X1    g342(.A1(new_n523), .A2(KEYINPUT97), .A3(new_n524), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(G134), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G122), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G116), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(KEYINPUT96), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(G116), .B2(new_n531), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n534), .A2(new_n349), .B1(new_n210), .B2(new_n527), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n530), .B(new_n535), .C1(new_n349), .C2(new_n534), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n349), .B1(new_n533), .B2(KEYINPUT14), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n537), .A2(new_n534), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n527), .B(new_n210), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n534), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n392), .A2(G217), .A3(new_n286), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n543), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n536), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT98), .ZN(new_n548));
  INV_X1    g362(.A(G478), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(KEYINPUT15), .ZN(new_n550));
  XOR2_X1   g364(.A(new_n548), .B(new_n550), .Z(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n490), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n285), .A2(new_n286), .A3(G214), .ZN(new_n554));
  OR2_X1    g368(.A1(new_n554), .A2(G143), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n189), .A3(new_n191), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(new_n205), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT17), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n555), .A2(new_n556), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G131), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n557), .A2(new_n205), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n553), .B(new_n559), .C1(new_n563), .C2(KEYINPUT17), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n560), .A2(KEYINPUT18), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n558), .A2(KEYINPUT18), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n479), .B(new_n190), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n565), .A2(new_n566), .A3(new_n567), .A4(new_n562), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(G113), .B(G122), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(new_n342), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n563), .A2(KEYINPUT95), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n479), .B(KEYINPUT19), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n190), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n561), .A2(new_n577), .A3(new_n562), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n574), .A2(new_n484), .A3(new_n576), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n571), .B1(new_n579), .B2(new_n568), .ZN(new_n580));
  OR2_X1    g394(.A1(new_n573), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT20), .ZN(new_n582));
  INV_X1    g396(.A(G475), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n188), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n583), .B(new_n188), .C1(new_n573), .C2(new_n580), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT20), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n569), .B(new_n571), .ZN(new_n588));
  OAI21_X1  g402(.A(G475), .B1(new_n588), .B2(G902), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n552), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n336), .A2(new_n459), .A3(new_n522), .A4(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  OAI21_X1  g407(.A(new_n188), .B1(new_n308), .B2(new_n311), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(G472), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n312), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n396), .B1(new_n385), .B2(new_n390), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(new_n598), .A3(new_n522), .ZN(new_n599));
  INV_X1    g413(.A(new_n450), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n447), .B2(new_n448), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT99), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n536), .A2(new_n541), .A3(new_n545), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n545), .B1(new_n536), .B2(new_n541), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n544), .A2(KEYINPUT33), .A3(new_n546), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n607), .A3(new_n188), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(G478), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT100), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n547), .A2(new_n549), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n610), .B1(new_n609), .B2(new_n611), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n590), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n602), .A2(new_n456), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n599), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT34), .B(G104), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  INV_X1    g434(.A(new_n590), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n552), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n602), .A2(new_n456), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n599), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT35), .B(G107), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  INV_X1    g441(.A(new_n458), .ZN(new_n628));
  INV_X1    g442(.A(new_n591), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n486), .A2(new_n493), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n498), .A2(KEYINPUT36), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT101), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n630), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n520), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n518), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n635), .A2(KEYINPUT102), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(KEYINPUT102), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n629), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n597), .A2(new_n628), .A3(new_n638), .A4(new_n598), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  AOI21_X1  g455(.A(new_n398), .B1(new_n637), .B2(new_n636), .ZN(new_n642));
  AOI21_X1  g456(.A(KEYINPUT99), .B1(new_n449), .B2(new_n450), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n644));
  AOI211_X1 g458(.A(new_n644), .B(new_n600), .C1(new_n447), .C2(new_n448), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(G900), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n455), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n452), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n622), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n336), .A2(new_n642), .A3(new_n646), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  XNOR2_X1  g468(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n650), .B(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT40), .B1(new_n398), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n635), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT40), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n598), .A2(new_n660), .A3(new_n656), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n658), .A2(new_n450), .A3(new_n659), .A4(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n291), .B1(new_n327), .B2(new_n295), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n188), .B1(new_n310), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(G472), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n314), .A2(new_n319), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n621), .A2(new_n551), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n449), .B(KEYINPUT38), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n670));
  OR3_X1    g484(.A1(new_n662), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n670), .B1(new_n662), .B2(new_n669), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n234), .ZN(G45));
  NOR2_X1   g488(.A1(new_n615), .A2(new_n651), .ZN(new_n675));
  AND2_X1   g489(.A1(new_n675), .A2(new_n646), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n336), .A2(new_n676), .A3(new_n642), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  NAND2_X1  g492(.A1(new_n383), .A2(new_n188), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n384), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n395), .ZN(new_n683));
  INV_X1    g497(.A(new_n681), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n383), .A2(new_n188), .A3(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n616), .A2(new_n336), .A3(new_n522), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT41), .B(G113), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G15));
  NAND4_X1  g504(.A1(new_n623), .A2(new_n336), .A3(new_n522), .A4(new_n687), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G116), .ZN(G18));
  NOR3_X1   g506(.A1(new_n602), .A2(new_n686), .A3(new_n456), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n336), .A3(new_n638), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  OAI21_X1  g509(.A(new_n292), .B1(new_n328), .B2(new_n301), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n298), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n310), .A2(new_n279), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n187), .B(new_n188), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n595), .A2(new_n522), .A3(new_n667), .A4(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT106), .B1(new_n701), .B2(new_n693), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n383), .A2(new_n188), .A3(new_n684), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n684), .B1(new_n383), .B2(new_n188), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n646), .A2(new_n705), .A3(new_n457), .A4(new_n683), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT106), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n700), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n531), .ZN(G24));
  AOI22_X1  g524(.A1(new_n316), .A2(KEYINPUT31), .B1(KEYINPUT73), .B2(new_n304), .ZN(new_n711));
  AOI21_X1  g525(.A(G902), .B1(new_n711), .B2(new_n315), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n635), .B(new_n699), .C1(new_n712), .C2(new_n187), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n602), .A2(new_n686), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n675), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G125), .ZN(G27));
  AOI21_X1  g531(.A(new_n187), .B1(new_n325), .B2(new_n331), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT75), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n319), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n712), .A2(KEYINPUT110), .A3(KEYINPUT32), .A4(new_n187), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n719), .A2(new_n721), .A3(new_n314), .A4(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n449), .A2(new_n600), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(new_n590), .A3(new_n614), .A4(new_n650), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n391), .A2(new_n683), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT107), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n395), .B1(new_n385), .B2(new_n390), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n725), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  AND4_X1   g545(.A1(KEYINPUT42), .A2(new_n723), .A3(new_n522), .A4(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n336), .A2(new_n522), .ZN(new_n734));
  INV_X1    g548(.A(new_n725), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n728), .A2(new_n729), .ZN(new_n736));
  AOI211_X1 g550(.A(KEYINPUT107), .B(new_n395), .C1(new_n385), .C2(new_n390), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n733), .B1(new_n734), .B2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n731), .A2(KEYINPUT108), .A3(new_n336), .A4(new_n522), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n732), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n205), .ZN(G33));
  NAND2_X1  g559(.A1(new_n727), .A2(new_n730), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n652), .A2(new_n724), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n746), .A2(new_n336), .A3(new_n522), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  NOR2_X1   g564(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n612), .A2(new_n590), .A3(new_n613), .ZN(new_n753));
  AND2_X1   g567(.A1(KEYINPUT111), .A2(KEYINPUT43), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n614), .A2(new_n621), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n751), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n596), .A3(new_n635), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n758), .A2(new_n596), .A3(KEYINPUT44), .A4(new_n635), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n724), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n389), .A2(KEYINPUT45), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT45), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n387), .B2(new_n388), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n768), .A3(G469), .ZN(new_n769));
  INV_X1    g583(.A(new_n386), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(KEYINPUT46), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n385), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT46), .B1(new_n769), .B2(new_n770), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n683), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(new_n657), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n761), .A2(KEYINPUT112), .A3(new_n724), .A4(new_n762), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n765), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT113), .B(G137), .Z(new_n779));
  XNOR2_X1  g593(.A(new_n778), .B(new_n779), .ZN(G39));
  OR2_X1    g594(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n774), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n336), .A2(new_n522), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n774), .A2(KEYINPUT114), .A3(KEYINPUT47), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n784), .A2(new_n735), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  NAND2_X1  g602(.A1(new_n687), .A2(new_n724), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n522), .A2(new_n452), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n789), .A2(new_n666), .A3(new_n615), .A4(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n723), .A2(new_n522), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n758), .A2(new_n452), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n789), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT48), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(G952), .A3(new_n286), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n789), .A2(new_n666), .A3(new_n790), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n798), .B(new_n621), .C1(new_n613), .C2(new_n612), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n794), .A2(new_n714), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n784), .A2(new_n786), .B1(new_n396), .B2(new_n705), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n522), .B(new_n699), .C1(new_n712), .C2(new_n187), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n649), .B1(new_n755), .B2(new_n757), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n804), .A3(new_n724), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT118), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n799), .B(new_n800), .C1(new_n801), .C2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n793), .A2(new_n802), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n668), .A2(new_n450), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n687), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT50), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT117), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g628(.A(KEYINPUT117), .B(KEYINPUT51), .C1(new_n807), .C2(new_n811), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n791), .B(new_n797), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n458), .B1(new_n615), .B2(new_n622), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n597), .A2(new_n598), .A3(new_n522), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n592), .A2(new_n639), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n629), .A2(new_n651), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n336), .A2(new_n642), .A3(new_n724), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n746), .A2(new_n714), .A3(new_n735), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n749), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n820), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n653), .A2(new_n677), .A3(new_n716), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n391), .A2(new_n659), .A3(new_n683), .A4(new_n650), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT115), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n646), .A2(new_n667), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n666), .A2(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT52), .B1(new_n827), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n653), .A2(new_n677), .A3(new_n716), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n829), .A2(new_n831), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT52), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n826), .B1(new_n833), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n688), .A2(new_n691), .A3(new_n694), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n709), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n840), .B1(new_n841), .B2(new_n732), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n817), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n592), .A2(new_n639), .A3(new_n819), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n822), .A2(new_n823), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n749), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n836), .B1(new_n834), .B2(new_n835), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n827), .A2(KEYINPUT52), .A3(new_n832), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n688), .A2(new_n691), .A3(new_n694), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n702), .A2(new_n708), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n744), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n849), .A2(new_n853), .A3(KEYINPUT53), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n843), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT54), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT116), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n857), .B1(new_n744), .B2(new_n852), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n840), .B(KEYINPUT116), .C1(new_n841), .C2(new_n732), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(new_n849), .A3(KEYINPUT53), .A4(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(new_n843), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n808), .A2(new_n715), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n816), .A2(new_n856), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n451), .A2(new_n286), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n705), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n867), .A2(KEYINPUT49), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n450), .B1(new_n867), .B2(KEYINPUT49), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n868), .A2(new_n869), .A3(new_n668), .A4(new_n756), .ZN(new_n870));
  INV_X1    g684(.A(new_n666), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n870), .A2(new_n397), .A3(new_n522), .A4(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n866), .A2(new_n872), .ZN(G75));
  NAND2_X1  g687(.A1(new_n419), .A2(new_n421), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(new_n427), .Z(new_n875));
  XNOR2_X1  g689(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n875), .B(new_n876), .Z(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n188), .B1(new_n860), .B2(new_n843), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(G210), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI211_X1 g696(.A(KEYINPUT56), .B(new_n877), .C1(new_n879), .C2(G210), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n286), .A2(G952), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G51));
  NAND2_X1  g699(.A1(new_n770), .A2(KEYINPUT57), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n770), .A2(KEYINPUT57), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n860), .A2(new_n861), .A3(new_n843), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n861), .B1(new_n860), .B2(new_n843), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n886), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n383), .ZN(new_n891));
  INV_X1    g705(.A(new_n769), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n879), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n884), .B1(new_n891), .B2(new_n893), .ZN(G54));
  NAND2_X1  g708(.A1(new_n860), .A2(new_n843), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n896));
  INV_X1    g710(.A(new_n581), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT120), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n884), .B1(new_n896), .B2(new_n897), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n900), .B(new_n188), .C1(new_n860), .C2(new_n843), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n902), .A3(G475), .A4(new_n581), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n898), .A2(new_n899), .A3(new_n903), .ZN(G60));
  INV_X1    g718(.A(new_n884), .ZN(new_n905));
  XNOR2_X1  g719(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n549), .A2(new_n188), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n906), .B(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(new_n856), .B2(new_n862), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n606), .A2(new_n607), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n905), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n889), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n910), .B(new_n908), .C1(new_n913), .C2(new_n862), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(G63));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n916));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT60), .Z(new_n918));
  NAND3_X1  g732(.A1(new_n895), .A2(new_n633), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n905), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n504), .B1(new_n895), .B2(new_n918), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n921), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(KEYINPUT61), .A3(new_n905), .A4(new_n919), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n924), .ZN(G66));
  INV_X1    g739(.A(new_n424), .ZN(new_n926));
  OAI21_X1  g740(.A(G953), .B1(new_n454), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n852), .A2(new_n820), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n927), .B1(new_n928), .B2(G953), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n874), .B1(G898), .B2(new_n286), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G69));
  NAND2_X1  g745(.A1(new_n778), .A2(new_n827), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n276), .A2(new_n249), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n575), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n776), .A2(new_n792), .A3(new_n830), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n744), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n939), .A2(new_n938), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n941), .A2(new_n749), .A3(new_n787), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n934), .A2(new_n937), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT62), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n673), .B2(new_n834), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n671), .A2(new_n827), .A3(KEYINPUT62), .A4(new_n672), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n778), .A2(new_n787), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n734), .B1(new_n615), .B2(new_n622), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n949), .A2(new_n598), .A3(new_n656), .A4(new_n724), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n947), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(G953), .B1(new_n951), .B2(new_n936), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n647), .B1(new_n936), .B2(new_n338), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n286), .B1(new_n937), .B2(G227), .ZN(new_n954));
  AOI22_X1  g768(.A1(new_n943), .A2(new_n952), .B1(new_n953), .B2(new_n954), .ZN(G72));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT63), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n843), .B2(new_n854), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n324), .A2(new_n291), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n310), .B1(new_n959), .B2(KEYINPUT126), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(KEYINPUT126), .B2(new_n959), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n884), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT125), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n947), .A2(new_n948), .A3(new_n928), .A4(new_n950), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n957), .B(KEYINPUT124), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n324), .A2(new_n292), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n967), .ZN(new_n969));
  AOI211_X1 g783(.A(KEYINPUT125), .B(new_n969), .C1(new_n964), .C2(new_n965), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n962), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n324), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n934), .A2(new_n928), .A3(new_n940), .A4(new_n942), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n972), .B(new_n291), .C1(new_n973), .C2(new_n965), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n971), .A2(new_n974), .ZN(G57));
endmodule


