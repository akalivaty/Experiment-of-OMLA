//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n550, new_n551, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n564, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT66), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  INV_X1    g030(.A(G2105), .ZN(new_n456));
  NAND3_X1  g031(.A1(new_n456), .A2(G101), .A3(G2104), .ZN(new_n457));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n457), .B(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n460), .A2(G137), .A3(new_n456), .ZN(new_n461));
  AOI22_X1  g036(.A1(new_n460), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(new_n459), .B(new_n461), .C1(new_n462), .C2(new_n456), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G160));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n460), .A2(KEYINPUT68), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(new_n472), .A3(G2105), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n471), .A2(new_n472), .A3(new_n456), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n456), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  AND2_X1   g057(.A1(G126), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n465), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  NOR2_X1   g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n460), .A2(new_n483), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n456), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n460), .A2(KEYINPUT4), .A3(G138), .A4(new_n456), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G164));
  XNOR2_X1  g069(.A(KEYINPUT6), .B(G651), .ZN(new_n495));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G543), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n495), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G88), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n495), .A2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G50), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n497), .A2(new_n499), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G62), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(new_n508), .B(KEYINPUT69), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n505), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G166));
  AOI22_X1  g088(.A1(new_n495), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n497), .A2(new_n499), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n502), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n516), .B1(G51), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(new_n520), .ZN(G286));
  INV_X1    g096(.A(G286), .ZN(G168));
  AOI22_X1  g097(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G90), .ZN(new_n526));
  INV_X1    g101(.A(G52), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n500), .A2(new_n526), .B1(new_n502), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(KEYINPUT70), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n529), .A2(KEYINPUT70), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n525), .B1(new_n531), .B2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  NAND2_X1  g109(.A1(G68), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G56), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n515), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(KEYINPUT71), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(KEYINPUT71), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n538), .A2(G651), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G81), .ZN(new_n541));
  INV_X1    g116(.A(G43), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n500), .A2(new_n541), .B1(new_n502), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(G188));
  INV_X1    g127(.A(new_n500), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G91), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  INV_X1    g130(.A(G53), .ZN(new_n556));
  OAI211_X1 g131(.A(KEYINPUT72), .B(new_n555), .C1(new_n502), .C2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n554), .B(new_n557), .C1(new_n524), .C2(new_n558), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT72), .B(KEYINPUT9), .Z(new_n560));
  NOR3_X1   g135(.A1(new_n502), .A2(new_n560), .A3(new_n556), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G299));
  NAND3_X1  g138(.A1(new_n505), .A2(new_n511), .A3(KEYINPUT73), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n524), .B1(new_n507), .B2(new_n509), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n566), .B2(new_n504), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G303));
  NAND2_X1  g143(.A1(new_n553), .A2(G87), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n517), .A2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  AND3_X1   g147(.A1(new_n497), .A2(new_n499), .A3(G61), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT74), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n576), .A2(G73), .A3(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n506), .A2(G86), .A3(new_n495), .ZN(new_n580));
  AND2_X1   g155(.A1(KEYINPUT6), .A2(G651), .ZN(new_n581));
  NOR2_X1   g156(.A1(KEYINPUT6), .A2(G651), .ZN(new_n582));
  OAI211_X1 g157(.A(G48), .B(G543), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(KEYINPUT75), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n495), .A2(new_n585), .A3(G48), .A4(G543), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n579), .A2(new_n580), .A3(new_n584), .A4(new_n586), .ZN(G305));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  INV_X1    g163(.A(G72), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n515), .A2(new_n588), .B1(new_n589), .B2(new_n496), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n590), .A2(KEYINPUT76), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(KEYINPUT76), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n591), .A2(G651), .A3(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n553), .A2(G85), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n517), .A2(G47), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n594), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n595), .A2(new_n596), .A3(new_n597), .A4(new_n598), .ZN(G290));
  AND3_X1   g174(.A1(new_n506), .A2(G92), .A3(new_n495), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n515), .B2(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(G54), .A2(new_n517), .B1(new_n604), .B2(G651), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G171), .B2(new_n607), .ZN(G284));
  OAI21_X1  g184(.A(new_n608), .B1(G171), .B2(new_n607), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n562), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(G868), .B2(new_n562), .ZN(G280));
  INV_X1    g188(.A(new_n606), .ZN(new_n614));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT78), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(G868), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(G868), .B2(new_n546), .ZN(G323));
  XOR2_X1   g195(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n621));
  XNOR2_X1  g196(.A(G323), .B(new_n621), .ZN(G282));
  NAND2_X1  g197(.A1(new_n474), .A2(G123), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n477), .A2(G135), .ZN(new_n624));
  OR2_X1    g199(.A1(G99), .A2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n625), .B(G2104), .C1(G111), .C2(new_n456), .ZN(new_n626));
  AND3_X1   g201(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2096), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n456), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT80), .B(G2100), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n628), .A2(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2435), .ZN(new_n636));
  XOR2_X1   g211(.A(G2427), .B(G2438), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT14), .ZN(new_n639));
  XOR2_X1   g214(.A(G2451), .B(G2454), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n644), .B(new_n645), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G14), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2072), .B(G2078), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(KEYINPUT17), .ZN(new_n653));
  AOI211_X1 g228(.A(new_n649), .B(new_n652), .C1(new_n653), .C2(new_n651), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT81), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  INV_X1    g232(.A(new_n653), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(new_n649), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n655), .B(new_n657), .C1(new_n651), .C2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT82), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1991), .B(G1996), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT21), .ZN(new_n667));
  XOR2_X1   g242(.A(G1956), .B(G2474), .Z(new_n668));
  XOR2_X1   g243(.A(G1961), .B(G1966), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT83), .ZN(new_n671));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT84), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n668), .A2(new_n669), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(new_n670), .ZN(new_n679));
  MUX2_X1   g254(.A(new_n679), .B(new_n678), .S(new_n673), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n676), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n681), .B1(new_n676), .B2(new_n680), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n667), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n676), .A2(new_n680), .ZN(new_n686));
  INV_X1    g261(.A(new_n681), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n667), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n682), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1981), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT22), .ZN(new_n692));
  AND3_X1   g267(.A1(new_n685), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n692), .B1(new_n685), .B2(new_n690), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NOR2_X1   g272(.A1(G301), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G1961), .ZN(new_n699));
  NOR2_X1   g274(.A1(G5), .A2(G16), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(G29), .A2(G32), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n474), .A2(G129), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n477), .A2(G141), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT26), .Z(new_n706));
  NAND3_X1  g281(.A1(new_n456), .A2(G105), .A3(G2104), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT93), .Z(new_n708));
  NAND4_X1  g283(.A1(new_n703), .A2(new_n704), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n702), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n701), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n477), .A2(G139), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(new_n456), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n456), .A2(G103), .A3(G2104), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT25), .Z(new_n718));
  AND3_X1   g293(.A1(new_n714), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G29), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n720), .B(G2072), .C1(G29), .C2(G33), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  AND2_X1   g297(.A1(KEYINPUT87), .A2(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(KEYINPUT87), .A2(G29), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT24), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(G34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(G34), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n463), .B2(new_n710), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n720), .B1(G29), .B2(G33), .ZN(new_n734));
  INV_X1    g309(.A(G2072), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AND3_X1   g311(.A1(new_n713), .A2(new_n722), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n627), .A2(new_n725), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT95), .Z(new_n739));
  OAI21_X1  g314(.A(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n726), .A2(G27), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G164), .B2(new_n726), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT96), .B(G2078), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT97), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n742), .B(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(G28), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(G28), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n747), .A2(new_n748), .A3(new_n710), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n739), .A2(new_n740), .A3(new_n745), .A4(new_n749), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n711), .A2(new_n712), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT31), .B(G11), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n697), .A2(G21), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G168), .B2(new_n697), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT94), .B(G1966), .Z(new_n757));
  INV_X1    g332(.A(new_n757), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n756), .B(new_n758), .ZN(new_n759));
  NAND4_X1  g334(.A1(new_n737), .A2(new_n753), .A3(new_n754), .A4(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT98), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT99), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n726), .A2(G35), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G162), .B2(new_n726), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT29), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G2090), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n763), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n766), .A2(KEYINPUT99), .A3(G2090), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n697), .A2(G4), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n614), .B2(new_n697), .ZN(new_n772));
  INV_X1    g347(.A(G1348), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n762), .A2(new_n769), .A3(new_n770), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n760), .A2(new_n761), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n766), .A2(G2090), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n697), .A2(G19), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n546), .B2(new_n697), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G1341), .Z(new_n781));
  MUX2_X1   g356(.A(G6), .B(G305), .S(G16), .Z(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT32), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1981), .ZN(new_n784));
  OAI21_X1  g359(.A(KEYINPUT90), .B1(G16), .B2(G23), .ZN(new_n785));
  OR3_X1    g360(.A1(KEYINPUT90), .A2(G16), .A3(G23), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n785), .B(new_n786), .C1(G288), .C2(new_n697), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT33), .B(G1976), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n697), .A2(G22), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n697), .ZN(new_n791));
  AND2_X1   g366(.A1(new_n791), .A2(G1971), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n791), .A2(G1971), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n789), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n784), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT34), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G16), .A2(G24), .ZN(new_n798));
  XNOR2_X1  g373(.A(G290), .B(KEYINPUT89), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(G16), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(G1986), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n726), .A2(G25), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n474), .A2(G119), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT88), .Z(new_n804));
  OR2_X1    g379(.A1(G95), .A2(G2105), .ZN(new_n805));
  INV_X1    g380(.A(G107), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n465), .B1(new_n806), .B2(G2105), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n477), .A2(G131), .B1(new_n805), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n804), .A2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n802), .B1(new_n810), .B2(new_n726), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT35), .B(G1991), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n811), .B(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n797), .A2(new_n801), .A3(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n816));
  NAND2_X1  g391(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n815), .A2(new_n817), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n778), .A2(new_n781), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n697), .A2(KEYINPUT23), .A3(G20), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT23), .ZN(new_n822));
  INV_X1    g397(.A(G20), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n823), .B2(G16), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n821), .B(new_n824), .C1(new_n562), .C2(new_n697), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1956), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n474), .A2(G128), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n477), .A2(G140), .ZN(new_n828));
  NOR2_X1   g403(.A1(G104), .A2(G2105), .ZN(new_n829));
  OAI21_X1  g404(.A(G2104), .B1(new_n456), .B2(G116), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n827), .B(new_n828), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G29), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n726), .A2(KEYINPUT28), .A3(G26), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT28), .B1(new_n726), .B2(G26), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G2067), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n820), .A2(new_n826), .A3(new_n837), .ZN(G311));
  AND3_X1   g413(.A1(new_n778), .A2(new_n818), .A3(new_n819), .ZN(new_n839));
  INV_X1    g414(.A(new_n826), .ZN(new_n840));
  INV_X1    g415(.A(new_n837), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .A4(new_n781), .ZN(G150));
  AOI22_X1  g417(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(new_n524), .ZN(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  INV_X1    g420(.A(G55), .ZN(new_n846));
  OAI22_X1  g421(.A1(new_n500), .A2(new_n845), .B1(new_n502), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n546), .A2(new_n849), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n545), .A2(new_n848), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n606), .A2(new_n615), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n852), .B1(new_n859), .B2(G860), .ZN(G145));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n466), .A2(new_n468), .A3(new_n483), .ZN(new_n862));
  OAI21_X1  g437(.A(G2104), .B1(new_n456), .B2(G114), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(new_n486), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n861), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n484), .A2(G2105), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n487), .A2(new_n866), .A3(G2104), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n466), .A2(new_n468), .A3(new_n483), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n868), .A3(KEYINPUT101), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n491), .A2(new_n492), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n831), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n709), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n719), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G142), .ZN(new_n877));
  OR3_X1    g452(.A1(new_n476), .A2(KEYINPUT102), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n474), .A2(G130), .ZN(new_n879));
  OR2_X1    g454(.A1(G106), .A2(G2105), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n880), .B(G2104), .C1(G118), .C2(new_n456), .ZN(new_n881));
  OAI21_X1  g456(.A(KEYINPUT102), .B1(new_n476), .B2(new_n877), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n878), .A2(new_n879), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n630), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(new_n809), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n885), .A2(KEYINPUT103), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(KEYINPUT103), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n876), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n875), .A2(new_n886), .A3(new_n887), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n481), .B(G160), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n627), .ZN(new_n893));
  AOI21_X1  g468(.A(G37), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  INV_X1    g470(.A(new_n885), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n890), .B(new_n895), .C1(new_n896), .C2(new_n875), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g474(.A1(new_n849), .A2(new_n607), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n606), .A2(new_n562), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n901), .A2(KEYINPUT105), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(KEYINPUT105), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n614), .A2(G299), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n904), .B(new_n908), .ZN(new_n909));
  AND2_X1   g484(.A1(new_n902), .A2(new_n903), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n907), .B1(new_n911), .B2(new_n906), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n618), .B(new_n855), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n911), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n916), .B(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n512), .B(G288), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(G305), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(G290), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n917), .B2(KEYINPUT42), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n919), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n900), .B1(new_n924), .B2(new_n607), .ZN(G295));
  OAI21_X1  g500(.A(new_n900), .B1(new_n924), .B2(new_n607), .ZN(G331));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n928));
  XNOR2_X1  g503(.A(G301), .B(G168), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n855), .ZN(new_n930));
  NAND2_X1  g505(.A1(G171), .A2(G286), .ZN(new_n931));
  NAND2_X1  g506(.A1(G301), .A2(G168), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n853), .A3(new_n854), .A4(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n928), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT108), .B1(new_n929), .B2(new_n855), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(KEYINPUT41), .B2(new_n905), .ZN(new_n937));
  INV_X1    g512(.A(new_n905), .ZN(new_n938));
  OAI22_X1  g513(.A1(new_n934), .A2(new_n935), .B1(new_n938), .B2(new_n906), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n930), .A2(new_n933), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n937), .A2(KEYINPUT41), .B1(new_n941), .B2(new_n911), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n927), .B1(new_n942), .B2(new_n922), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n936), .A2(new_n911), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n912), .A2(new_n940), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n922), .A3(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n946), .B(KEYINPUT110), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT43), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n946), .B(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n936), .A2(new_n911), .B1(new_n912), .B2(new_n940), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n927), .B1(new_n952), .B2(new_n922), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT109), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n955), .B(new_n927), .C1(new_n952), .C2(new_n922), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n950), .A2(new_n951), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n948), .A2(new_n957), .A3(KEYINPUT44), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n951), .B1(new_n943), .B2(new_n947), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n950), .A2(KEYINPUT43), .A3(new_n954), .A4(new_n956), .ZN(new_n960));
  XNOR2_X1  g535(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G1956), .ZN(new_n964));
  XNOR2_X1  g539(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1384), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n966), .B1(new_n872), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G40), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n463), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n493), .A2(new_n971), .A3(new_n967), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n964), .B1(new_n968), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(G113), .A2(G2104), .ZN(new_n975));
  INV_X1    g550(.A(G125), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(new_n469), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G2105), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n978), .A2(G40), .A3(new_n461), .A4(new_n459), .ZN(new_n979));
  AOI21_X1  g554(.A(G1384), .B1(new_n870), .B2(new_n871), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(new_n980), .B2(KEYINPUT45), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n493), .A2(new_n967), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT56), .B(G2072), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n981), .A2(new_n985), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT57), .ZN(new_n988));
  NOR2_X1   g563(.A1(G299), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n562), .A2(KEYINPUT57), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n974), .B(new_n987), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n872), .A2(new_n967), .A3(new_n966), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n982), .A2(KEYINPUT50), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n992), .A2(new_n970), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n980), .A2(new_n970), .ZN(new_n995));
  OAI22_X1  g570(.A1(new_n994), .A2(G1348), .B1(G2067), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n991), .A2(new_n614), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n987), .A2(new_n974), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n562), .B(new_n988), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT59), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n872), .A2(KEYINPUT45), .A3(new_n967), .ZN(new_n1003));
  INV_X1    g578(.A(G1996), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n970), .A4(new_n985), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n981), .A2(KEYINPUT119), .A3(new_n1004), .A4(new_n985), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT58), .B(G1341), .Z(new_n1009));
  NAND2_X1  g584(.A1(new_n995), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT121), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n546), .A2(KEYINPUT120), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1012), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1002), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT121), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(KEYINPUT59), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT122), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT61), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1000), .A2(new_n991), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1022), .A2(KEYINPUT61), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n992), .A2(new_n970), .A3(new_n993), .ZN(new_n1027));
  INV_X1    g602(.A(new_n995), .ZN(new_n1028));
  INV_X1    g603(.A(G2067), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1027), .A2(new_n773), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n606), .B(KEYINPUT123), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(KEYINPUT60), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n614), .A2(KEYINPUT123), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT60), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1033), .B1(new_n996), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n996), .A2(new_n1034), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1000), .A2(new_n991), .A3(new_n1022), .A4(KEYINPUT61), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1026), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1001), .B1(new_n1021), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G2078), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n981), .A2(new_n1041), .A3(new_n985), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1042), .A2(new_n1043), .B1(new_n699), .B2(new_n1027), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n493), .A2(new_n967), .A3(new_n983), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n970), .B(new_n1045), .C1(new_n980), .C2(KEYINPUT45), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(KEYINPUT53), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1044), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g623(.A(G301), .B(KEYINPUT54), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1046), .A2(new_n758), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n992), .A2(new_n732), .A3(new_n970), .A4(new_n993), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT124), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT124), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(new_n1055), .A3(new_n1052), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1054), .A2(G168), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G8), .ZN(new_n1058));
  INV_X1    g633(.A(G8), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1058), .A2(KEYINPUT51), .B1(G286), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(G8), .B1(new_n1053), .B2(G286), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1062), .A2(KEYINPUT51), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1050), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n995), .A2(G8), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT113), .B(G1981), .Z(new_n1067));
  NOR2_X1   g642(.A1(G305), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G305), .A2(G1981), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(G305), .A2(KEYINPUT114), .A3(G1981), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1068), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1066), .B1(new_n1073), .B2(KEYINPUT49), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1068), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1072), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT114), .B1(G305), .B2(G1981), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT49), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(KEYINPUT115), .A3(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1065), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(KEYINPUT49), .B(new_n1075), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT116), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1085), .A2(KEYINPUT116), .A3(KEYINPUT49), .A4(new_n1075), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1065), .ZN(new_n1088));
  INV_X1    g663(.A(G1976), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(G288), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1081), .A2(new_n1087), .B1(KEYINPUT52), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT52), .B1(G288), .B2(new_n1089), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1088), .B(new_n1092), .C1(new_n1089), .C2(G288), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1003), .A2(new_n970), .A3(new_n985), .ZN(new_n1095));
  INV_X1    g670(.A(G1971), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n994), .A2(new_n768), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(G303), .A2(G8), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT55), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT55), .ZN(new_n1100));
  NAND3_X1  g675(.A1(G303), .A2(new_n1100), .A3(G8), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  OR3_X1    g677(.A1(new_n1097), .A2(new_n1102), .A3(new_n1059), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  AND2_X1   g679(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n867), .A2(new_n868), .A3(KEYINPUT101), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT101), .B1(new_n867), .B2(new_n868), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n491), .A2(new_n492), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n967), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n965), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1111), .A2(new_n1112), .A3(new_n970), .A4(new_n972), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT117), .B1(new_n968), .B2(new_n973), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1114), .A3(new_n768), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1105), .B1(new_n1117), .B2(G8), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1094), .A2(new_n1104), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1049), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n980), .A2(new_n983), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n981), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1120), .B(new_n1044), .C1(new_n1047), .C2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1040), .A2(new_n1064), .A3(new_n1119), .A4(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1062), .A2(G286), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1102), .B1(new_n1097), .B2(new_n1059), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1091), .A2(new_n1093), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(new_n1088), .A3(new_n1087), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1090), .A2(KEYINPUT52), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1130), .A2(new_n1131), .A3(new_n1093), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1053), .A2(new_n1133), .A3(G8), .A4(G168), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1103), .B1(new_n1118), .B2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1128), .A2(KEYINPUT63), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g711(.A(G1976), .B(G288), .C1(new_n1081), .C2(new_n1087), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1088), .B1(new_n1137), .B2(new_n1068), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT118), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1130), .A2(new_n1131), .A3(new_n1093), .A4(new_n1127), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1126), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT63), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1143));
  AND4_X1   g718(.A1(KEYINPUT118), .A2(new_n1138), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1125), .B1(new_n1139), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1125), .B(KEYINPUT125), .C1(new_n1139), .C2(new_n1144), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1149));
  OR2_X1    g724(.A1(new_n1149), .A2(KEYINPUT62), .ZN(new_n1150));
  AOI21_X1  g725(.A(G301), .B1(new_n1149), .B2(KEYINPUT62), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1150), .A2(new_n1151), .A3(new_n1119), .A4(new_n1048), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1147), .A2(new_n1148), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n810), .A2(new_n813), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n831), .B(new_n1029), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n709), .B(new_n1004), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n809), .A2(new_n812), .ZN(new_n1158));
  NOR3_X1   g733(.A1(new_n1154), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  OR2_X1    g734(.A1(G290), .A2(G1986), .ZN(new_n1160));
  NAND2_X1  g735(.A1(G290), .A2(G1986), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1122), .A2(new_n979), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1153), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1163), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1160), .A2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT48), .Z(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n1166), .B2(new_n1159), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1155), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1163), .B1(new_n1170), .B2(new_n709), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT46), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1172), .B1(new_n1166), .B2(G1996), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1163), .A2(KEYINPUT46), .A3(new_n1004), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1171), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1175), .B(KEYINPUT47), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1158), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1177), .A2(new_n1157), .B1(G2067), .B2(new_n831), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1163), .ZN(new_n1179));
  AND3_X1   g754(.A1(new_n1169), .A2(new_n1176), .A3(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1165), .A2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g756(.A1(new_n664), .A2(KEYINPUT126), .A3(G319), .ZN(new_n1183));
  NAND2_X1  g757(.A1(new_n664), .A2(G319), .ZN(new_n1184));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g760(.A1(new_n695), .A2(new_n647), .A3(new_n1183), .A4(new_n1186), .ZN(new_n1187));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n1188));
  OR2_X1    g762(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI22_X1  g763(.A1(new_n1187), .A2(new_n1188), .B1(new_n894), .B2(new_n897), .ZN(new_n1190));
  AND4_X1   g764(.A1(new_n959), .A2(new_n1189), .A3(new_n1190), .A4(new_n960), .ZN(G308));
  NAND4_X1  g765(.A1(new_n1189), .A2(new_n1190), .A3(new_n959), .A4(new_n960), .ZN(G225));
endmodule


