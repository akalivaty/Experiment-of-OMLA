//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:51 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1142, new_n1143, new_n1144, new_n1145, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1194, new_n1195;
  NOR4_X1   g000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g002(.A(G1), .ZN(new_n203));
  INV_X1    g003(.A(G20), .ZN(new_n204));
  NOR2_X1   g004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g005(.A(new_n205), .ZN(new_n206));
  INV_X1    g006(.A(G116), .ZN(new_n207));
  INV_X1    g007(.A(G270), .ZN(new_n208));
  NOR2_X1   g008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g009(.A1(G97), .A2(G257), .ZN(new_n210));
  INV_X1    g010(.A(G68), .ZN(new_n211));
  INV_X1    g011(.A(G238), .ZN(new_n212));
  INV_X1    g012(.A(G87), .ZN(new_n213));
  INV_X1    g013(.A(G250), .ZN(new_n214));
  OAI221_X1 g014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g015(.A(new_n209), .B(new_n215), .C1(G107), .C2(G264), .ZN(new_n216));
  INV_X1    g016(.A(G50), .ZN(new_n217));
  INV_X1    g017(.A(G226), .ZN(new_n218));
  INV_X1    g018(.A(G77), .ZN(new_n219));
  INV_X1    g019(.A(G244), .ZN(new_n220));
  OAI221_X1 g020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g021(.A(G58), .ZN(new_n222));
  INV_X1    g022(.A(G232), .ZN(new_n223));
  NOR2_X1   g023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g024(.A(new_n206), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g026(.A1(new_n206), .A2(G13), .ZN(new_n227));
  OAI211_X1 g027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  NOR2_X1   g029(.A1(G58), .A2(G68), .ZN(new_n230));
  INV_X1    g030(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  NAND2_X1  g032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR3_X1   g033(.A1(new_n232), .A2(new_n204), .A3(new_n233), .ZN(new_n234));
  NOR3_X1   g034(.A1(new_n226), .A2(new_n229), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g040(.A(new_n240), .B(G264), .ZN(new_n241));
  XNOR2_X1  g041(.A(new_n241), .B(new_n208), .ZN(new_n242));
  XNOR2_X1  g042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g043(.A(G87), .B(G97), .ZN(new_n244));
  INV_X1    g044(.A(G107), .ZN(new_n245));
  XNOR2_X1  g045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g046(.A(new_n246), .B(new_n207), .ZN(new_n247));
  XOR2_X1   g047(.A(G68), .B(G77), .Z(new_n248));
  XOR2_X1   g048(.A(G50), .B(G58), .Z(new_n249));
  XNOR2_X1  g049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  INV_X1    g053(.A(G33), .ZN(new_n254));
  NAND2_X1  g054(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  AND2_X1   g055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g056(.A1(new_n256), .A2(G1698), .ZN(new_n257));
  XNOR2_X1  g057(.A(new_n257), .B(KEYINPUT64), .ZN(new_n258));
  NAND2_X1  g058(.A1(new_n258), .A2(G223), .ZN(new_n259));
  NAND2_X1  g059(.A1(new_n253), .A2(new_n255), .ZN(new_n260));
  NAND2_X1  g060(.A1(new_n260), .A2(G77), .ZN(new_n261));
  NOR2_X1   g061(.A1(new_n260), .A2(G1698), .ZN(new_n262));
  NAND2_X1  g062(.A1(new_n262), .A2(G222), .ZN(new_n263));
  NAND3_X1  g063(.A1(new_n259), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g064(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n265));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g066(.A(G41), .ZN(new_n267));
  INV_X1    g067(.A(G45), .ZN(new_n268));
  AOI21_X1  g068(.A(G1), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g069(.A1(new_n269), .A2(G274), .ZN(new_n270));
  NOR2_X1   g070(.A1(new_n265), .A2(new_n269), .ZN(new_n271));
  NAND2_X1  g071(.A1(new_n271), .A2(G226), .ZN(new_n272));
  NAND3_X1  g072(.A1(new_n266), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g073(.A(new_n273), .ZN(new_n274));
  INV_X1    g074(.A(G179), .ZN(new_n275));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g076(.A(G20), .B1(new_n231), .B2(G50), .ZN(new_n277));
  INV_X1    g077(.A(G150), .ZN(new_n278));
  NOR2_X1   g078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g080(.A1(new_n204), .A2(G33), .ZN(new_n281));
  XNOR2_X1  g081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  OAI221_X1 g082(.A(new_n277), .B1(new_n278), .B2(new_n280), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g083(.A(new_n233), .ZN(new_n284));
  AOI21_X1  g084(.A(new_n284), .B1(new_n205), .B2(G33), .ZN(new_n285));
  INV_X1    g085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g086(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g087(.A1(new_n204), .A2(G1), .ZN(new_n288));
  NOR2_X1   g088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g089(.A1(new_n289), .A2(G50), .ZN(new_n290));
  NAND2_X1  g090(.A1(new_n288), .A2(G13), .ZN(new_n291));
  OAI211_X1 g091(.A(new_n287), .B(new_n290), .C1(G50), .C2(new_n291), .ZN(new_n292));
  OAI211_X1 g092(.A(new_n276), .B(new_n292), .C1(G169), .C2(new_n274), .ZN(new_n293));
  INV_X1    g093(.A(new_n270), .ZN(new_n294));
  NAND2_X1  g094(.A1(new_n258), .A2(G238), .ZN(new_n295));
  AOI22_X1  g095(.A1(new_n262), .A2(G232), .B1(G107), .B2(new_n260), .ZN(new_n296));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g097(.A(new_n294), .B1(new_n297), .B2(new_n265), .ZN(new_n298));
  NAND2_X1  g098(.A1(new_n271), .A2(G244), .ZN(new_n299));
  AND2_X1   g099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n275), .ZN(new_n301));
  OAI22_X1  g101(.A1(new_n282), .A2(new_n280), .B1(new_n204), .B2(new_n219), .ZN(new_n302));
  XNOR2_X1  g102(.A(new_n302), .B(KEYINPUT65), .ZN(new_n303));
  XOR2_X1   g103(.A(KEYINPUT15), .B(G87), .Z(new_n304));
  INV_X1    g104(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g105(.A(new_n303), .B1(new_n281), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g106(.A1(new_n285), .A2(new_n291), .ZN(new_n307));
  NAND2_X1  g107(.A1(new_n307), .A2(KEYINPUT66), .ZN(new_n308));
  INV_X1    g108(.A(KEYINPUT66), .ZN(new_n309));
  NAND3_X1  g109(.A1(new_n285), .A2(new_n309), .A3(new_n291), .ZN(new_n310));
  AOI21_X1  g110(.A(new_n288), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AOI22_X1  g111(.A1(new_n306), .A2(new_n286), .B1(G77), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g112(.A(new_n312), .B1(G77), .B2(new_n291), .ZN(new_n313));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n314));
  INV_X1    g114(.A(G169), .ZN(new_n315));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  INV_X1    g117(.A(KEYINPUT10), .ZN(new_n318));
  NAND2_X1  g118(.A1(new_n274), .A2(G190), .ZN(new_n319));
  XNOR2_X1  g119(.A(new_n292), .B(KEYINPUT9), .ZN(new_n320));
  AND2_X1   g120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g121(.A(G200), .ZN(new_n322));
  NOR2_X1   g122(.A1(new_n274), .A2(new_n322), .ZN(new_n323));
  INV_X1    g123(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g124(.A(new_n318), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g125(.A1(new_n319), .A2(new_n320), .ZN(new_n326));
  NOR3_X1   g126(.A1(new_n326), .A2(new_n323), .A3(KEYINPUT10), .ZN(new_n327));
  OAI211_X1 g127(.A(new_n293), .B(new_n317), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  NAND2_X1  g128(.A1(G33), .A2(G97), .ZN(new_n329));
  NAND2_X1  g129(.A1(new_n223), .A2(G1698), .ZN(new_n330));
  OAI21_X1  g130(.A(new_n330), .B1(G226), .B2(G1698), .ZN(new_n331));
  OAI21_X1  g131(.A(new_n329), .B1(new_n331), .B2(new_n260), .ZN(new_n332));
  AOI21_X1  g132(.A(new_n294), .B1(new_n332), .B2(new_n265), .ZN(new_n333));
  INV_X1    g133(.A(new_n271), .ZN(new_n334));
  OAI21_X1  g134(.A(new_n333), .B1(new_n212), .B2(new_n334), .ZN(new_n335));
  OR2_X1    g135(.A1(new_n335), .A2(KEYINPUT13), .ZN(new_n336));
  NAND2_X1  g136(.A1(new_n335), .A2(KEYINPUT13), .ZN(new_n337));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g138(.A1(new_n338), .A2(G169), .ZN(new_n339));
  NAND2_X1  g139(.A1(new_n339), .A2(KEYINPUT14), .ZN(new_n340));
  INV_X1    g140(.A(KEYINPUT14), .ZN(new_n341));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n341), .A3(G169), .ZN(new_n342));
  OAI211_X1 g142(.A(new_n340), .B(new_n342), .C1(new_n275), .C2(new_n338), .ZN(new_n343));
  NAND2_X1  g143(.A1(new_n311), .A2(G68), .ZN(new_n344));
  INV_X1    g144(.A(new_n291), .ZN(new_n345));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n211), .ZN(new_n346));
  XNOR2_X1  g146(.A(new_n346), .B(KEYINPUT12), .ZN(new_n347));
  NAND2_X1  g147(.A1(new_n279), .A2(G50), .ZN(new_n348));
  XNOR2_X1  g148(.A(new_n348), .B(KEYINPUT67), .ZN(new_n349));
  OAI22_X1  g149(.A1(new_n281), .A2(new_n219), .B1(new_n204), .B2(G68), .ZN(new_n350));
  OAI21_X1  g150(.A(new_n286), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g151(.A1(new_n351), .A2(KEYINPUT11), .ZN(new_n352));
  NOR2_X1   g152(.A1(new_n351), .A2(KEYINPUT11), .ZN(new_n353));
  OAI211_X1 g153(.A(new_n344), .B(new_n347), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g154(.A1(new_n343), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g155(.A1(new_n338), .A2(G200), .ZN(new_n356));
  INV_X1    g156(.A(new_n354), .ZN(new_n357));
  INV_X1    g157(.A(G190), .ZN(new_n358));
  OAI211_X1 g158(.A(new_n356), .B(new_n357), .C1(new_n358), .C2(new_n338), .ZN(new_n359));
  NAND2_X1  g159(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  INV_X1    g160(.A(KEYINPUT68), .ZN(new_n361));
  OAI21_X1  g161(.A(new_n361), .B1(new_n252), .B2(G33), .ZN(new_n362));
  NAND3_X1  g162(.A1(new_n254), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n363));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n253), .ZN(new_n365));
  INV_X1    g165(.A(KEYINPUT7), .ZN(new_n366));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n366), .A3(new_n204), .ZN(new_n367));
  AOI22_X1  g167(.A1(new_n362), .A2(new_n363), .B1(new_n252), .B2(G33), .ZN(new_n368));
  OAI21_X1  g168(.A(KEYINPUT7), .B1(new_n368), .B2(G20), .ZN(new_n369));
  NAND3_X1  g169(.A1(new_n367), .A2(new_n369), .A3(G68), .ZN(new_n370));
  AND2_X1   g170(.A1(G58), .A2(G68), .ZN(new_n371));
  OAI21_X1  g171(.A(G20), .B1(new_n371), .B2(new_n230), .ZN(new_n372));
  NAND2_X1  g172(.A1(new_n279), .A2(G159), .ZN(new_n373));
  AND3_X1   g173(.A1(new_n372), .A2(KEYINPUT69), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g174(.A(KEYINPUT69), .B1(new_n372), .B2(new_n373), .ZN(new_n375));
  NOR2_X1   g175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g176(.A1(new_n370), .A2(KEYINPUT16), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g177(.A1(new_n377), .A2(KEYINPUT70), .ZN(new_n378));
  INV_X1    g178(.A(KEYINPUT16), .ZN(new_n379));
  INV_X1    g179(.A(new_n376), .ZN(new_n380));
  OAI21_X1  g180(.A(new_n366), .B1(new_n256), .B2(G20), .ZN(new_n381));
  NAND3_X1  g181(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n382));
  AOI21_X1  g182(.A(new_n211), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g183(.A(new_n379), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  INV_X1    g184(.A(KEYINPUT70), .ZN(new_n385));
  NAND4_X1  g185(.A1(new_n370), .A2(new_n385), .A3(KEYINPUT16), .A4(new_n376), .ZN(new_n386));
  NAND4_X1  g186(.A1(new_n378), .A2(new_n286), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  INV_X1    g187(.A(new_n282), .ZN(new_n388));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n291), .ZN(new_n389));
  AOI21_X1  g189(.A(new_n389), .B1(new_n289), .B2(new_n388), .ZN(new_n390));
  NAND2_X1  g190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  OR2_X1    g191(.A1(G223), .A2(G1698), .ZN(new_n392));
  NAND2_X1  g192(.A1(new_n218), .A2(G1698), .ZN(new_n393));
  NAND4_X1  g193(.A1(new_n364), .A2(new_n253), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g194(.A1(G33), .A2(G87), .ZN(new_n395));
  NAND2_X1  g195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n265), .ZN(new_n397));
  AOI21_X1  g197(.A(new_n294), .B1(new_n271), .B2(G232), .ZN(new_n398));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n275), .A3(new_n398), .ZN(new_n399));
  INV_X1    g199(.A(KEYINPUT71), .ZN(new_n400));
  INV_X1    g200(.A(new_n265), .ZN(new_n401));
  AOI21_X1  g201(.A(new_n401), .B1(new_n394), .B2(new_n395), .ZN(new_n402));
  INV_X1    g202(.A(new_n269), .ZN(new_n403));
  NAND3_X1  g203(.A1(new_n401), .A2(G232), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n270), .ZN(new_n405));
  OAI21_X1  g205(.A(new_n315), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  AND3_X1   g206(.A1(new_n399), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g207(.A(new_n400), .B1(new_n399), .B2(new_n406), .ZN(new_n408));
  NOR3_X1   g208(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT72), .ZN(new_n409));
  INV_X1    g209(.A(KEYINPUT72), .ZN(new_n410));
  AOI21_X1  g210(.A(G169), .B1(new_n397), .B2(new_n398), .ZN(new_n411));
  NOR3_X1   g211(.A1(new_n402), .A2(new_n405), .A3(G179), .ZN(new_n412));
  OAI21_X1  g212(.A(KEYINPUT71), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n400), .A3(new_n406), .ZN(new_n414));
  AOI21_X1  g214(.A(new_n410), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g215(.A(new_n391), .B1(new_n409), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g216(.A(KEYINPUT73), .B(KEYINPUT18), .ZN(new_n417));
  NAND2_X1  g217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g218(.A1(new_n397), .A2(new_n398), .ZN(new_n419));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n322), .ZN(new_n420));
  OAI21_X1  g220(.A(new_n420), .B1(G190), .B2(new_n419), .ZN(new_n421));
  XOR2_X1   g221(.A(KEYINPUT74), .B(KEYINPUT17), .Z(new_n422));
  INV_X1    g222(.A(new_n422), .ZN(new_n423));
  NAND4_X1  g223(.A1(new_n387), .A2(new_n390), .A3(new_n421), .A4(new_n423), .ZN(new_n424));
  AND3_X1   g224(.A1(new_n387), .A2(new_n390), .A3(new_n421), .ZN(new_n425));
  NOR2_X1   g225(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n426));
  OAI21_X1  g226(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g227(.A(new_n417), .ZN(new_n428));
  OAI211_X1 g228(.A(new_n391), .B(new_n428), .C1(new_n409), .C2(new_n415), .ZN(new_n429));
  NAND3_X1  g229(.A1(new_n418), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NOR2_X1   g230(.A1(new_n300), .A2(new_n322), .ZN(new_n431));
  NOR2_X1   g231(.A1(new_n314), .A2(new_n358), .ZN(new_n432));
  NOR3_X1   g232(.A1(new_n431), .A2(new_n432), .A3(new_n313), .ZN(new_n433));
  NOR4_X1   g233(.A1(new_n328), .A2(new_n360), .A3(new_n430), .A4(new_n433), .ZN(new_n434));
  NOR2_X1   g234(.A1(new_n204), .A2(G107), .ZN(new_n435));
  XNOR2_X1  g235(.A(new_n435), .B(KEYINPUT23), .ZN(new_n436));
  NAND3_X1  g236(.A1(new_n204), .A2(G33), .A3(G116), .ZN(new_n437));
  INV_X1    g237(.A(KEYINPUT22), .ZN(new_n438));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n213), .ZN(new_n439));
  NAND3_X1  g239(.A1(new_n368), .A2(new_n204), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g240(.A1(new_n253), .A2(new_n255), .A3(new_n204), .A4(G87), .ZN(new_n441));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n438), .ZN(new_n442));
  AND3_X1   g242(.A1(new_n440), .A2(KEYINPUT83), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g243(.A(KEYINPUT83), .B1(new_n440), .B2(new_n442), .ZN(new_n444));
  OAI211_X1 g244(.A(new_n436), .B(new_n437), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  INV_X1    g245(.A(KEYINPUT24), .ZN(new_n446));
  NAND2_X1  g246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g247(.A1(new_n440), .A2(new_n442), .ZN(new_n448));
  INV_X1    g248(.A(KEYINPUT83), .ZN(new_n449));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g250(.A1(new_n440), .A2(KEYINPUT83), .A3(new_n442), .ZN(new_n451));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g252(.A1(new_n452), .A2(KEYINPUT24), .A3(new_n436), .A4(new_n437), .ZN(new_n453));
  NAND3_X1  g253(.A1(new_n447), .A2(new_n453), .A3(new_n286), .ZN(new_n454));
  OAI211_X1 g254(.A(new_n285), .B(new_n291), .C1(G1), .C2(new_n254), .ZN(new_n455));
  INV_X1    g255(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g256(.A1(new_n456), .A2(G107), .ZN(new_n457));
  NOR2_X1   g257(.A1(new_n291), .A2(G107), .ZN(new_n458));
  XNOR2_X1  g258(.A(new_n458), .B(KEYINPUT25), .ZN(new_n459));
  NAND3_X1  g259(.A1(new_n454), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  INV_X1    g260(.A(G1698), .ZN(new_n461));
  OAI21_X1  g261(.A(new_n368), .B1(G257), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g262(.A1(G250), .A2(G1698), .ZN(new_n463));
  INV_X1    g263(.A(G294), .ZN(new_n464));
  OAI22_X1  g264(.A1(new_n462), .A2(new_n463), .B1(new_n254), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g265(.A1(new_n267), .A2(KEYINPUT5), .ZN(new_n466));
  INV_X1    g266(.A(KEYINPUT76), .ZN(new_n467));
  XNOR2_X1  g267(.A(new_n466), .B(new_n467), .ZN(new_n468));
  OAI211_X1 g268(.A(new_n203), .B(G45), .C1(new_n267), .C2(KEYINPUT5), .ZN(new_n469));
  NOR2_X1   g269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n265), .ZN(new_n471));
  AOI22_X1  g271(.A1(new_n265), .A2(new_n465), .B1(new_n471), .B2(G264), .ZN(new_n472));
  XOR2_X1   g272(.A(new_n469), .B(KEYINPUT75), .Z(new_n473));
  NOR2_X1   g273(.A1(new_n468), .A2(new_n265), .ZN(new_n474));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n474), .A3(G274), .ZN(new_n475));
  AOI21_X1  g275(.A(G169), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g276(.A1(new_n472), .A2(new_n475), .ZN(new_n477));
  AOI21_X1  g277(.A(new_n476), .B1(new_n275), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g278(.A1(new_n460), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g279(.A1(new_n479), .A2(KEYINPUT84), .ZN(new_n480));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n481));
  NAND3_X1  g281(.A1(new_n460), .A2(new_n481), .A3(new_n478), .ZN(new_n482));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR3_X1   g283(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n484));
  XNOR2_X1  g284(.A(new_n484), .B(KEYINPUT78), .ZN(new_n485));
  INV_X1    g285(.A(KEYINPUT19), .ZN(new_n486));
  OAI21_X1  g286(.A(new_n204), .B1(new_n329), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g288(.A(G97), .ZN(new_n489));
  OAI21_X1  g289(.A(new_n486), .B1(new_n281), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g290(.A1(new_n368), .A2(new_n204), .A3(G68), .ZN(new_n491));
  NAND3_X1  g291(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g292(.A1(new_n492), .A2(KEYINPUT79), .ZN(new_n493));
  INV_X1    g293(.A(KEYINPUT79), .ZN(new_n494));
  NAND4_X1  g294(.A1(new_n488), .A2(new_n494), .A3(new_n490), .A4(new_n491), .ZN(new_n495));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n286), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g296(.A1(new_n305), .A2(new_n345), .ZN(new_n497));
  NAND2_X1  g297(.A1(new_n456), .A2(new_n304), .ZN(new_n498));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OR2_X1    g299(.A1(new_n499), .A2(KEYINPUT80), .ZN(new_n500));
  OR3_X1    g300(.A1(new_n268), .A2(G1), .A3(G274), .ZN(new_n501));
  AND2_X1   g301(.A1(new_n401), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g302(.A(new_n214), .B1(new_n268), .B2(G1), .ZN(new_n503));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g304(.A1(G238), .A2(G1698), .ZN(new_n505));
  AOI21_X1  g305(.A(new_n505), .B1(new_n220), .B2(G1698), .ZN(new_n506));
  AOI22_X1  g306(.A1(new_n368), .A2(new_n506), .B1(G33), .B2(G116), .ZN(new_n507));
  OAI21_X1  g307(.A(new_n504), .B1(new_n507), .B2(new_n401), .ZN(new_n508));
  NAND2_X1  g308(.A1(new_n508), .A2(G169), .ZN(new_n509));
  OAI21_X1  g309(.A(new_n509), .B1(new_n275), .B2(new_n508), .ZN(new_n510));
  NAND2_X1  g310(.A1(new_n499), .A2(KEYINPUT80), .ZN(new_n511));
  NAND3_X1  g311(.A1(new_n500), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AND2_X1   g312(.A1(new_n496), .A2(new_n497), .ZN(new_n513));
  INV_X1    g313(.A(new_n508), .ZN(new_n514));
  NAND3_X1  g314(.A1(new_n514), .A2(KEYINPUT81), .A3(G190), .ZN(new_n515));
  INV_X1    g315(.A(KEYINPUT81), .ZN(new_n516));
  OAI21_X1  g316(.A(new_n516), .B1(new_n508), .B2(new_n358), .ZN(new_n517));
  NAND2_X1  g317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g318(.A1(new_n456), .A2(G87), .ZN(new_n519));
  NAND2_X1  g319(.A1(new_n508), .A2(G200), .ZN(new_n520));
  NAND4_X1  g320(.A1(new_n513), .A2(new_n518), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  AND2_X1   g321(.A1(new_n512), .A2(new_n521), .ZN(new_n522));
  INV_X1    g322(.A(KEYINPUT77), .ZN(new_n523));
  INV_X1    g323(.A(KEYINPUT4), .ZN(new_n524));
  OAI21_X1  g324(.A(new_n524), .B1(new_n365), .B2(new_n220), .ZN(new_n525));
  NAND2_X1  g325(.A1(G33), .A2(G283), .ZN(new_n526));
  OAI21_X1  g326(.A(KEYINPUT4), .B1(new_n260), .B2(new_n214), .ZN(new_n527));
  NAND2_X1  g327(.A1(new_n527), .A2(G1698), .ZN(new_n528));
  NAND3_X1  g328(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .ZN(new_n529));
  NAND4_X1  g329(.A1(new_n525), .A2(new_n526), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n265), .ZN(new_n531));
  NAND2_X1  g331(.A1(new_n471), .A2(G257), .ZN(new_n532));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n475), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g333(.A(new_n523), .B1(new_n533), .B2(new_n358), .ZN(new_n534));
  INV_X1    g334(.A(new_n475), .ZN(new_n535));
  AOI21_X1  g335(.A(new_n535), .B1(new_n265), .B2(new_n530), .ZN(new_n536));
  NAND4_X1  g336(.A1(new_n536), .A2(KEYINPUT77), .A3(G190), .A4(new_n532), .ZN(new_n537));
  NOR2_X1   g337(.A1(new_n291), .A2(G97), .ZN(new_n538));
  NOR2_X1   g338(.A1(new_n455), .A2(new_n489), .ZN(new_n539));
  NOR2_X1   g339(.A1(new_n280), .A2(new_n219), .ZN(new_n540));
  INV_X1    g340(.A(new_n540), .ZN(new_n541));
  NAND3_X1  g341(.A1(new_n245), .A2(KEYINPUT6), .A3(G97), .ZN(new_n542));
  NOR2_X1   g342(.A1(new_n489), .A2(new_n245), .ZN(new_n543));
  NOR2_X1   g343(.A1(G97), .A2(G107), .ZN(new_n544));
  NOR2_X1   g344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g345(.A(new_n542), .B1(new_n545), .B2(KEYINPUT6), .ZN(new_n546));
  NAND2_X1  g346(.A1(new_n546), .A2(G20), .ZN(new_n547));
  AND2_X1   g347(.A1(new_n381), .A2(new_n382), .ZN(new_n548));
  OAI211_X1 g348(.A(new_n541), .B(new_n547), .C1(new_n548), .C2(new_n245), .ZN(new_n549));
  AOI211_X1 g349(.A(new_n538), .B(new_n539), .C1(new_n549), .C2(new_n286), .ZN(new_n550));
  NAND2_X1  g350(.A1(new_n533), .A2(G200), .ZN(new_n551));
  NAND4_X1  g351(.A1(new_n534), .A2(new_n537), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  AOI21_X1  g352(.A(new_n539), .B1(new_n549), .B2(new_n286), .ZN(new_n553));
  INV_X1    g353(.A(new_n538), .ZN(new_n554));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g355(.A1(new_n533), .A2(new_n315), .ZN(new_n556));
  OAI211_X1 g356(.A(new_n555), .B(new_n556), .C1(G179), .C2(new_n533), .ZN(new_n557));
  NAND3_X1  g357(.A1(new_n472), .A2(G190), .A3(new_n475), .ZN(new_n558));
  NAND4_X1  g358(.A1(new_n454), .A2(new_n457), .A3(new_n459), .A4(new_n558), .ZN(new_n559));
  NOR2_X1   g359(.A1(new_n477), .A2(new_n322), .ZN(new_n560));
  OAI211_X1 g360(.A(new_n552), .B(new_n557), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  OAI211_X1 g361(.A(new_n526), .B(new_n204), .C1(G33), .C2(new_n489), .ZN(new_n562));
  INV_X1    g362(.A(KEYINPUT82), .ZN(new_n563));
  XNOR2_X1  g363(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND2_X1  g364(.A1(new_n207), .A2(G20), .ZN(new_n565));
  NAND3_X1  g365(.A1(new_n564), .A2(new_n286), .A3(new_n565), .ZN(new_n566));
  INV_X1    g366(.A(KEYINPUT20), .ZN(new_n567));
  XNOR2_X1  g367(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NOR2_X1   g368(.A1(new_n291), .A2(G116), .ZN(new_n569));
  INV_X1    g369(.A(new_n569), .ZN(new_n570));
  AOI22_X1  g370(.A1(new_n308), .A2(new_n310), .B1(new_n203), .B2(G33), .ZN(new_n571));
  NAND2_X1  g371(.A1(new_n571), .A2(G116), .ZN(new_n572));
  NAND3_X1  g372(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g373(.A(new_n368), .B1(G264), .B2(new_n461), .ZN(new_n574));
  NOR2_X1   g374(.A1(G257), .A2(G1698), .ZN(new_n575));
  INV_X1    g375(.A(G303), .ZN(new_n576));
  OAI22_X1  g376(.A1(new_n574), .A2(new_n575), .B1(new_n576), .B2(new_n256), .ZN(new_n577));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n265), .ZN(new_n578));
  NAND2_X1  g378(.A1(new_n471), .A2(G270), .ZN(new_n579));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n475), .ZN(new_n580));
  NAND3_X1  g380(.A1(new_n573), .A2(G169), .A3(new_n580), .ZN(new_n581));
  INV_X1    g381(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g383(.A1(new_n580), .A2(new_n275), .ZN(new_n584));
  NAND2_X1  g384(.A1(new_n573), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g385(.A1(new_n568), .A2(new_n570), .A3(new_n572), .ZN(new_n586));
  OR2_X1    g386(.A1(new_n580), .A2(new_n358), .ZN(new_n587));
  NAND2_X1  g387(.A1(new_n580), .A2(G200), .ZN(new_n588));
  NAND3_X1  g388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND4_X1  g389(.A1(new_n573), .A2(KEYINPUT21), .A3(G169), .A4(new_n580), .ZN(new_n590));
  NAND4_X1  g390(.A1(new_n583), .A2(new_n585), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NOR2_X1   g391(.A1(new_n561), .A2(new_n591), .ZN(new_n592));
  AND4_X1   g392(.A1(new_n434), .A2(new_n483), .A3(new_n522), .A4(new_n592), .ZN(G372));
  INV_X1    g393(.A(new_n293), .ZN(new_n594));
  NOR2_X1   g394(.A1(new_n325), .A2(new_n327), .ZN(new_n595));
  INV_X1    g395(.A(new_n427), .ZN(new_n596));
  AND3_X1   g396(.A1(new_n301), .A2(new_n313), .A3(new_n316), .ZN(new_n597));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n359), .ZN(new_n598));
  AOI21_X1  g398(.A(new_n596), .B1(new_n598), .B2(new_n355), .ZN(new_n599));
  NAND2_X1  g399(.A1(new_n413), .A2(new_n414), .ZN(new_n600));
  NAND2_X1  g400(.A1(new_n391), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g401(.A(new_n601), .B(KEYINPUT18), .ZN(new_n602));
  NOR2_X1   g402(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g403(.A(new_n595), .B1(new_n603), .B2(KEYINPUT85), .ZN(new_n604));
  INV_X1    g404(.A(KEYINPUT85), .ZN(new_n605));
  OAI21_X1  g405(.A(new_n605), .B1(new_n599), .B2(new_n602), .ZN(new_n606));
  AOI21_X1  g406(.A(new_n594), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  INV_X1    g407(.A(new_n557), .ZN(new_n608));
  INV_X1    g408(.A(KEYINPUT26), .ZN(new_n609));
  NAND2_X1  g409(.A1(new_n499), .A2(new_n510), .ZN(new_n610));
  NAND4_X1  g410(.A1(new_n608), .A2(new_n609), .A3(new_n521), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n610), .ZN(new_n612));
  INV_X1    g412(.A(new_n479), .ZN(new_n613));
  NAND3_X1  g413(.A1(new_n583), .A2(new_n585), .A3(new_n590), .ZN(new_n614));
  OR2_X1    g414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g415(.A1(new_n521), .A2(new_n610), .ZN(new_n616));
  NOR2_X1   g416(.A1(new_n561), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g417(.A(new_n612), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g418(.A1(new_n522), .A2(new_n608), .ZN(new_n619));
  NAND2_X1  g419(.A1(new_n619), .A2(KEYINPUT26), .ZN(new_n620));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g421(.A1(new_n434), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n622), .ZN(G369));
  INV_X1    g423(.A(G13), .ZN(new_n624));
  NOR2_X1   g424(.A1(new_n624), .A2(G20), .ZN(new_n625));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n203), .ZN(new_n626));
  OR2_X1    g426(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n627));
  NAND2_X1  g427(.A1(new_n626), .A2(KEYINPUT27), .ZN(new_n628));
  NAND3_X1  g428(.A1(new_n627), .A2(G213), .A3(new_n628), .ZN(new_n629));
  INV_X1    g429(.A(G343), .ZN(new_n630));
  NOR2_X1   g430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g431(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g432(.A1(new_n586), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g434(.A(new_n634), .B(KEYINPUT86), .Z(new_n635));
  OAI21_X1  g435(.A(new_n635), .B1(new_n591), .B2(new_n633), .ZN(new_n636));
  NAND2_X1  g436(.A1(new_n460), .A2(new_n631), .ZN(new_n637));
  OAI211_X1 g437(.A(new_n483), .B(new_n637), .C1(new_n560), .C2(new_n559), .ZN(new_n638));
  OAI21_X1  g438(.A(new_n638), .B1(new_n479), .B2(new_n632), .ZN(new_n639));
  NAND3_X1  g439(.A1(new_n636), .A2(G330), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g440(.A(new_n640), .B(KEYINPUT87), .ZN(new_n641));
  NAND2_X1  g441(.A1(new_n614), .A2(new_n632), .ZN(new_n642));
  XNOR2_X1  g442(.A(new_n642), .B(KEYINPUT88), .ZN(new_n643));
  AND2_X1   g443(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g444(.A(new_n644), .B1(new_n613), .B2(new_n632), .ZN(new_n645));
  NAND2_X1  g445(.A1(new_n641), .A2(new_n645), .ZN(G399));
  INV_X1    g446(.A(KEYINPUT89), .ZN(new_n647));
  INV_X1    g447(.A(new_n227), .ZN(new_n648));
  OAI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(G41), .ZN(new_n649));
  NAND3_X1  g449(.A1(new_n227), .A2(KEYINPUT89), .A3(new_n267), .ZN(new_n650));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g451(.A1(new_n651), .A2(G1), .ZN(new_n652));
  OR2_X1    g452(.A1(new_n485), .A2(G116), .ZN(new_n653));
  OAI22_X1  g453(.A1(new_n652), .A2(new_n653), .B1(new_n232), .B2(new_n651), .ZN(new_n654));
  XNOR2_X1  g454(.A(new_n654), .B(KEYINPUT28), .ZN(new_n655));
  NAND4_X1  g455(.A1(new_n592), .A2(new_n483), .A3(new_n522), .A4(new_n632), .ZN(new_n656));
  AND2_X1   g456(.A1(new_n472), .A2(new_n514), .ZN(new_n657));
  INV_X1    g457(.A(new_n533), .ZN(new_n658));
  NAND3_X1  g458(.A1(new_n584), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g459(.A(KEYINPUT30), .ZN(new_n660));
  NAND2_X1  g460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g461(.A1(new_n584), .A2(new_n657), .A3(new_n658), .A4(KEYINPUT30), .ZN(new_n662));
  AND2_X1   g462(.A1(new_n580), .A2(new_n508), .ZN(new_n663));
  NAND2_X1  g463(.A1(new_n472), .A2(new_n475), .ZN(new_n664));
  NAND4_X1  g464(.A1(new_n663), .A2(new_n275), .A3(new_n664), .A4(new_n533), .ZN(new_n665));
  NAND3_X1  g465(.A1(new_n661), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n631), .ZN(new_n667));
  INV_X1    g467(.A(KEYINPUT31), .ZN(new_n668));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g469(.A1(new_n666), .A2(KEYINPUT31), .A3(new_n631), .ZN(new_n670));
  NAND3_X1  g470(.A1(new_n656), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g471(.A(KEYINPUT90), .ZN(new_n672));
  AND3_X1   g472(.A1(new_n671), .A2(new_n672), .A3(G330), .ZN(new_n673));
  AOI21_X1  g473(.A(new_n672), .B1(new_n671), .B2(G330), .ZN(new_n674));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g475(.A(new_n483), .ZN(new_n676));
  OAI21_X1  g476(.A(new_n617), .B1(new_n676), .B2(new_n614), .ZN(new_n677));
  NAND3_X1  g477(.A1(new_n522), .A2(new_n609), .A3(new_n608), .ZN(new_n678));
  OAI21_X1  g478(.A(KEYINPUT26), .B1(new_n616), .B2(new_n557), .ZN(new_n679));
  AND2_X1   g479(.A1(new_n679), .A2(new_n610), .ZN(new_n680));
  NAND3_X1  g480(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g481(.A1(new_n681), .A2(KEYINPUT29), .A3(new_n632), .ZN(new_n682));
  AOI21_X1  g482(.A(new_n631), .B1(new_n618), .B2(new_n620), .ZN(new_n683));
  OAI21_X1  g483(.A(new_n682), .B1(KEYINPUT29), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g484(.A1(new_n675), .A2(new_n684), .ZN(new_n685));
  INV_X1    g485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g486(.A(new_n655), .B1(new_n686), .B2(G1), .ZN(G364));
  NOR2_X1   g487(.A1(G13), .A2(G33), .ZN(new_n688));
  INV_X1    g488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g489(.A1(new_n689), .A2(G20), .ZN(new_n690));
  INV_X1    g490(.A(new_n690), .ZN(new_n691));
  OR2_X1    g491(.A1(new_n636), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g492(.A(new_n204), .B1(KEYINPUT92), .B2(new_n315), .ZN(new_n693));
  OAI21_X1  g493(.A(new_n693), .B1(KEYINPUT92), .B2(new_n315), .ZN(new_n694));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n284), .ZN(new_n695));
  INV_X1    g495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g496(.A1(new_n204), .A2(new_n358), .ZN(new_n697));
  NAND3_X1  g497(.A1(new_n697), .A2(G179), .A3(new_n322), .ZN(new_n698));
  INV_X1    g498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g499(.A1(new_n204), .A2(G190), .ZN(new_n700));
  NOR2_X1   g500(.A1(G179), .A2(G200), .ZN(new_n701));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g502(.A(new_n702), .ZN(new_n703));
  AOI22_X1  g503(.A1(new_n699), .A2(G322), .B1(new_n703), .B2(G329), .ZN(new_n704));
  AOI21_X1  g504(.A(new_n204), .B1(new_n701), .B2(G190), .ZN(new_n705));
  NOR2_X1   g505(.A1(new_n322), .A2(G179), .ZN(new_n706));
  NAND2_X1  g506(.A1(new_n697), .A2(new_n706), .ZN(new_n707));
  OAI221_X1 g507(.A(new_n704), .B1(new_n464), .B2(new_n705), .C1(new_n576), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g508(.A1(new_n700), .A2(new_n706), .ZN(new_n709));
  INV_X1    g509(.A(G283), .ZN(new_n710));
  NOR2_X1   g510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g511(.A(new_n700), .ZN(new_n712));
  NOR3_X1   g512(.A1(new_n712), .A2(new_n275), .A3(G200), .ZN(new_n713));
  AND2_X1   g513(.A1(new_n713), .A2(G311), .ZN(new_n714));
  NOR4_X1   g514(.A1(new_n708), .A2(new_n256), .A3(new_n711), .A4(new_n714), .ZN(new_n715));
  INV_X1    g515(.A(G326), .ZN(new_n716));
  NOR2_X1   g516(.A1(new_n275), .A2(new_n322), .ZN(new_n717));
  NAND2_X1  g517(.A1(new_n697), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n700), .ZN(new_n719));
  XNOR2_X1  g519(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n720));
  XNOR2_X1  g520(.A(new_n720), .B(G317), .ZN(new_n721));
  OAI221_X1 g521(.A(new_n715), .B1(new_n716), .B2(new_n718), .C1(new_n719), .C2(new_n721), .ZN(new_n722));
  XOR2_X1   g522(.A(new_n722), .B(KEYINPUT96), .Z(new_n723));
  OR2_X1    g523(.A1(new_n713), .A2(KEYINPUT93), .ZN(new_n724));
  NAND2_X1  g524(.A1(new_n713), .A2(KEYINPUT93), .ZN(new_n725));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI22_X1  g526(.A1(new_n726), .A2(new_n219), .B1(new_n222), .B2(new_n698), .ZN(new_n727));
  INV_X1    g527(.A(KEYINPUT94), .ZN(new_n728));
  OR2_X1    g528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g529(.A(new_n707), .ZN(new_n730));
  NAND2_X1  g530(.A1(new_n730), .A2(G87), .ZN(new_n731));
  NOR2_X1   g531(.A1(new_n705), .A2(new_n489), .ZN(new_n732));
  OAI22_X1  g532(.A1(new_n718), .A2(new_n217), .B1(new_n719), .B2(new_n211), .ZN(new_n733));
  NAND2_X1  g533(.A1(new_n703), .A2(G159), .ZN(new_n734));
  AOI211_X1 g534(.A(new_n732), .B(new_n733), .C1(KEYINPUT32), .C2(new_n734), .ZN(new_n735));
  NAND3_X1  g535(.A1(new_n729), .A2(new_n731), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g536(.A1(new_n727), .A2(new_n728), .ZN(new_n737));
  OAI21_X1  g537(.A(new_n737), .B1(new_n245), .B2(new_n709), .ZN(new_n738));
  NOR2_X1   g538(.A1(new_n734), .A2(KEYINPUT32), .ZN(new_n739));
  NOR4_X1   g539(.A1(new_n736), .A2(new_n738), .A3(new_n260), .A4(new_n739), .ZN(new_n740));
  OAI21_X1  g540(.A(new_n696), .B1(new_n723), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g541(.A(new_n652), .B1(G45), .B2(new_n625), .ZN(new_n742));
  NAND2_X1  g542(.A1(new_n250), .A2(G45), .ZN(new_n743));
  NOR2_X1   g543(.A1(new_n648), .A2(new_n368), .ZN(new_n744));
  OAI211_X1 g544(.A(new_n743), .B(new_n744), .C1(G45), .C2(new_n232), .ZN(new_n745));
  NAND3_X1  g545(.A1(new_n227), .A2(G355), .A3(new_n256), .ZN(new_n746));
  OAI211_X1 g546(.A(new_n745), .B(new_n746), .C1(G116), .C2(new_n227), .ZN(new_n747));
  XOR2_X1   g547(.A(new_n747), .B(KEYINPUT91), .Z(new_n748));
  NOR2_X1   g548(.A1(new_n696), .A2(new_n690), .ZN(new_n749));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g550(.A1(new_n692), .A2(new_n741), .A3(new_n742), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g551(.A1(new_n636), .A2(G330), .ZN(new_n752));
  NAND2_X1  g552(.A1(new_n636), .A2(G330), .ZN(new_n753));
  INV_X1    g553(.A(new_n742), .ZN(new_n754));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g555(.A(new_n751), .B1(new_n752), .B2(new_n755), .ZN(G396));
  NAND2_X1  g556(.A1(new_n313), .A2(new_n631), .ZN(new_n757));
  INV_X1    g557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g558(.A(new_n317), .B1(new_n433), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g559(.A1(new_n317), .A2(new_n631), .ZN(new_n760));
  INV_X1    g560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g562(.A1(new_n675), .A2(new_n762), .ZN(new_n763));
  INV_X1    g563(.A(new_n762), .ZN(new_n764));
  OAI21_X1  g564(.A(new_n764), .B1(new_n673), .B2(new_n674), .ZN(new_n765));
  NAND2_X1  g565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g566(.A(new_n766), .B(new_n683), .Z(new_n767));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n742), .ZN(new_n768));
  NOR2_X1   g568(.A1(new_n764), .A2(new_n689), .ZN(new_n769));
  INV_X1    g569(.A(G132), .ZN(new_n770));
  OAI21_X1  g570(.A(new_n368), .B1(new_n770), .B2(new_n702), .ZN(new_n771));
  INV_X1    g571(.A(new_n719), .ZN(new_n772));
  AOI22_X1  g572(.A1(new_n699), .A2(G143), .B1(new_n772), .B2(G150), .ZN(new_n773));
  INV_X1    g573(.A(G137), .ZN(new_n774));
  INV_X1    g574(.A(G159), .ZN(new_n775));
  OAI221_X1 g575(.A(new_n773), .B1(new_n774), .B2(new_n718), .C1(new_n726), .C2(new_n775), .ZN(new_n776));
  XOR2_X1   g576(.A(new_n776), .B(KEYINPUT34), .Z(new_n777));
  INV_X1    g577(.A(new_n709), .ZN(new_n778));
  AOI211_X1 g578(.A(new_n771), .B(new_n777), .C1(G68), .C2(new_n778), .ZN(new_n779));
  OAI221_X1 g579(.A(new_n779), .B1(new_n217), .B2(new_n707), .C1(new_n222), .C2(new_n705), .ZN(new_n780));
  AOI21_X1  g580(.A(new_n732), .B1(G294), .B2(new_n699), .ZN(new_n781));
  XOR2_X1   g581(.A(new_n781), .B(KEYINPUT97), .Z(new_n782));
  INV_X1    g582(.A(new_n726), .ZN(new_n783));
  AOI211_X1 g583(.A(new_n256), .B(new_n782), .C1(G116), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g584(.A1(new_n703), .A2(G311), .ZN(new_n785));
  NAND2_X1  g585(.A1(new_n778), .A2(G87), .ZN(new_n786));
  OAI22_X1  g586(.A1(new_n718), .A2(new_n576), .B1(new_n719), .B2(new_n710), .ZN(new_n787));
  AOI21_X1  g587(.A(new_n787), .B1(G107), .B2(new_n730), .ZN(new_n788));
  NAND4_X1  g588(.A1(new_n784), .A2(new_n785), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g589(.A(new_n695), .B1(new_n780), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g590(.A1(new_n696), .A2(G77), .A3(new_n688), .ZN(new_n791));
  NOR4_X1   g591(.A1(new_n769), .A2(new_n790), .A3(new_n754), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g592(.A1(new_n768), .A2(new_n792), .ZN(new_n793));
  INV_X1    g593(.A(new_n793), .ZN(G384));
  NAND3_X1  g594(.A1(new_n378), .A2(new_n286), .A3(new_n386), .ZN(new_n795));
  AOI21_X1  g595(.A(KEYINPUT16), .B1(new_n370), .B2(new_n376), .ZN(new_n796));
  OAI21_X1  g596(.A(new_n390), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g597(.A(new_n629), .ZN(new_n798));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g600(.A1(new_n430), .A2(new_n800), .ZN(new_n801));
  INV_X1    g601(.A(KEYINPUT37), .ZN(new_n802));
  NAND3_X1  g602(.A1(new_n387), .A2(new_n390), .A3(new_n421), .ZN(new_n803));
  NAND2_X1  g603(.A1(new_n391), .A2(new_n798), .ZN(new_n804));
  NAND4_X1  g604(.A1(new_n416), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g605(.A1(new_n797), .A2(new_n600), .ZN(new_n806));
  AND3_X1   g606(.A1(new_n799), .A2(new_n806), .A3(new_n803), .ZN(new_n807));
  OAI21_X1  g607(.A(new_n805), .B1(new_n807), .B2(new_n802), .ZN(new_n808));
  AND3_X1   g608(.A1(new_n801), .A2(new_n808), .A3(KEYINPUT38), .ZN(new_n809));
  NAND2_X1  g609(.A1(new_n805), .A2(KEYINPUT100), .ZN(new_n810));
  NAND3_X1  g610(.A1(new_n601), .A2(new_n804), .A3(new_n803), .ZN(new_n811));
  NAND2_X1  g611(.A1(new_n811), .A2(KEYINPUT37), .ZN(new_n812));
  AOI21_X1  g612(.A(new_n629), .B1(new_n387), .B2(new_n390), .ZN(new_n813));
  NOR2_X1   g613(.A1(new_n425), .A2(new_n813), .ZN(new_n814));
  INV_X1    g614(.A(KEYINPUT100), .ZN(new_n815));
  NAND4_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n802), .A4(new_n416), .ZN(new_n816));
  NAND3_X1  g616(.A1(new_n810), .A2(new_n812), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g617(.A1(new_n817), .A2(KEYINPUT101), .ZN(new_n818));
  OAI21_X1  g618(.A(new_n813), .B1(new_n602), .B2(new_n596), .ZN(new_n819));
  INV_X1    g619(.A(KEYINPUT101), .ZN(new_n820));
  NAND4_X1  g620(.A1(new_n810), .A2(new_n820), .A3(new_n812), .A4(new_n816), .ZN(new_n821));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  INV_X1    g622(.A(KEYINPUT38), .ZN(new_n823));
  AOI21_X1  g623(.A(new_n809), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g624(.A(new_n824), .ZN(new_n825));
  OAI211_X1 g625(.A(new_n355), .B(new_n359), .C1(new_n357), .C2(new_n632), .ZN(new_n826));
  NAND3_X1  g626(.A1(new_n343), .A2(new_n354), .A3(new_n631), .ZN(new_n827));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g628(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n762), .ZN(new_n830));
  INV_X1    g630(.A(KEYINPUT105), .ZN(new_n831));
  XNOR2_X1  g631(.A(new_n670), .B(new_n831), .ZN(new_n832));
  INV_X1    g632(.A(KEYINPUT104), .ZN(new_n833));
  NAND2_X1  g633(.A1(new_n669), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g634(.A1(new_n667), .A2(KEYINPUT104), .A3(new_n668), .ZN(new_n835));
  NAND4_X1  g635(.A1(new_n832), .A2(new_n656), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  NAND4_X1  g636(.A1(new_n825), .A2(KEYINPUT40), .A3(new_n830), .A4(new_n836), .ZN(new_n837));
  INV_X1    g637(.A(KEYINPUT40), .ZN(new_n838));
  NAND2_X1  g638(.A1(new_n830), .A2(new_n836), .ZN(new_n839));
  AOI21_X1  g639(.A(KEYINPUT38), .B1(new_n801), .B2(new_n808), .ZN(new_n840));
  NOR2_X1   g640(.A1(new_n809), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g641(.A(new_n838), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g642(.A1(new_n837), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g643(.A1(new_n843), .A2(G330), .ZN(new_n844));
  AND2_X1   g644(.A1(new_n836), .A2(G330), .ZN(new_n845));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n434), .ZN(new_n846));
  NAND2_X1  g646(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g647(.A1(new_n843), .A2(new_n434), .A3(new_n836), .ZN(new_n848));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g649(.A(new_n434), .B(new_n682), .C1(KEYINPUT29), .C2(new_n683), .ZN(new_n850));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n607), .ZN(new_n851));
  XNOR2_X1  g651(.A(new_n851), .B(KEYINPUT103), .ZN(new_n852));
  XNOR2_X1  g652(.A(new_n849), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g653(.A1(new_n822), .A2(new_n823), .ZN(new_n854));
  INV_X1    g654(.A(KEYINPUT39), .ZN(new_n855));
  INV_X1    g655(.A(new_n809), .ZN(new_n856));
  NAND3_X1  g656(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g657(.A(KEYINPUT102), .ZN(new_n858));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g659(.A1(new_n824), .A2(KEYINPUT102), .A3(new_n855), .ZN(new_n860));
  INV_X1    g660(.A(KEYINPUT99), .ZN(new_n861));
  OAI21_X1  g661(.A(new_n861), .B1(new_n841), .B2(new_n855), .ZN(new_n862));
  OAI211_X1 g662(.A(KEYINPUT99), .B(KEYINPUT39), .C1(new_n809), .C2(new_n840), .ZN(new_n863));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g664(.A1(new_n859), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g665(.A1(new_n355), .A2(new_n631), .ZN(new_n866));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g667(.A(new_n760), .B1(new_n683), .B2(new_n759), .ZN(new_n868));
  NOR3_X1   g668(.A1(new_n868), .A2(new_n841), .A3(new_n829), .ZN(new_n869));
  AOI21_X1  g669(.A(new_n869), .B1(new_n602), .B2(new_n629), .ZN(new_n870));
  NAND2_X1  g670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g671(.A(new_n853), .B(new_n871), .ZN(new_n872));
  OAI21_X1  g672(.A(new_n872), .B1(new_n203), .B2(new_n625), .ZN(new_n873));
  OAI21_X1  g673(.A(G77), .B1(new_n222), .B2(new_n211), .ZN(new_n874));
  OAI22_X1  g674(.A1(new_n232), .A2(new_n874), .B1(G50), .B2(new_n211), .ZN(new_n875));
  NAND3_X1  g675(.A1(new_n875), .A2(G1), .A3(new_n624), .ZN(new_n876));
  OAI211_X1 g676(.A(G20), .B(new_n284), .C1(new_n546), .C2(KEYINPUT35), .ZN(new_n877));
  AOI211_X1 g677(.A(new_n207), .B(new_n877), .C1(KEYINPUT35), .C2(new_n546), .ZN(new_n878));
  XNOR2_X1  g678(.A(KEYINPUT98), .B(KEYINPUT36), .ZN(new_n879));
  XNOR2_X1  g679(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND3_X1  g680(.A1(new_n873), .A2(new_n876), .A3(new_n880), .ZN(G367));
  INV_X1    g681(.A(KEYINPUT42), .ZN(new_n882));
  AOI22_X1  g682(.A1(new_n644), .A2(new_n882), .B1(new_n676), .B2(new_n632), .ZN(new_n883));
  OAI21_X1  g683(.A(new_n552), .B1(new_n550), .B2(new_n632), .ZN(new_n884));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n557), .ZN(new_n885));
  INV_X1    g685(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g687(.A1(new_n557), .A2(new_n631), .ZN(new_n888));
  AOI21_X1  g688(.A(new_n882), .B1(new_n644), .B2(new_n885), .ZN(new_n889));
  NOR3_X1   g689(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g690(.A(new_n632), .B1(new_n513), .B2(new_n519), .ZN(new_n891));
  MUX2_X1   g691(.A(new_n616), .B(new_n610), .S(new_n891), .Z(new_n892));
  INV_X1    g692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g693(.A(new_n890), .B1(KEYINPUT43), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g694(.A1(new_n886), .A2(new_n888), .ZN(new_n895));
  INV_X1    g695(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g696(.A1(new_n641), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g697(.A(new_n894), .B(new_n897), .ZN(new_n898));
  NOR2_X1   g698(.A1(new_n893), .A2(KEYINPUT43), .ZN(new_n899));
  XOR2_X1   g699(.A(new_n898), .B(new_n899), .Z(new_n900));
  XOR2_X1   g700(.A(new_n651), .B(KEYINPUT106), .Z(new_n901));
  XOR2_X1   g701(.A(new_n901), .B(KEYINPUT41), .Z(new_n902));
  INV_X1    g702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g703(.A1(new_n645), .A2(new_n895), .ZN(new_n904));
  XOR2_X1   g704(.A(new_n904), .B(KEYINPUT45), .Z(new_n905));
  OAI211_X1 g705(.A(KEYINPUT107), .B(KEYINPUT44), .C1(new_n645), .C2(new_n895), .ZN(new_n906));
  XNOR2_X1  g706(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n907));
  OR3_X1    g707(.A1(new_n645), .A2(new_n895), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g708(.A1(new_n905), .A2(new_n906), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g709(.A1(new_n641), .A2(KEYINPUT108), .ZN(new_n910));
  OR2_X1    g710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n910), .ZN(new_n912));
  XNOR2_X1  g712(.A(new_n753), .B(new_n639), .ZN(new_n913));
  XNOR2_X1  g713(.A(new_n913), .B(new_n643), .ZN(new_n914));
  INV_X1    g714(.A(new_n914), .ZN(new_n915));
  NAND4_X1  g715(.A1(new_n911), .A2(new_n686), .A3(new_n912), .A4(new_n915), .ZN(new_n916));
  AOI21_X1  g716(.A(new_n903), .B1(new_n916), .B2(new_n686), .ZN(new_n917));
  AOI21_X1  g717(.A(new_n203), .B1(new_n625), .B2(G45), .ZN(new_n918));
  INV_X1    g718(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g719(.A(new_n900), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g720(.A1(new_n707), .A2(new_n222), .ZN(new_n921));
  AOI22_X1  g721(.A1(G159), .A2(new_n772), .B1(new_n703), .B2(G137), .ZN(new_n922));
  NAND2_X1  g722(.A1(new_n778), .A2(G77), .ZN(new_n923));
  OAI211_X1 g723(.A(new_n922), .B(new_n923), .C1(new_n278), .C2(new_n698), .ZN(new_n924));
  INV_X1    g724(.A(new_n718), .ZN(new_n925));
  AOI211_X1 g725(.A(new_n921), .B(new_n924), .C1(G143), .C2(new_n925), .ZN(new_n926));
  INV_X1    g726(.A(new_n705), .ZN(new_n927));
  NAND2_X1  g727(.A1(new_n927), .A2(G68), .ZN(new_n928));
  NAND2_X1  g728(.A1(new_n783), .A2(G50), .ZN(new_n929));
  NAND4_X1  g729(.A1(new_n926), .A2(new_n256), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  AOI21_X1  g730(.A(KEYINPUT46), .B1(new_n730), .B2(G116), .ZN(new_n931));
  NAND3_X1  g731(.A1(new_n730), .A2(KEYINPUT46), .A3(G116), .ZN(new_n932));
  XOR2_X1   g732(.A(new_n932), .B(KEYINPUT109), .Z(new_n933));
  AOI211_X1 g733(.A(new_n931), .B(new_n933), .C1(G294), .C2(new_n772), .ZN(new_n934));
  INV_X1    g734(.A(KEYINPUT110), .ZN(new_n935));
  NAND2_X1  g735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g736(.A1(new_n778), .A2(G97), .ZN(new_n937));
  NAND2_X1  g737(.A1(new_n703), .A2(G317), .ZN(new_n938));
  AOI22_X1  g738(.A1(new_n699), .A2(G303), .B1(new_n927), .B2(G107), .ZN(new_n939));
  NAND2_X1  g739(.A1(new_n925), .A2(G311), .ZN(new_n940));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n365), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g741(.A(new_n941), .B1(new_n783), .B2(G283), .ZN(new_n942));
  NAND4_X1  g742(.A1(new_n936), .A2(new_n937), .A3(new_n938), .A4(new_n942), .ZN(new_n943));
  NOR2_X1   g743(.A1(new_n934), .A2(new_n935), .ZN(new_n944));
  OAI21_X1  g744(.A(new_n930), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g745(.A(new_n945), .B(KEYINPUT47), .ZN(new_n946));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n696), .ZN(new_n947));
  NAND2_X1  g747(.A1(new_n892), .A2(new_n690), .ZN(new_n948));
  INV_X1    g748(.A(new_n744), .ZN(new_n949));
  OAI221_X1 g749(.A(new_n749), .B1(new_n227), .B2(new_n305), .C1(new_n242), .C2(new_n949), .ZN(new_n950));
  NAND4_X1  g750(.A1(new_n947), .A2(new_n742), .A3(new_n948), .A4(new_n950), .ZN(new_n951));
  NAND2_X1  g751(.A1(new_n920), .A2(new_n951), .ZN(G387));
  NAND2_X1  g752(.A1(new_n915), .A2(new_n686), .ZN(new_n953));
  INV_X1    g753(.A(new_n651), .ZN(new_n954));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g755(.A(new_n955), .B(KEYINPUT112), .ZN(new_n956));
  OAI21_X1  g756(.A(new_n956), .B1(new_n686), .B2(new_n915), .ZN(new_n957));
  NAND2_X1  g757(.A1(new_n915), .A2(new_n919), .ZN(new_n958));
  NOR2_X1   g758(.A1(new_n702), .A2(new_n278), .ZN(new_n959));
  AOI22_X1  g759(.A1(new_n713), .A2(G68), .B1(new_n925), .B2(G159), .ZN(new_n960));
  NAND2_X1  g760(.A1(new_n730), .A2(G77), .ZN(new_n961));
  NAND2_X1  g761(.A1(new_n927), .A2(new_n304), .ZN(new_n962));
  NAND3_X1  g762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g763(.A(new_n368), .B1(new_n217), .B2(new_n698), .ZN(new_n964));
  OAI21_X1  g764(.A(new_n937), .B1(new_n282), .B2(new_n719), .ZN(new_n965));
  OR4_X1    g765(.A1(new_n959), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  AOI22_X1  g766(.A1(new_n699), .A2(G317), .B1(new_n772), .B2(G311), .ZN(new_n967));
  INV_X1    g767(.A(G322), .ZN(new_n968));
  OAI221_X1 g768(.A(new_n967), .B1(new_n968), .B2(new_n718), .C1(new_n726), .C2(new_n576), .ZN(new_n969));
  XNOR2_X1  g769(.A(new_n969), .B(KEYINPUT48), .ZN(new_n970));
  OAI221_X1 g770(.A(new_n970), .B1(new_n710), .B2(new_n705), .C1(new_n464), .C2(new_n707), .ZN(new_n971));
  XOR2_X1   g771(.A(new_n971), .B(KEYINPUT49), .Z(new_n972));
  OAI221_X1 g772(.A(new_n365), .B1(new_n207), .B2(new_n709), .C1(new_n716), .C2(new_n702), .ZN(new_n973));
  OAI21_X1  g773(.A(new_n966), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g774(.A(new_n974), .B(KEYINPUT111), .ZN(new_n975));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n696), .ZN(new_n976));
  OR2_X1    g776(.A1(new_n639), .A2(new_n691), .ZN(new_n977));
  NAND2_X1  g777(.A1(new_n388), .A2(new_n217), .ZN(new_n978));
  XNOR2_X1  g778(.A(new_n978), .B(KEYINPUT50), .ZN(new_n979));
  NOR2_X1   g779(.A1(new_n211), .A2(new_n219), .ZN(new_n980));
  NOR4_X1   g780(.A1(new_n979), .A2(new_n653), .A3(G45), .A4(new_n980), .ZN(new_n981));
  OAI21_X1  g781(.A(new_n744), .B1(new_n239), .B2(new_n268), .ZN(new_n982));
  NAND3_X1  g782(.A1(new_n653), .A2(new_n227), .A3(new_n256), .ZN(new_n983));
  AOI21_X1  g783(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g784(.A1(new_n227), .A2(G107), .ZN(new_n985));
  OAI21_X1  g785(.A(new_n749), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND4_X1  g786(.A1(new_n976), .A2(new_n742), .A3(new_n977), .A4(new_n986), .ZN(new_n987));
  NAND3_X1  g787(.A1(new_n957), .A2(new_n958), .A3(new_n987), .ZN(G393));
  INV_X1    g788(.A(new_n641), .ZN(new_n989));
  XNOR2_X1  g789(.A(new_n909), .B(new_n989), .ZN(new_n990));
  NAND2_X1  g790(.A1(new_n990), .A2(new_n953), .ZN(new_n991));
  NAND2_X1  g791(.A1(new_n991), .A2(KEYINPUT114), .ZN(new_n992));
  INV_X1    g792(.A(KEYINPUT114), .ZN(new_n993));
  NAND3_X1  g793(.A1(new_n990), .A2(new_n993), .A3(new_n953), .ZN(new_n994));
  NAND4_X1  g794(.A1(new_n992), .A2(new_n954), .A3(new_n916), .A4(new_n994), .ZN(new_n995));
  OR2_X1    g795(.A1(new_n990), .A2(new_n918), .ZN(new_n996));
  NAND2_X1  g796(.A1(new_n896), .A2(new_n690), .ZN(new_n997));
  AOI22_X1  g797(.A1(new_n699), .A2(G311), .B1(new_n925), .B2(G317), .ZN(new_n998));
  XNOR2_X1  g798(.A(new_n998), .B(KEYINPUT113), .ZN(new_n999));
  XNOR2_X1  g799(.A(new_n999), .B(KEYINPUT52), .ZN(new_n1000));
  NAND2_X1  g800(.A1(new_n713), .A2(G294), .ZN(new_n1001));
  AOI21_X1  g801(.A(new_n256), .B1(new_n778), .B2(G107), .ZN(new_n1002));
  OAI22_X1  g802(.A1(new_n719), .A2(new_n576), .B1(new_n702), .B2(new_n968), .ZN(new_n1003));
  AOI21_X1  g803(.A(new_n1003), .B1(G283), .B2(new_n730), .ZN(new_n1004));
  NAND4_X1  g804(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g805(.A(new_n1005), .B1(G116), .B2(new_n927), .ZN(new_n1006));
  OAI22_X1  g806(.A1(new_n698), .A2(new_n775), .B1(new_n718), .B2(new_n278), .ZN(new_n1007));
  XOR2_X1   g807(.A(new_n1007), .B(KEYINPUT51), .Z(new_n1008));
  AOI21_X1  g808(.A(new_n1008), .B1(G143), .B2(new_n703), .ZN(new_n1009));
  NAND2_X1  g809(.A1(new_n783), .A2(new_n388), .ZN(new_n1010));
  OAI221_X1 g810(.A(new_n368), .B1(new_n707), .B2(new_n211), .C1(new_n217), .C2(new_n719), .ZN(new_n1011));
  AOI21_X1  g811(.A(new_n1011), .B1(G77), .B2(new_n927), .ZN(new_n1012));
  AND4_X1   g812(.A1(new_n786), .A2(new_n1009), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1013));
  OAI21_X1  g813(.A(new_n696), .B1(new_n1006), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g814(.A1(new_n247), .A2(new_n744), .ZN(new_n1015));
  OAI211_X1 g815(.A(new_n1015), .B(new_n749), .C1(new_n489), .C2(new_n227), .ZN(new_n1016));
  NAND4_X1  g816(.A1(new_n997), .A2(new_n742), .A3(new_n1014), .A4(new_n1016), .ZN(new_n1017));
  NAND3_X1  g817(.A1(new_n995), .A2(new_n996), .A3(new_n1017), .ZN(G390));
  OAI22_X1  g818(.A1(new_n719), .A2(new_n774), .B1(new_n705), .B2(new_n775), .ZN(new_n1019));
  XOR2_X1   g819(.A(KEYINPUT54), .B(G143), .Z(new_n1020));
  AOI21_X1  g820(.A(new_n1019), .B1(new_n783), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g821(.A(new_n1021), .B(KEYINPUT118), .ZN(new_n1022));
  INV_X1    g822(.A(G128), .ZN(new_n1023));
  INV_X1    g823(.A(G125), .ZN(new_n1024));
  OAI22_X1  g824(.A1(new_n718), .A2(new_n1023), .B1(new_n702), .B2(new_n1024), .ZN(new_n1025));
  NOR3_X1   g825(.A1(new_n707), .A2(KEYINPUT53), .A3(new_n278), .ZN(new_n1026));
  NOR4_X1   g826(.A1(new_n1022), .A2(new_n260), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  OAI21_X1  g827(.A(KEYINPUT53), .B1(new_n707), .B2(new_n278), .ZN(new_n1028));
  NAND2_X1  g828(.A1(new_n778), .A2(G50), .ZN(new_n1029));
  NAND2_X1  g829(.A1(new_n699), .A2(G132), .ZN(new_n1030));
  NAND4_X1  g830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  OAI221_X1 g831(.A(new_n731), .B1(new_n219), .B2(new_n705), .C1(new_n464), .C2(new_n702), .ZN(new_n1032));
  OAI22_X1  g832(.A1(new_n698), .A2(new_n207), .B1(new_n709), .B2(new_n211), .ZN(new_n1033));
  OAI21_X1  g833(.A(new_n260), .B1(new_n718), .B2(new_n710), .ZN(new_n1034));
  NOR3_X1   g834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OAI221_X1 g835(.A(new_n1035), .B1(new_n489), .B2(new_n726), .C1(new_n245), .C2(new_n719), .ZN(new_n1036));
  AOI21_X1  g836(.A(new_n695), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g837(.A1(new_n696), .A2(new_n688), .ZN(new_n1038));
  AOI211_X1 g838(.A(new_n754), .B(new_n1037), .C1(new_n282), .C2(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g839(.A(new_n1039), .B(KEYINPUT119), .ZN(new_n1040));
  OAI21_X1  g840(.A(new_n1040), .B1(new_n865), .B2(new_n689), .ZN(new_n1041));
  XNOR2_X1  g841(.A(new_n1041), .B(KEYINPUT120), .ZN(new_n1042));
  INV_X1    g842(.A(new_n866), .ZN(new_n1043));
  OAI21_X1  g843(.A(new_n1043), .B1(new_n868), .B2(new_n829), .ZN(new_n1044));
  NAND4_X1  g844(.A1(new_n859), .A2(new_n860), .A3(new_n864), .A4(new_n1044), .ZN(new_n1045));
  AND2_X1   g845(.A1(new_n681), .A2(new_n632), .ZN(new_n1046));
  AOI21_X1  g846(.A(new_n760), .B1(new_n1046), .B2(new_n759), .ZN(new_n1047));
  OAI211_X1 g847(.A(new_n1043), .B(new_n825), .C1(new_n1047), .C2(new_n829), .ZN(new_n1048));
  NAND2_X1  g848(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  AND3_X1   g849(.A1(new_n830), .A2(new_n836), .A3(G330), .ZN(new_n1050));
  NAND2_X1  g850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g851(.A1(new_n1051), .A2(KEYINPUT115), .ZN(new_n1052));
  OAI211_X1 g852(.A(new_n764), .B(new_n828), .C1(new_n673), .C2(new_n674), .ZN(new_n1053));
  NAND3_X1  g853(.A1(new_n1045), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g854(.A(KEYINPUT115), .ZN(new_n1055));
  NAND3_X1  g855(.A1(new_n1049), .A2(new_n1055), .A3(new_n1050), .ZN(new_n1056));
  NAND3_X1  g856(.A1(new_n1052), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  OAI21_X1  g857(.A(new_n1042), .B1(new_n1057), .B2(new_n918), .ZN(new_n1058));
  NAND3_X1  g858(.A1(new_n836), .A2(G330), .A3(new_n764), .ZN(new_n1059));
  NAND2_X1  g859(.A1(new_n1059), .A2(new_n829), .ZN(new_n1060));
  NAND3_X1  g860(.A1(new_n1053), .A2(new_n1047), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g861(.A(new_n1050), .B1(new_n765), .B2(new_n829), .ZN(new_n1062));
  OAI21_X1  g862(.A(new_n1061), .B1(new_n1062), .B2(new_n868), .ZN(new_n1063));
  INV_X1    g863(.A(KEYINPUT116), .ZN(new_n1064));
  NAND2_X1  g864(.A1(new_n846), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g865(.A1(new_n845), .A2(KEYINPUT116), .A3(new_n434), .ZN(new_n1066));
  AOI21_X1  g866(.A(new_n851), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g867(.A(KEYINPUT117), .ZN(new_n1068));
  AND3_X1   g868(.A1(new_n1063), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g869(.A(new_n1068), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1070));
  NOR2_X1   g870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g871(.A1(new_n1057), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g872(.A1(new_n1072), .A2(new_n651), .ZN(new_n1073));
  NAND2_X1  g873(.A1(new_n1057), .A2(new_n1071), .ZN(new_n1074));
  AOI21_X1  g874(.A(new_n1058), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g875(.A(new_n1075), .ZN(G378));
  OAI21_X1  g876(.A(new_n1067), .B1(new_n1057), .B2(new_n1071), .ZN(new_n1077));
  INV_X1    g877(.A(KEYINPUT122), .ZN(new_n1078));
  NAND2_X1  g878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g879(.A1(new_n595), .A2(new_n594), .ZN(new_n1080));
  XOR2_X1   g880(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1081));
  XNOR2_X1  g881(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  NAND2_X1  g882(.A1(new_n292), .A2(new_n798), .ZN(new_n1083));
  XNOR2_X1  g883(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  NAND2_X1  g884(.A1(new_n844), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g885(.A(new_n1084), .ZN(new_n1086));
  NAND3_X1  g886(.A1(new_n1086), .A2(G330), .A3(new_n843), .ZN(new_n1087));
  NAND2_X1  g887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g888(.A(new_n871), .ZN(new_n1089));
  XNOR2_X1  g889(.A(new_n1088), .B(new_n1089), .ZN(new_n1090));
  OAI211_X1 g890(.A(KEYINPUT122), .B(new_n1067), .C1(new_n1057), .C2(new_n1071), .ZN(new_n1091));
  NAND3_X1  g891(.A1(new_n1079), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g892(.A(KEYINPUT57), .ZN(new_n1093));
  NAND2_X1  g893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g894(.A1(new_n1079), .A2(KEYINPUT57), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1095));
  NAND3_X1  g895(.A1(new_n1094), .A2(new_n954), .A3(new_n1095), .ZN(new_n1096));
  AOI22_X1  g896(.A1(new_n1086), .A2(new_n688), .B1(new_n217), .B2(new_n1038), .ZN(new_n1097));
  AOI21_X1  g897(.A(G41), .B1(new_n925), .B2(G116), .ZN(new_n1098));
  NAND3_X1  g898(.A1(new_n1098), .A2(new_n365), .A3(new_n961), .ZN(new_n1099));
  OAI221_X1 g899(.A(new_n928), .B1(new_n222), .B2(new_n709), .C1(new_n710), .C2(new_n702), .ZN(new_n1100));
  AOI211_X1 g900(.A(new_n1099), .B(new_n1100), .C1(new_n304), .C2(new_n713), .ZN(new_n1101));
  OAI221_X1 g901(.A(new_n1101), .B1(new_n489), .B2(new_n719), .C1(new_n245), .C2(new_n698), .ZN(new_n1102));
  XOR2_X1   g902(.A(new_n1102), .B(KEYINPUT58), .Z(new_n1103));
  AOI22_X1  g903(.A1(new_n713), .A2(G137), .B1(new_n699), .B2(G128), .ZN(new_n1104));
  NAND2_X1  g904(.A1(new_n925), .A2(G125), .ZN(new_n1105));
  AOI22_X1  g905(.A1(new_n730), .A2(new_n1020), .B1(new_n927), .B2(G150), .ZN(new_n1106));
  NAND3_X1  g906(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g907(.A(new_n1107), .B1(G132), .B2(new_n772), .ZN(new_n1108));
  INV_X1    g908(.A(KEYINPUT59), .ZN(new_n1109));
  AOI21_X1  g909(.A(G33), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g910(.A(G41), .B1(new_n703), .B2(G124), .ZN(new_n1111));
  OAI211_X1 g911(.A(new_n1110), .B(new_n1111), .C1(new_n775), .C2(new_n709), .ZN(new_n1112));
  NOR2_X1   g912(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1113));
  AOI21_X1  g913(.A(G41), .B1(new_n368), .B2(G33), .ZN(new_n1114));
  OAI22_X1  g914(.A1(new_n1112), .A2(new_n1113), .B1(G50), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g915(.A(new_n696), .B1(new_n1103), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g916(.A1(new_n1097), .A2(new_n742), .A3(new_n1116), .ZN(new_n1117));
  XOR2_X1   g917(.A(new_n1117), .B(KEYINPUT121), .Z(new_n1118));
  AOI21_X1  g918(.A(new_n1118), .B1(new_n919), .B2(new_n1090), .ZN(new_n1119));
  NAND2_X1  g919(.A1(new_n1096), .A2(new_n1119), .ZN(G375));
  OR2_X1    g920(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1121));
  NAND3_X1  g921(.A1(new_n1071), .A2(new_n902), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g922(.A1(new_n1038), .A2(new_n211), .ZN(new_n1123));
  NOR2_X1   g923(.A1(new_n828), .A2(new_n689), .ZN(new_n1124));
  OAI21_X1  g924(.A(new_n962), .B1(new_n710), .B2(new_n698), .ZN(new_n1125));
  XOR2_X1   g925(.A(new_n1125), .B(KEYINPUT123), .Z(new_n1126));
  NOR2_X1   g926(.A1(new_n718), .A2(new_n464), .ZN(new_n1127));
  OAI221_X1 g927(.A(new_n923), .B1(new_n207), .B2(new_n719), .C1(new_n576), .C2(new_n702), .ZN(new_n1128));
  NOR4_X1   g928(.A1(new_n1126), .A2(new_n256), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OAI221_X1 g929(.A(new_n1129), .B1(new_n489), .B2(new_n707), .C1(new_n245), .C2(new_n726), .ZN(new_n1130));
  AOI21_X1  g930(.A(new_n365), .B1(new_n772), .B2(new_n1020), .ZN(new_n1131));
  OAI21_X1  g931(.A(new_n1131), .B1(new_n222), .B2(new_n709), .ZN(new_n1132));
  OAI22_X1  g932(.A1(new_n718), .A2(new_n770), .B1(new_n707), .B2(new_n775), .ZN(new_n1133));
  AOI21_X1  g933(.A(new_n1133), .B1(G150), .B2(new_n713), .ZN(new_n1134));
  OAI21_X1  g934(.A(new_n1134), .B1(new_n217), .B2(new_n705), .ZN(new_n1135));
  AOI211_X1 g935(.A(new_n1132), .B(new_n1135), .C1(G128), .C2(new_n703), .ZN(new_n1136));
  OAI21_X1  g936(.A(new_n1136), .B1(new_n774), .B2(new_n698), .ZN(new_n1137));
  AOI21_X1  g937(.A(new_n695), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1138));
  NOR3_X1   g938(.A1(new_n1124), .A2(new_n754), .A3(new_n1138), .ZN(new_n1139));
  AOI22_X1  g939(.A1(new_n1063), .A2(new_n919), .B1(new_n1123), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g940(.A1(new_n1122), .A2(new_n1140), .ZN(G381));
  OR2_X1    g941(.A1(G390), .A2(G387), .ZN(new_n1142));
  NOR3_X1   g942(.A1(new_n1142), .A2(G396), .A3(G393), .ZN(new_n1143));
  NAND3_X1  g943(.A1(new_n1096), .A2(new_n1075), .A3(new_n1119), .ZN(new_n1144));
  NOR3_X1   g944(.A1(new_n1144), .A2(G384), .A3(G381), .ZN(new_n1145));
  NAND2_X1  g945(.A1(new_n1143), .A2(new_n1145), .ZN(G407));
  INV_X1    g946(.A(new_n1144), .ZN(new_n1147));
  NAND2_X1  g947(.A1(new_n630), .A2(G213), .ZN(new_n1148));
  INV_X1    g948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  OR2_X1    g950(.A1(new_n1150), .A2(KEYINPUT124), .ZN(new_n1151));
  NAND2_X1  g951(.A1(new_n1150), .A2(KEYINPUT124), .ZN(new_n1152));
  NAND4_X1  g952(.A1(G407), .A2(new_n1151), .A3(G213), .A4(new_n1152), .ZN(G409));
  AOI21_X1  g953(.A(new_n1149), .B1(G375), .B2(G378), .ZN(new_n1154));
  NAND4_X1  g954(.A1(new_n1079), .A2(new_n902), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1155));
  NAND3_X1  g955(.A1(new_n1119), .A2(new_n1155), .A3(new_n1075), .ZN(new_n1156));
  NAND2_X1  g956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g957(.A1(new_n1121), .A2(KEYINPUT125), .ZN(new_n1158));
  XNOR2_X1  g958(.A(new_n1158), .B(KEYINPUT60), .ZN(new_n1159));
  INV_X1    g959(.A(new_n1121), .ZN(new_n1160));
  OAI21_X1  g960(.A(new_n954), .B1(new_n1071), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g961(.A(new_n1140), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  AND2_X1   g962(.A1(new_n1162), .A2(new_n793), .ZN(new_n1163));
  NOR2_X1   g963(.A1(new_n1162), .A2(new_n793), .ZN(new_n1164));
  NOR2_X1   g964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AND2_X1   g965(.A1(new_n1149), .A2(G2897), .ZN(new_n1166));
  XNOR2_X1  g966(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  AOI21_X1  g967(.A(KEYINPUT61), .B1(new_n1157), .B2(new_n1167), .ZN(new_n1168));
  AND4_X1   g968(.A1(KEYINPUT62), .A2(new_n1154), .A3(new_n1165), .A4(new_n1156), .ZN(new_n1169));
  AOI21_X1  g969(.A(new_n1075), .B1(new_n1096), .B2(new_n1119), .ZN(new_n1170));
  INV_X1    g970(.A(new_n1156), .ZN(new_n1171));
  NOR3_X1   g971(.A1(new_n1170), .A2(new_n1149), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g972(.A(KEYINPUT62), .B1(new_n1172), .B2(new_n1165), .ZN(new_n1173));
  OAI21_X1  g973(.A(new_n1168), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g974(.A(KEYINPUT127), .ZN(new_n1175));
  NAND2_X1  g975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g976(.A(G390), .B(G387), .ZN(new_n1177));
  XNOR2_X1  g977(.A(G393), .B(G396), .ZN(new_n1178));
  INV_X1    g978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g980(.A1(G390), .A2(G387), .ZN(new_n1181));
  NAND3_X1  g981(.A1(new_n1142), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  NAND2_X1  g982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g983(.A(new_n1168), .B(KEYINPUT127), .C1(new_n1169), .C2(new_n1173), .ZN(new_n1184));
  NAND3_X1  g984(.A1(new_n1176), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g985(.A1(new_n1172), .A2(new_n1165), .ZN(new_n1186));
  INV_X1    g986(.A(new_n1186), .ZN(new_n1187));
  AOI21_X1  g987(.A(new_n1183), .B1(KEYINPUT63), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g988(.A(KEYINPUT63), .ZN(new_n1189));
  AOI21_X1  g989(.A(KEYINPUT126), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  AND3_X1   g990(.A1(new_n1186), .A2(KEYINPUT126), .A3(new_n1189), .ZN(new_n1191));
  OAI211_X1 g991(.A(new_n1188), .B(new_n1168), .C1(new_n1190), .C2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g992(.A1(new_n1185), .A2(new_n1192), .ZN(G405));
  NOR2_X1   g993(.A1(new_n1147), .A2(new_n1170), .ZN(new_n1194));
  XNOR2_X1  g994(.A(new_n1194), .B(new_n1165), .ZN(new_n1195));
  XNOR2_X1  g995(.A(new_n1195), .B(new_n1183), .ZN(G402));
endmodule


