//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1158, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT66), .ZN(G319));
  XNOR2_X1  g031(.A(KEYINPUT3), .B(G2104), .ZN(new_n457));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n457), .A2(G137), .A3(new_n458), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n458), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(KEYINPUT67), .B(G125), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n462), .B1(new_n470), .B2(G2105), .ZN(G160));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n458), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n477));
  INV_X1    g052(.A(G136), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n457), .A2(new_n458), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n475), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(G138), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n483), .B(new_n484), .C1(new_n464), .C2(new_n463), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n484), .B1(new_n457), .B2(new_n483), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n458), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n457), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT68), .B1(new_n488), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n483), .B1(new_n463), .B2(new_n464), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(new_n485), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n474), .A2(G126), .B1(new_n489), .B2(new_n491), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n511), .A2(new_n514), .ZN(G166));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT70), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(new_n509), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n518), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n519), .ZN(new_n524));
  INV_X1    g099(.A(G89), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n525), .B2(new_n507), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G168));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  INV_X1    g103(.A(G52), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n507), .A2(new_n528), .B1(new_n509), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n513), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n530), .A2(new_n532), .ZN(G171));
  AND2_X1   g108(.A1(new_n505), .A2(new_n506), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n506), .A2(G543), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT71), .B(G43), .Z(new_n536));
  AOI22_X1  g111(.A1(G81), .A2(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n513), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  NAND4_X1  g116(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND4_X1  g119(.A1(G319), .A2(G483), .A3(G661), .A4(new_n544), .ZN(G188));
  NAND2_X1  g120(.A1(G78), .A2(G543), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT72), .ZN(new_n547));
  INV_X1    g122(.A(new_n505), .ZN(new_n548));
  INV_X1    g123(.A(G65), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT73), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n547), .B(new_n552), .C1(new_n548), .C2(new_n549), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(G651), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT9), .B1(new_n509), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n506), .A2(new_n557), .A3(G53), .A4(G543), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n556), .A2(new_n558), .B1(G91), .B2(new_n534), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n554), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  INV_X1    g136(.A(G168), .ZN(G286));
  INV_X1    g137(.A(G166), .ZN(G303));
  OR2_X1    g138(.A1(new_n505), .A2(G74), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n564), .A2(G651), .B1(new_n535), .B2(G49), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n534), .A2(G87), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(G288));
  NAND3_X1  g142(.A1(new_n506), .A2(G48), .A3(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT75), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n506), .A2(new_n570), .A3(G48), .A4(G543), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n569), .A2(new_n571), .B1(new_n534), .B2(G86), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n505), .A2(G61), .ZN(new_n573));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n575), .A2(KEYINPUT74), .A3(G651), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n513), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n572), .A2(new_n576), .A3(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(G85), .A2(new_n534), .B1(new_n535), .B2(G47), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n513), .B2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n534), .A2(G92), .ZN(new_n585));
  XOR2_X1   g160(.A(new_n585), .B(KEYINPUT10), .Z(new_n586));
  NAND2_X1  g161(.A1(new_n535), .A2(KEYINPUT76), .ZN(new_n587));
  INV_X1    g162(.A(G54), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n588), .B1(new_n509), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(G79), .A2(G543), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT77), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n548), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n587), .A2(new_n590), .B1(new_n594), .B2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n586), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n584), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n584), .B1(new_n597), .B2(G868), .ZN(G321));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G299), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G168), .B2(new_n600), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(G168), .B2(new_n600), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  NOR2_X1   g180(.A1(new_n540), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n597), .A2(new_n604), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT78), .Z(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n457), .A2(new_n460), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT13), .ZN(new_n613));
  INV_X1    g188(.A(G2100), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n474), .A2(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n458), .A2(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  INV_X1    g194(.A(G135), .ZN(new_n620));
  OAI221_X1 g195(.A(new_n617), .B1(new_n618), .B2(new_n619), .C1(new_n620), .C2(new_n479), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(G156));
  INV_X1    g198(.A(KEYINPUT14), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2427), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n627), .B2(new_n626), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n629), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(G14), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n634), .A2(new_n635), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n640), .A2(new_n641), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(KEYINPUT80), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(new_n645), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n646), .A2(KEYINPUT17), .ZN(new_n649));
  OAI221_X1 g224(.A(new_n642), .B1(new_n644), .B2(new_n645), .C1(new_n648), .C2(new_n649), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n642), .A2(new_n643), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT79), .B(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2096), .B(G2100), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT81), .ZN(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT82), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT20), .Z(new_n666));
  OR2_X1    g241(.A1(new_n659), .A2(new_n661), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n664), .A3(new_n662), .ZN(new_n668));
  OAI211_X1 g243(.A(new_n666), .B(new_n668), .C1(new_n664), .C2(new_n667), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT83), .ZN(new_n670));
  XOR2_X1   g245(.A(G1981), .B(G1986), .Z(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n670), .B(new_n675), .ZN(G229));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G23), .ZN(new_n678));
  INV_X1    g253(.A(G288), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n678), .B1(new_n679), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT33), .ZN(new_n681));
  INV_X1    g256(.A(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(G6), .A2(G16), .ZN(new_n684));
  INV_X1    g259(.A(G305), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(G16), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT32), .B(G1981), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n688), .A2(KEYINPUT84), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n677), .A2(G22), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n677), .ZN(new_n691));
  INV_X1    g266(.A(G1971), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT85), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n688), .A2(KEYINPUT84), .ZN(new_n695));
  NOR4_X1   g270(.A1(new_n683), .A2(new_n689), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT34), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  MUX2_X1   g274(.A(G24), .B(G290), .S(G16), .Z(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(G1986), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n474), .A2(G119), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n458), .A2(G107), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n704));
  INV_X1    g279(.A(G131), .ZN(new_n705));
  OAI221_X1 g280(.A(new_n702), .B1(new_n703), .B2(new_n704), .C1(new_n705), .C2(new_n479), .ZN(new_n706));
  MUX2_X1   g281(.A(G25), .B(new_n706), .S(G29), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND4_X1  g284(.A1(new_n698), .A2(new_n699), .A3(new_n701), .A4(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G27), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G164), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2078), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT92), .ZN(new_n717));
  INV_X1    g292(.A(G34), .ZN(new_n718));
  AOI21_X1  g293(.A(G29), .B1(new_n718), .B2(KEYINPUT24), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(KEYINPUT24), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G160), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(new_n713), .ZN(new_n722));
  INV_X1    g297(.A(G2084), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT89), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n717), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n474), .A2(G128), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n458), .A2(G116), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n729));
  INV_X1    g304(.A(G140), .ZN(new_n730));
  OAI221_X1 g305(.A(new_n727), .B1(new_n728), .B2(new_n729), .C1(new_n730), .C2(new_n479), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT86), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n713), .A2(G26), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT87), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G2067), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n677), .A2(G20), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT23), .Z(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G299), .B2(G16), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1956), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n713), .A2(G35), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT93), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G162), .B2(new_n713), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT29), .B(G2090), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n677), .A2(G5), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G171), .B2(new_n677), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1961), .ZN(new_n751));
  INV_X1    g326(.A(G2072), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n713), .A2(G33), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT88), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT25), .ZN(new_n756));
  INV_X1    g331(.A(G139), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n457), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  OAI221_X1 g333(.A(new_n756), .B1(new_n757), .B2(new_n479), .C1(new_n458), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n753), .B1(new_n759), .B2(G29), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n751), .B1(new_n752), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n739), .A2(new_n743), .A3(new_n748), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n540), .A2(G16), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G16), .B2(G19), .ZN(new_n764));
  INV_X1    g339(.A(G1341), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n760), .A2(new_n752), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n713), .A2(G32), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT90), .B(KEYINPUT26), .Z(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n460), .A2(G105), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(G129), .ZN(new_n774));
  INV_X1    g349(.A(G141), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n774), .A2(new_n493), .B1(new_n479), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n768), .B1(new_n777), .B2(new_n713), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT27), .B(G1996), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT31), .B(G11), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT91), .B(G28), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(KEYINPUT30), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(KEYINPUT30), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n783), .A2(new_n713), .A3(new_n784), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n781), .B(new_n785), .C1(new_n621), .C2(new_n713), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n764), .B2(new_n765), .ZN(new_n787));
  AND4_X1   g362(.A1(new_n766), .A2(new_n767), .A3(new_n780), .A4(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G168), .A2(new_n677), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n677), .B2(G21), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n677), .A2(G4), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n597), .B2(new_n677), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n791), .A2(G1966), .B1(new_n793), .B2(G1348), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(G1348), .ZN(new_n795));
  INV_X1    g370(.A(G1966), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n790), .A2(new_n796), .B1(new_n723), .B2(new_n722), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n788), .A2(new_n794), .A3(new_n795), .A4(new_n797), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n712), .A2(new_n726), .A3(new_n762), .A4(new_n798), .ZN(G311));
  OR4_X1    g374(.A1(new_n712), .A2(new_n726), .A3(new_n762), .A4(new_n798), .ZN(G150));
  INV_X1    g375(.A(KEYINPUT94), .ZN(new_n801));
  INV_X1    g376(.A(G93), .ZN(new_n802));
  INV_X1    g377(.A(G55), .ZN(new_n803));
  OAI22_X1  g378(.A1(new_n507), .A2(new_n802), .B1(new_n509), .B2(new_n803), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n805), .A2(new_n513), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n540), .B1(new_n801), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n801), .B2(new_n808), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n540), .A2(KEYINPUT94), .A3(new_n807), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT38), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n597), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n816));
  INV_X1    g391(.A(G860), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n807), .A2(new_n817), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT37), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(G145));
  NAND2_X1  g397(.A1(new_n499), .A2(new_n501), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n731), .B(new_n823), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n759), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n777), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n706), .B(KEYINPUT96), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n612), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n474), .A2(G130), .ZN(new_n829));
  NOR3_X1   g404(.A1(new_n458), .A2(KEYINPUT95), .A3(G118), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT95), .B1(new_n458), .B2(G118), .ZN(new_n831));
  OR2_X1    g406(.A1(G106), .A2(G2105), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n831), .A2(G2104), .A3(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G142), .ZN(new_n834));
  OAI221_X1 g409(.A(new_n829), .B1(new_n830), .B2(new_n833), .C1(new_n834), .C2(new_n479), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n828), .B(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n826), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n826), .A2(new_n836), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(G160), .B(new_n621), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G162), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n836), .A2(new_n826), .A3(KEYINPUT97), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n842), .B1(new_n836), .B2(new_n826), .ZN(new_n845));
  AOI21_X1  g420(.A(G37), .B1(new_n837), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g423(.A(KEYINPUT101), .B1(new_n807), .B2(G868), .ZN(new_n849));
  XNOR2_X1  g424(.A(G166), .B(KEYINPUT100), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n685), .ZN(new_n851));
  XNOR2_X1  g426(.A(G290), .B(G288), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT42), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n810), .A2(new_n811), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n607), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n596), .B(G299), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT41), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n596), .A2(new_n554), .A3(new_n559), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n860), .B(new_n861), .C1(new_n859), .C2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(KEYINPUT99), .B(KEYINPUT41), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n858), .B1(new_n866), .B2(new_n856), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n600), .B1(new_n854), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n868), .B1(new_n854), .B2(new_n867), .ZN(new_n869));
  MUX2_X1   g444(.A(KEYINPUT101), .B(new_n849), .S(new_n869), .Z(G295));
  MUX2_X1   g445(.A(KEYINPUT101), .B(new_n849), .S(new_n869), .Z(G331));
  NAND3_X1  g446(.A1(G168), .A2(KEYINPUT102), .A3(G171), .ZN(new_n872));
  NAND2_X1  g447(.A1(G171), .A2(KEYINPUT102), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n874));
  NAND2_X1  g449(.A1(G301), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(G286), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n812), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n872), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n855), .ZN(new_n879));
  AOI22_X1  g454(.A1(new_n863), .A2(new_n865), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n879), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n881), .A2(new_n857), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n853), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n886));
  INV_X1    g461(.A(G37), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n853), .B1(new_n880), .B2(new_n882), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT103), .ZN(new_n890));
  AOI21_X1  g465(.A(G37), .B1(new_n883), .B2(new_n884), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n891), .A2(new_n892), .A3(new_n886), .A4(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n860), .B1(new_n859), .B2(new_n862), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n881), .A2(KEYINPUT41), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n857), .B1(new_n881), .B2(new_n864), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n853), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n891), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n895), .B1(new_n900), .B2(KEYINPUT43), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n894), .A2(KEYINPUT104), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT104), .B1(new_n894), .B2(new_n901), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n900), .A2(KEYINPUT43), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n886), .B1(new_n891), .B2(new_n888), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI22_X1  g481(.A1(new_n902), .A2(new_n903), .B1(new_n906), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g482(.A(KEYINPUT123), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT53), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n470), .A2(G2105), .ZN(new_n910));
  INV_X1    g485(.A(new_n462), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(G40), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(G1384), .B1(new_n499), .B2(new_n501), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT45), .ZN(new_n915));
  AOI21_X1  g490(.A(G1384), .B1(new_n496), .B2(new_n502), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n913), .B(new_n915), .C1(new_n916), .C2(KEYINPUT45), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n909), .B1(new_n917), .B2(G2078), .ZN(new_n918));
  XNOR2_X1  g493(.A(KEYINPUT121), .B(G1961), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT50), .ZN(new_n920));
  INV_X1    g495(.A(G1384), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n503), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n914), .A2(new_n920), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n923), .A2(G40), .A3(G160), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n919), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT122), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT45), .B1(new_n823), .B2(new_n921), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n927), .A2(new_n912), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n500), .B1(new_n499), .B2(new_n501), .ZN(new_n930));
  OAI211_X1 g505(.A(KEYINPUT45), .B(new_n921), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n909), .A2(G2078), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n925), .A2(new_n926), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n926), .B1(new_n925), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n918), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(G171), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n913), .B(new_n923), .C1(new_n916), .C2(new_n920), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n915), .A2(new_n932), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n938), .A2(new_n919), .B1(new_n928), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n918), .A3(G301), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT54), .B1(new_n937), .B2(new_n941), .ZN(new_n942));
  OAI211_X1 g517(.A(G301), .B(new_n918), .C1(new_n934), .C2(new_n935), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT54), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n918), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(G171), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT55), .ZN(new_n948));
  INV_X1    g523(.A(G8), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n948), .B1(G166), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g525(.A(KEYINPUT55), .B(G8), .C1(new_n511), .C2(new_n514), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g527(.A(G160), .B(G40), .C1(new_n914), .C2(new_n920), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(new_n916), .B2(new_n920), .ZN(new_n954));
  INV_X1    g529(.A(G2090), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n692), .A2(new_n917), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n952), .B1(new_n956), .B2(new_n949), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT49), .ZN(new_n958));
  INV_X1    g533(.A(G1981), .ZN(new_n959));
  AND2_X1   g534(.A1(new_n576), .A2(new_n579), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n960), .B2(new_n572), .ZN(new_n961));
  AND4_X1   g536(.A1(new_n959), .A2(new_n572), .A3(new_n576), .A4(new_n579), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(G160), .A2(new_n914), .A3(G40), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(new_n949), .ZN(new_n966));
  NAND2_X1  g541(.A1(G305), .A2(G1981), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n960), .A2(new_n959), .A3(new_n572), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n968), .A3(KEYINPUT49), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n963), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n565), .A2(G1976), .A3(new_n566), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n964), .A2(G8), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n964), .A2(KEYINPUT107), .A3(G8), .A4(new_n971), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(KEYINPUT52), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT52), .B1(G288), .B2(new_n682), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n966), .A2(new_n971), .A3(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n970), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n950), .A2(KEYINPUT106), .A3(new_n951), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT106), .B1(new_n950), .B2(new_n951), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n915), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n921), .B1(new_n929), .B2(new_n930), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n983), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(G1971), .B1(new_n986), .B2(new_n913), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n938), .A2(G2090), .ZN(new_n988));
  OAI211_X1 g563(.A(G8), .B(new_n982), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n957), .A2(new_n979), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n947), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n942), .A2(new_n991), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n922), .A2(G2084), .A3(new_n924), .ZN(new_n993));
  AOI21_X1  g568(.A(G1966), .B1(new_n928), .B2(new_n931), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT119), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n928), .A2(new_n931), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n796), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n912), .B1(new_n920), .B2(new_n914), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n999), .A3(new_n723), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT119), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(G286), .B1(new_n995), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(new_n949), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT120), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n997), .A2(new_n1001), .A3(new_n1000), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1001), .B1(new_n997), .B2(new_n1000), .ZN(new_n1009));
  OAI21_X1  g584(.A(G168), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT120), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1011), .A3(new_n1005), .ZN(new_n1012));
  OAI21_X1  g587(.A(G8), .B1(new_n993), .B2(new_n994), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1013), .B(new_n1004), .C1(new_n949), .C2(G168), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1007), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n995), .A2(G8), .A3(G286), .A4(new_n1002), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n992), .A2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n920), .B(new_n921), .C1(new_n929), .C2(new_n930), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n823), .A2(new_n921), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT50), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n913), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1956), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n985), .A2(new_n984), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT56), .B(G2072), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(new_n913), .A3(new_n915), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n1029));
  AOI211_X1 g604(.A(KEYINPUT111), .B(new_n1029), .C1(new_n554), .C2(new_n559), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(KEYINPUT111), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1029), .A2(KEYINPUT111), .ZN(new_n1032));
  AND4_X1   g607(.A1(new_n554), .A2(new_n559), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1028), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT61), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1024), .A2(new_n1027), .A3(new_n1034), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1036), .A2(KEYINPUT117), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1042), .A2(new_n1037), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1040), .A2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n912), .A2(G1996), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1045), .B(new_n915), .C1(new_n916), .C2(KEYINPUT45), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1025), .A2(KEYINPUT112), .A3(new_n915), .A4(new_n1045), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(G1341), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n964), .A2(KEYINPUT114), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT114), .B1(new_n964), .B2(new_n1051), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1048), .A2(new_n1049), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(new_n540), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1058), .A2(KEYINPUT115), .A3(KEYINPUT116), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1055), .A2(new_n540), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1055), .A2(new_n540), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT115), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1059), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT118), .B1(new_n1044), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1042), .A2(new_n1037), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1039), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1055), .A2(new_n540), .A3(new_n1060), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n1055), .B2(new_n540), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1069), .A2(new_n1070), .A3(new_n1059), .A4(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G1348), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n938), .A2(new_n1076), .B1(new_n738), .B2(new_n965), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1077), .A2(KEYINPUT60), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(KEYINPUT60), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n597), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(KEYINPUT60), .A3(new_n596), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1065), .A2(new_n1075), .A3(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1036), .B1(new_n1077), .B2(new_n596), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1085), .A2(new_n1038), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1018), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1013), .A2(G286), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n990), .A2(KEYINPUT110), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT63), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1089), .A2(new_n957), .A3(new_n989), .A4(new_n979), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT110), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n987), .A2(new_n988), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n952), .B1(new_n1096), .B2(new_n949), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1013), .A2(new_n1091), .A3(G286), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1097), .A2(new_n1098), .A3(new_n989), .A4(new_n979), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n989), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n979), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n679), .A2(new_n682), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(KEYINPUT108), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n970), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n968), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT109), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n949), .B(new_n965), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1107), .B2(new_n1106), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1100), .A2(new_n1102), .A3(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n908), .B1(new_n1088), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1102), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1074), .B(new_n1059), .C1(new_n1043), .C2(new_n1040), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1082), .B1(new_n1114), .B2(KEYINPUT118), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1086), .B1(new_n1115), .B2(new_n1075), .ZN(new_n1116));
  OAI211_X1 g691(.A(KEYINPUT123), .B(new_n1113), .C1(new_n1116), .C2(new_n1018), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n990), .A2(G171), .A3(new_n936), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1111), .A2(new_n1117), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n913), .A2(new_n927), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n731), .B(G2067), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(new_n1126), .B(KEYINPUT105), .Z(new_n1127));
  XNOR2_X1  g702(.A(new_n777), .B(G1996), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n708), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n706), .B(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1129), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(G290), .A2(G1986), .ZN(new_n1133));
  AND2_X1   g708(.A1(G290), .A2(G1986), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1124), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1122), .A2(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n1123), .A2(G1996), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT46), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT124), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1125), .A2(new_n773), .A3(new_n776), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1141), .B(new_n1142), .C1(new_n1123), .C2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT47), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1124), .A2(new_n1133), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1149));
  XNOR2_X1  g724(.A(new_n1148), .B(new_n1149), .ZN(new_n1150));
  OR2_X1    g725(.A1(new_n706), .A2(new_n1130), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1129), .A2(new_n1151), .B1(G2067), .B2(new_n731), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1132), .A2(new_n1150), .B1(new_n1152), .B2(new_n1124), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1147), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1137), .A2(new_n1155), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g731(.A1(new_n656), .A2(new_n455), .ZN(new_n1158));
  NOR3_X1   g732(.A1(G229), .A2(G401), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g733(.A1(new_n847), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g734(.A1(new_n906), .A2(new_n1160), .ZN(G308));
  INV_X1    g735(.A(G308), .ZN(G225));
endmodule


