

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n568), .A2(n527), .ZN(n804) );
  XNOR2_X1 U553 ( .A(n596), .B(KEYINPUT27), .ZN(n597) );
  INV_X1 U554 ( .A(n649), .ZN(n676) );
  AND2_X1 U555 ( .A1(n683), .A2(n682), .ZN(n684) );
  AND2_X1 U556 ( .A1(n592), .A2(n591), .ZN(n774) );
  AND2_X2 U557 ( .A1(n541), .A2(G2105), .ZN(n893) );
  BUF_X1 U558 ( .A(n543), .Z(n541) );
  NAND2_X2 U559 ( .A1(G8), .A2(n676), .ZN(n675) );
  XNOR2_X1 U560 ( .A(n634), .B(n633), .ZN(n636) );
  AND2_X1 U561 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U562 ( .A1(n647), .A2(n932), .ZN(n595) );
  INV_X1 U563 ( .A(KEYINPUT28), .ZN(n605) );
  NOR2_X1 U564 ( .A1(n641), .A2(n640), .ZN(n642) );
  INV_X1 U565 ( .A(G2105), .ZN(n536) );
  INV_X1 U566 ( .A(G2104), .ZN(n535) );
  INV_X1 U567 ( .A(KEYINPUT23), .ZN(n544) );
  XOR2_X1 U568 ( .A(n656), .B(n655), .Z(n518) );
  OR2_X1 U569 ( .A1(n675), .A2(n716), .ZN(n519) );
  AND2_X1 U570 ( .A1(n676), .A2(G1341), .ZN(n520) );
  AND2_X1 U571 ( .A1(n767), .A2(n1013), .ZN(n521) );
  AND2_X1 U572 ( .A1(n649), .A2(G1996), .ZN(n609) );
  INV_X1 U573 ( .A(KEYINPUT94), .ZN(n633) );
  NOR2_X1 U574 ( .A1(n636), .A2(n635), .ZN(n639) );
  INV_X1 U575 ( .A(n647), .ZN(n648) );
  NOR2_X1 U576 ( .A1(G168), .A2(n518), .ZN(n659) );
  INV_X1 U577 ( .A(n736), .ZN(n594) );
  AND2_X2 U578 ( .A1(n735), .A2(n594), .ZN(n649) );
  NOR2_X1 U579 ( .A1(n774), .A2(G1384), .ZN(n593) );
  XNOR2_X1 U580 ( .A(G2104), .B(KEYINPUT66), .ZN(n540) );
  INV_X1 U581 ( .A(KEYINPUT100), .ZN(n713) );
  NAND2_X1 U582 ( .A1(G160), .A2(G40), .ZN(n736) );
  NOR2_X1 U583 ( .A1(G651), .A2(n568), .ZN(n799) );
  XNOR2_X1 U584 ( .A(n545), .B(n544), .ZN(n546) );
  BUF_X1 U585 ( .A(n774), .Z(G164) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n568) );
  NAND2_X1 U587 ( .A1(G51), .A2(n799), .ZN(n524) );
  INV_X1 U588 ( .A(G651), .ZN(n527) );
  NOR2_X1 U589 ( .A1(G543), .A2(n527), .ZN(n522) );
  XOR2_X2 U590 ( .A(KEYINPUT1), .B(n522), .Z(n800) );
  NAND2_X1 U591 ( .A1(G63), .A2(n800), .ZN(n523) );
  NAND2_X1 U592 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U593 ( .A(KEYINPUT6), .B(n525), .ZN(n532) );
  NOR2_X1 U594 ( .A1(G543), .A2(G651), .ZN(n803) );
  NAND2_X1 U595 ( .A1(n803), .A2(G89), .ZN(n526) );
  XNOR2_X1 U596 ( .A(n526), .B(KEYINPUT4), .ZN(n529) );
  NAND2_X1 U597 ( .A1(G76), .A2(n804), .ZN(n528) );
  NAND2_X1 U598 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U599 ( .A(n530), .B(KEYINPUT5), .Z(n531) );
  NOR2_X1 U600 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U601 ( .A(KEYINPUT7), .B(n533), .Z(n534) );
  XOR2_X1 U602 ( .A(KEYINPUT75), .B(n534), .Z(G168) );
  AND2_X1 U603 ( .A1(G2105), .A2(G2104), .ZN(n892) );
  NAND2_X1 U604 ( .A1(n892), .A2(G113), .ZN(n539) );
  NAND2_X1 U605 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X2 U606 ( .A(n537), .B(KEYINPUT17), .ZN(n888) );
  NAND2_X1 U607 ( .A1(n888), .A2(G137), .ZN(n538) );
  NAND2_X1 U608 ( .A1(n539), .A2(n538), .ZN(n549) );
  INV_X1 U609 ( .A(n540), .ZN(n543) );
  NAND2_X1 U610 ( .A1(G125), .A2(n893), .ZN(n542) );
  XOR2_X1 U611 ( .A(KEYINPUT67), .B(n542), .Z(n547) );
  NOR2_X2 U612 ( .A1(n543), .A2(G2105), .ZN(n584) );
  BUF_X2 U613 ( .A(n584), .Z(n889) );
  NAND2_X1 U614 ( .A1(G101), .A2(n889), .ZN(n545) );
  NAND2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X2 U616 ( .A1(n549), .A2(n548), .ZN(G160) );
  NAND2_X1 U617 ( .A1(G52), .A2(n799), .ZN(n551) );
  NAND2_X1 U618 ( .A1(G64), .A2(n800), .ZN(n550) );
  NAND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n803), .A2(G90), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n552), .B(KEYINPUT68), .ZN(n554) );
  NAND2_X1 U622 ( .A1(G77), .A2(n804), .ZN(n553) );
  NAND2_X1 U623 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U624 ( .A(KEYINPUT9), .B(n555), .Z(n556) );
  NOR2_X1 U625 ( .A1(n557), .A2(n556), .ZN(G171) );
  INV_X1 U626 ( .A(G171), .ZN(G301) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G88), .A2(n803), .ZN(n559) );
  NAND2_X1 U629 ( .A1(G75), .A2(n804), .ZN(n558) );
  NAND2_X1 U630 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U631 ( .A1(G50), .A2(n799), .ZN(n561) );
  NAND2_X1 U632 ( .A1(G62), .A2(n800), .ZN(n560) );
  NAND2_X1 U633 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U634 ( .A1(n563), .A2(n562), .ZN(G166) );
  INV_X1 U635 ( .A(G166), .ZN(G303) );
  NAND2_X1 U636 ( .A1(G49), .A2(n799), .ZN(n565) );
  NAND2_X1 U637 ( .A1(G74), .A2(G651), .ZN(n564) );
  NAND2_X1 U638 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U639 ( .A(KEYINPUT78), .B(n566), .ZN(n567) );
  NOR2_X1 U640 ( .A1(n800), .A2(n567), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n568), .A2(G87), .ZN(n569) );
  NAND2_X1 U642 ( .A1(n570), .A2(n569), .ZN(G288) );
  NAND2_X1 U643 ( .A1(G86), .A2(n803), .ZN(n572) );
  NAND2_X1 U644 ( .A1(G48), .A2(n799), .ZN(n571) );
  NAND2_X1 U645 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U646 ( .A1(n804), .A2(G73), .ZN(n573) );
  XOR2_X1 U647 ( .A(KEYINPUT2), .B(n573), .Z(n574) );
  NOR2_X1 U648 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n800), .A2(G61), .ZN(n576) );
  NAND2_X1 U650 ( .A1(n577), .A2(n576), .ZN(G305) );
  NAND2_X1 U651 ( .A1(G85), .A2(n803), .ZN(n579) );
  NAND2_X1 U652 ( .A1(G72), .A2(n804), .ZN(n578) );
  NAND2_X1 U653 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U654 ( .A1(G47), .A2(n799), .ZN(n581) );
  NAND2_X1 U655 ( .A1(G60), .A2(n800), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n581), .A2(n580), .ZN(n582) );
  OR2_X1 U657 ( .A1(n583), .A2(n582), .ZN(G290) );
  NAND2_X1 U658 ( .A1(n584), .A2(G102), .ZN(n585) );
  XNOR2_X1 U659 ( .A(n585), .B(KEYINPUT82), .ZN(n587) );
  NAND2_X1 U660 ( .A1(G138), .A2(n888), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U662 ( .A(n588), .B(KEYINPUT83), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G114), .A2(n892), .ZN(n590) );
  NAND2_X1 U664 ( .A1(G126), .A2(n893), .ZN(n589) );
  AND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U666 ( .A(n593), .B(KEYINPUT64), .ZN(n735) );
  XNOR2_X2 U667 ( .A(n649), .B(KEYINPUT90), .ZN(n647) );
  XNOR2_X1 U668 ( .A(G1956), .B(KEYINPUT91), .ZN(n932) );
  XNOR2_X1 U669 ( .A(n595), .B(KEYINPUT92), .ZN(n598) );
  NAND2_X1 U670 ( .A1(G2072), .A2(n647), .ZN(n596) );
  NOR2_X2 U671 ( .A1(n598), .A2(n597), .ZN(n607) );
  NAND2_X1 U672 ( .A1(G53), .A2(n799), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G65), .A2(n800), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U675 ( .A1(G91), .A2(n803), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G78), .A2(n804), .ZN(n601) );
  NAND2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n1009) );
  NOR2_X1 U679 ( .A1(n607), .A2(n1009), .ZN(n606) );
  XNOR2_X1 U680 ( .A(n606), .B(n605), .ZN(n645) );
  NAND2_X1 U681 ( .A1(n607), .A2(n1009), .ZN(n643) );
  XNOR2_X1 U682 ( .A(KEYINPUT26), .B(KEYINPUT93), .ZN(n608) );
  XNOR2_X1 U683 ( .A(n609), .B(n608), .ZN(n621) );
  NAND2_X1 U684 ( .A1(G68), .A2(n804), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n803), .A2(G81), .ZN(n610) );
  XNOR2_X1 U686 ( .A(n610), .B(KEYINPUT12), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U688 ( .A(n613), .B(KEYINPUT13), .ZN(n615) );
  NAND2_X1 U689 ( .A1(G43), .A2(n799), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n800), .A2(G56), .ZN(n616) );
  XOR2_X1 U692 ( .A(KEYINPUT14), .B(n616), .Z(n617) );
  NOR2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U694 ( .A(KEYINPUT71), .B(n619), .ZN(n1025) );
  NOR2_X1 U695 ( .A1(n520), .A2(n1025), .ZN(n620) );
  XNOR2_X1 U696 ( .A(n622), .B(KEYINPUT65), .ZN(n638) );
  NAND2_X1 U697 ( .A1(G66), .A2(n800), .ZN(n629) );
  NAND2_X1 U698 ( .A1(G79), .A2(n804), .ZN(n624) );
  NAND2_X1 U699 ( .A1(G54), .A2(n799), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n803), .A2(G92), .ZN(n625) );
  XOR2_X1 U702 ( .A(KEYINPUT72), .B(n625), .Z(n626) );
  NOR2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n630), .B(KEYINPUT15), .ZN(n632) );
  XOR2_X1 U706 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n631) );
  XNOR2_X1 U707 ( .A(n632), .B(n631), .ZN(n1014) );
  NAND2_X1 U708 ( .A1(n676), .A2(G1348), .ZN(n634) );
  AND2_X1 U709 ( .A1(n647), .A2(G2067), .ZN(n635) );
  NOR2_X1 U710 ( .A1(n1014), .A2(n639), .ZN(n637) );
  NOR2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n641) );
  AND2_X1 U712 ( .A1(n1014), .A2(n639), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U715 ( .A(n646), .B(KEYINPUT29), .ZN(n653) );
  XOR2_X1 U716 ( .A(KEYINPUT25), .B(G2078), .Z(n964) );
  NOR2_X1 U717 ( .A1(n964), .A2(n648), .ZN(n651) );
  NOR2_X1 U718 ( .A1(n649), .A2(G1961), .ZN(n650) );
  NOR2_X1 U719 ( .A1(n651), .A2(n650), .ZN(n657) );
  NOR2_X1 U720 ( .A1(G301), .A2(n657), .ZN(n652) );
  NOR2_X1 U721 ( .A1(n653), .A2(n652), .ZN(n662) );
  XNOR2_X1 U722 ( .A(KEYINPUT95), .B(KEYINPUT30), .ZN(n656) );
  NOR2_X1 U723 ( .A1(G2084), .A2(n676), .ZN(n666) );
  NOR2_X1 U724 ( .A1(G1966), .A2(n675), .ZN(n663) );
  NOR2_X1 U725 ( .A1(n666), .A2(n663), .ZN(n654) );
  NAND2_X1 U726 ( .A1(n654), .A2(G8), .ZN(n655) );
  AND2_X1 U727 ( .A1(G301), .A2(n657), .ZN(n658) );
  NOR2_X1 U728 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n660), .B(KEYINPUT31), .ZN(n661) );
  NOR2_X2 U730 ( .A1(n662), .A2(n661), .ZN(n672) );
  XNOR2_X1 U731 ( .A(n672), .B(KEYINPUT96), .ZN(n664) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U733 ( .A(KEYINPUT97), .B(n665), .ZN(n668) );
  AND2_X1 U734 ( .A1(G8), .A2(n666), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n670) );
  INV_X1 U736 ( .A(KEYINPUT98), .ZN(n669) );
  XNOR2_X1 U737 ( .A(n670), .B(n669), .ZN(n697) );
  INV_X1 U738 ( .A(KEYINPUT96), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n672), .B(n671), .ZN(n674) );
  AND2_X1 U740 ( .A1(G286), .A2(G8), .ZN(n673) );
  NAND2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n683) );
  INV_X1 U742 ( .A(G8), .ZN(n681) );
  NOR2_X1 U743 ( .A1(G1971), .A2(n675), .ZN(n678) );
  NOR2_X1 U744 ( .A1(G2090), .A2(n676), .ZN(n677) );
  NOR2_X1 U745 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U746 ( .A1(n679), .A2(G303), .ZN(n680) );
  OR2_X1 U747 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U748 ( .A(n684), .B(KEYINPUT32), .ZN(n691) );
  AND2_X1 U749 ( .A1(n691), .A2(n675), .ZN(n685) );
  NAND2_X1 U750 ( .A1(n697), .A2(n685), .ZN(n690) );
  INV_X1 U751 ( .A(n675), .ZN(n688) );
  NOR2_X1 U752 ( .A1(G2090), .A2(G303), .ZN(n686) );
  NAND2_X1 U753 ( .A1(G8), .A2(n686), .ZN(n687) );
  OR2_X1 U754 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U755 ( .A1(n690), .A2(n689), .ZN(n712) );
  NAND2_X1 U756 ( .A1(G1976), .A2(G288), .ZN(n1023) );
  AND2_X1 U757 ( .A1(n691), .A2(n1023), .ZN(n696) );
  NOR2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n692) );
  XOR2_X1 U759 ( .A(KEYINPUT99), .B(n692), .Z(n702) );
  INV_X1 U760 ( .A(n702), .ZN(n1010) );
  NOR2_X1 U761 ( .A1(n675), .A2(n1010), .ZN(n693) );
  AND2_X1 U762 ( .A1(KEYINPUT33), .A2(n693), .ZN(n694) );
  XNOR2_X1 U763 ( .A(G1981), .B(G305), .ZN(n1019) );
  OR2_X1 U764 ( .A1(n694), .A2(n1019), .ZN(n699) );
  OR2_X1 U765 ( .A1(n675), .A2(n699), .ZN(n706) );
  INV_X1 U766 ( .A(n706), .ZN(n695) );
  AND2_X1 U767 ( .A1(n696), .A2(n695), .ZN(n698) );
  NAND2_X1 U768 ( .A1(n698), .A2(n697), .ZN(n710) );
  INV_X1 U769 ( .A(n699), .ZN(n700) );
  NAND2_X1 U770 ( .A1(n700), .A2(KEYINPUT33), .ZN(n708) );
  INV_X1 U771 ( .A(n1023), .ZN(n704) );
  NOR2_X1 U772 ( .A1(G1971), .A2(G303), .ZN(n701) );
  NOR2_X1 U773 ( .A1(n702), .A2(n701), .ZN(n703) );
  OR2_X1 U774 ( .A1(n704), .A2(n703), .ZN(n705) );
  OR2_X1 U775 ( .A1(n706), .A2(n705), .ZN(n707) );
  AND2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n714) );
  XNOR2_X1 U779 ( .A(n714), .B(n713), .ZN(n717) );
  NOR2_X1 U780 ( .A1(G1981), .A2(G305), .ZN(n715) );
  XOR2_X1 U781 ( .A(n715), .B(KEYINPUT24), .Z(n716) );
  NAND2_X1 U782 ( .A1(n717), .A2(n519), .ZN(n740) );
  NAND2_X1 U783 ( .A1(G107), .A2(n892), .ZN(n719) );
  NAND2_X1 U784 ( .A1(G131), .A2(n888), .ZN(n718) );
  NAND2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U786 ( .A1(G119), .A2(n893), .ZN(n721) );
  NAND2_X1 U787 ( .A1(G95), .A2(n889), .ZN(n720) );
  NAND2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n722) );
  OR2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n905) );
  NAND2_X1 U790 ( .A1(G1991), .A2(n905), .ZN(n734) );
  XOR2_X1 U791 ( .A(KEYINPUT87), .B(KEYINPUT38), .Z(n725) );
  NAND2_X1 U792 ( .A1(G105), .A2(n889), .ZN(n724) );
  XNOR2_X1 U793 ( .A(n725), .B(n724), .ZN(n732) );
  NAND2_X1 U794 ( .A1(G117), .A2(n892), .ZN(n727) );
  NAND2_X1 U795 ( .A1(G141), .A2(n888), .ZN(n726) );
  NAND2_X1 U796 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U797 ( .A1(n893), .A2(G129), .ZN(n728) );
  XOR2_X1 U798 ( .A(KEYINPUT86), .B(n728), .Z(n729) );
  NOR2_X1 U799 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U800 ( .A1(n732), .A2(n731), .ZN(n886) );
  NAND2_X1 U801 ( .A1(G1996), .A2(n886), .ZN(n733) );
  NAND2_X1 U802 ( .A1(n734), .A2(n733), .ZN(n983) );
  NOR2_X1 U803 ( .A1(n736), .A2(n735), .ZN(n767) );
  NAND2_X1 U804 ( .A1(n983), .A2(n767), .ZN(n737) );
  XOR2_X1 U805 ( .A(KEYINPUT88), .B(n737), .Z(n758) );
  XOR2_X1 U806 ( .A(n758), .B(KEYINPUT89), .Z(n738) );
  XNOR2_X1 U807 ( .A(G1986), .B(G290), .ZN(n1013) );
  NOR2_X1 U808 ( .A1(n738), .A2(n521), .ZN(n739) );
  NAND2_X1 U809 ( .A1(n740), .A2(n739), .ZN(n753) );
  NAND2_X1 U810 ( .A1(G104), .A2(n889), .ZN(n742) );
  NAND2_X1 U811 ( .A1(n888), .A2(G140), .ZN(n741) );
  NAND2_X1 U812 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U813 ( .A(n743), .B(KEYINPUT34), .ZN(n744) );
  XNOR2_X1 U814 ( .A(KEYINPUT84), .B(n744), .ZN(n749) );
  NAND2_X1 U815 ( .A1(G116), .A2(n892), .ZN(n746) );
  NAND2_X1 U816 ( .A1(G128), .A2(n893), .ZN(n745) );
  NAND2_X1 U817 ( .A1(n746), .A2(n745), .ZN(n747) );
  XOR2_X1 U818 ( .A(KEYINPUT35), .B(n747), .Z(n748) );
  NOR2_X1 U819 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U820 ( .A(KEYINPUT36), .B(n750), .ZN(n904) );
  XNOR2_X1 U821 ( .A(G2067), .B(KEYINPUT37), .ZN(n765) );
  NOR2_X1 U822 ( .A1(n904), .A2(n765), .ZN(n984) );
  NAND2_X1 U823 ( .A1(n984), .A2(n767), .ZN(n751) );
  XOR2_X1 U824 ( .A(KEYINPUT85), .B(n751), .Z(n764) );
  INV_X1 U825 ( .A(n764), .ZN(n752) );
  NOR2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n771) );
  NOR2_X1 U827 ( .A1(G1996), .A2(n886), .ZN(n754) );
  XOR2_X1 U828 ( .A(KEYINPUT101), .B(n754), .Z(n980) );
  NOR2_X1 U829 ( .A1(G1986), .A2(G290), .ZN(n756) );
  NOR2_X1 U830 ( .A1(G1991), .A2(n905), .ZN(n755) );
  XNOR2_X1 U831 ( .A(KEYINPUT102), .B(n755), .ZN(n990) );
  NOR2_X1 U832 ( .A1(n756), .A2(n990), .ZN(n757) );
  NOR2_X1 U833 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U834 ( .A(KEYINPUT103), .B(n759), .Z(n760) );
  NOR2_X1 U835 ( .A1(n980), .A2(n760), .ZN(n761) );
  XNOR2_X1 U836 ( .A(n761), .B(KEYINPUT104), .ZN(n762) );
  XNOR2_X1 U837 ( .A(n762), .B(KEYINPUT39), .ZN(n763) );
  NAND2_X1 U838 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U839 ( .A1(n904), .A2(n765), .ZN(n985) );
  NAND2_X1 U840 ( .A1(n766), .A2(n985), .ZN(n768) );
  NAND2_X1 U841 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U842 ( .A(n769), .B(KEYINPUT105), .ZN(n770) );
  NOR2_X2 U843 ( .A1(n771), .A2(n770), .ZN(n773) );
  INV_X1 U844 ( .A(KEYINPUT40), .ZN(n772) );
  XNOR2_X1 U845 ( .A(n773), .B(n772), .ZN(G329) );
  AND2_X1 U846 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U847 ( .A1(G111), .A2(n892), .ZN(n776) );
  NAND2_X1 U848 ( .A1(G135), .A2(n888), .ZN(n775) );
  NAND2_X1 U849 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U850 ( .A1(n893), .A2(G123), .ZN(n777) );
  XOR2_X1 U851 ( .A(KEYINPUT18), .B(n777), .Z(n778) );
  NOR2_X1 U852 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U853 ( .A1(n889), .A2(G99), .ZN(n780) );
  NAND2_X1 U854 ( .A1(n781), .A2(n780), .ZN(n987) );
  XNOR2_X1 U855 ( .A(G2096), .B(n987), .ZN(n782) );
  OR2_X1 U856 ( .A1(G2100), .A2(n782), .ZN(G156) );
  INV_X1 U857 ( .A(G57), .ZN(G237) );
  INV_X1 U858 ( .A(G132), .ZN(G219) );
  NAND2_X1 U859 ( .A1(G7), .A2(G661), .ZN(n783) );
  XNOR2_X1 U860 ( .A(n783), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U861 ( .A(G223), .B(KEYINPUT70), .Z(n835) );
  NAND2_X1 U862 ( .A1(n835), .A2(G567), .ZN(n784) );
  XOR2_X1 U863 ( .A(KEYINPUT11), .B(n784), .Z(G234) );
  INV_X1 U864 ( .A(G860), .ZN(n798) );
  OR2_X1 U865 ( .A1(n1025), .A2(n798), .ZN(G153) );
  INV_X1 U866 ( .A(n1014), .ZN(n863) );
  NOR2_X1 U867 ( .A1(n863), .A2(G868), .ZN(n786) );
  INV_X1 U868 ( .A(G868), .ZN(n787) );
  NOR2_X1 U869 ( .A1(n787), .A2(G301), .ZN(n785) );
  NOR2_X1 U870 ( .A1(n786), .A2(n785), .ZN(G284) );
  INV_X1 U871 ( .A(n1009), .ZN(G299) );
  NOR2_X1 U872 ( .A1(G286), .A2(n787), .ZN(n788) );
  XNOR2_X1 U873 ( .A(n788), .B(KEYINPUT76), .ZN(n790) );
  NOR2_X1 U874 ( .A1(G299), .A2(G868), .ZN(n789) );
  NOR2_X1 U875 ( .A1(n790), .A2(n789), .ZN(G297) );
  NAND2_X1 U876 ( .A1(n798), .A2(G559), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n791), .A2(n1014), .ZN(n792) );
  XNOR2_X1 U878 ( .A(n792), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U879 ( .A1(G868), .A2(n1025), .ZN(n793) );
  XOR2_X1 U880 ( .A(KEYINPUT77), .B(n793), .Z(n796) );
  NAND2_X1 U881 ( .A1(G868), .A2(n1014), .ZN(n794) );
  NOR2_X1 U882 ( .A1(G559), .A2(n794), .ZN(n795) );
  NOR2_X1 U883 ( .A1(n796), .A2(n795), .ZN(G282) );
  NAND2_X1 U884 ( .A1(n1014), .A2(G559), .ZN(n797) );
  XOR2_X1 U885 ( .A(n1025), .B(n797), .Z(n815) );
  NAND2_X1 U886 ( .A1(n798), .A2(n815), .ZN(n809) );
  NAND2_X1 U887 ( .A1(G55), .A2(n799), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G67), .A2(n800), .ZN(n801) );
  NAND2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n808) );
  NAND2_X1 U890 ( .A1(G93), .A2(n803), .ZN(n806) );
  NAND2_X1 U891 ( .A1(G80), .A2(n804), .ZN(n805) );
  NAND2_X1 U892 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U893 ( .A1(n808), .A2(n807), .ZN(n817) );
  XOR2_X1 U894 ( .A(n809), .B(n817), .Z(G145) );
  XNOR2_X1 U895 ( .A(n1009), .B(KEYINPUT19), .ZN(n811) );
  XNOR2_X1 U896 ( .A(G290), .B(G166), .ZN(n810) );
  XNOR2_X1 U897 ( .A(n811), .B(n810), .ZN(n812) );
  XOR2_X1 U898 ( .A(n817), .B(n812), .Z(n813) );
  XNOR2_X1 U899 ( .A(G305), .B(n813), .ZN(n814) );
  XNOR2_X1 U900 ( .A(n814), .B(G288), .ZN(n866) );
  XNOR2_X1 U901 ( .A(n815), .B(n866), .ZN(n816) );
  NAND2_X1 U902 ( .A1(n816), .A2(G868), .ZN(n819) );
  OR2_X1 U903 ( .A1(G868), .A2(n817), .ZN(n818) );
  NAND2_X1 U904 ( .A1(n819), .A2(n818), .ZN(G295) );
  NAND2_X1 U905 ( .A1(G2084), .A2(G2078), .ZN(n820) );
  XOR2_X1 U906 ( .A(KEYINPUT20), .B(n820), .Z(n821) );
  NAND2_X1 U907 ( .A1(G2090), .A2(n821), .ZN(n823) );
  XOR2_X1 U908 ( .A(KEYINPUT21), .B(KEYINPUT79), .Z(n822) );
  XNOR2_X1 U909 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U910 ( .A1(G2072), .A2(n824), .ZN(G158) );
  XNOR2_X1 U911 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U912 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  NOR2_X1 U913 ( .A1(G219), .A2(G220), .ZN(n826) );
  XNOR2_X1 U914 ( .A(KEYINPUT80), .B(KEYINPUT81), .ZN(n825) );
  XNOR2_X1 U915 ( .A(n826), .B(n825), .ZN(n827) );
  XNOR2_X1 U916 ( .A(KEYINPUT22), .B(n827), .ZN(n828) );
  NOR2_X1 U917 ( .A1(G218), .A2(n828), .ZN(n829) );
  NAND2_X1 U918 ( .A1(G96), .A2(n829), .ZN(n840) );
  NAND2_X1 U919 ( .A1(n840), .A2(G2106), .ZN(n833) );
  NAND2_X1 U920 ( .A1(G69), .A2(G120), .ZN(n830) );
  NOR2_X1 U921 ( .A1(G237), .A2(n830), .ZN(n831) );
  NAND2_X1 U922 ( .A1(G108), .A2(n831), .ZN(n841) );
  NAND2_X1 U923 ( .A1(n841), .A2(G567), .ZN(n832) );
  NAND2_X1 U924 ( .A1(n833), .A2(n832), .ZN(n842) );
  NAND2_X1 U925 ( .A1(G483), .A2(G661), .ZN(n834) );
  NOR2_X1 U926 ( .A1(n842), .A2(n834), .ZN(n839) );
  NAND2_X1 U927 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n835), .ZN(G217) );
  NAND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n836) );
  XOR2_X1 U930 ( .A(KEYINPUT108), .B(n836), .Z(n837) );
  NAND2_X1 U931 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U933 ( .A1(n839), .A2(n838), .ZN(G188) );
  INV_X1 U935 ( .A(G120), .ZN(G236) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  INV_X1 U939 ( .A(n842), .ZN(G319) );
  XOR2_X1 U940 ( .A(G2678), .B(KEYINPUT109), .Z(n844) );
  XNOR2_X1 U941 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U943 ( .A(KEYINPUT42), .B(G2072), .Z(n846) );
  XNOR2_X1 U944 ( .A(G2067), .B(G2090), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U946 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U947 ( .A(G2096), .B(G2100), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U949 ( .A(G2084), .B(G2078), .Z(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U951 ( .A(G1956), .B(G1961), .Z(n854) );
  XNOR2_X1 U952 ( .A(G1986), .B(G1996), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U954 ( .A(G1976), .B(G1971), .Z(n856) );
  XNOR2_X1 U955 ( .A(G1981), .B(G1966), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U957 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U958 ( .A(G2474), .B(KEYINPUT111), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n862) );
  XOR2_X1 U960 ( .A(G1991), .B(KEYINPUT41), .Z(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(G229) );
  XOR2_X1 U962 ( .A(KEYINPUT117), .B(G286), .Z(n865) );
  XNOR2_X1 U963 ( .A(G171), .B(n863), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n868) );
  XOR2_X1 U965 ( .A(n1025), .B(n866), .Z(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n869) );
  NOR2_X1 U967 ( .A1(G37), .A2(n869), .ZN(G397) );
  NAND2_X1 U968 ( .A1(G112), .A2(n892), .ZN(n871) );
  NAND2_X1 U969 ( .A1(G136), .A2(n888), .ZN(n870) );
  NAND2_X1 U970 ( .A1(n871), .A2(n870), .ZN(n877) );
  NAND2_X1 U971 ( .A1(G100), .A2(n889), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n872), .B(KEYINPUT112), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G124), .A2(n893), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n873), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U976 ( .A1(n877), .A2(n876), .ZN(G162) );
  NAND2_X1 U977 ( .A1(G118), .A2(n892), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G130), .A2(n893), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n885) );
  NAND2_X1 U980 ( .A1(n889), .A2(G106), .ZN(n880) );
  XOR2_X1 U981 ( .A(KEYINPUT113), .B(n880), .Z(n882) );
  NAND2_X1 U982 ( .A1(n888), .A2(G142), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  NOR2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n902) );
  NAND2_X1 U987 ( .A1(G139), .A2(n888), .ZN(n891) );
  NAND2_X1 U988 ( .A1(G103), .A2(n889), .ZN(n890) );
  NAND2_X1 U989 ( .A1(n891), .A2(n890), .ZN(n899) );
  NAND2_X1 U990 ( .A1(G115), .A2(n892), .ZN(n895) );
  NAND2_X1 U991 ( .A1(G127), .A2(n893), .ZN(n894) );
  NAND2_X1 U992 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U993 ( .A(KEYINPUT47), .B(n896), .Z(n897) );
  XNOR2_X1 U994 ( .A(KEYINPUT114), .B(n897), .ZN(n898) );
  NOR2_X1 U995 ( .A1(n899), .A2(n898), .ZN(n996) );
  XNOR2_X1 U996 ( .A(n996), .B(G162), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n900), .B(n987), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U999 ( .A(G164), .B(n903), .ZN(n911) );
  XNOR2_X1 U1000 ( .A(G160), .B(n904), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1002 ( .A(n907), .B(KEYINPUT48), .Z(n909) );
  XNOR2_X1 U1003 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1005 ( .A(n911), .B(n910), .Z(n912) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n912), .ZN(n913) );
  XNOR2_X1 U1007 ( .A(KEYINPUT116), .B(n913), .ZN(G395) );
  XNOR2_X1 U1008 ( .A(G2451), .B(G2443), .ZN(n923) );
  XOR2_X1 U1009 ( .A(G2446), .B(KEYINPUT106), .Z(n915) );
  XNOR2_X1 U1010 ( .A(G2438), .B(G2435), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n919) );
  XOR2_X1 U1012 ( .A(KEYINPUT107), .B(G2454), .Z(n917) );
  XNOR2_X1 U1013 ( .A(G1348), .B(G1341), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1015 ( .A(n919), .B(n918), .Z(n921) );
  XNOR2_X1 U1016 ( .A(G2430), .B(G2427), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n921), .B(n920), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(n923), .B(n922), .ZN(n924) );
  NAND2_X1 U1019 ( .A1(n924), .A2(G14), .ZN(n930) );
  NAND2_X1 U1020 ( .A1(G319), .A2(n930), .ZN(n927) );
  NOR2_X1 U1021 ( .A1(G227), .A2(G229), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT49), .B(n925), .ZN(n926) );
  NOR2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n929) );
  NOR2_X1 U1024 ( .A1(G397), .A2(G395), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(G225) );
  INV_X1 U1026 ( .A(G225), .ZN(G308) );
  INV_X1 U1027 ( .A(G96), .ZN(G221) );
  INV_X1 U1028 ( .A(G108), .ZN(G238) );
  INV_X1 U1029 ( .A(n930), .ZN(G401) );
  XOR2_X1 U1030 ( .A(G1348), .B(KEYINPUT59), .Z(n931) );
  XNOR2_X1 U1031 ( .A(G4), .B(n931), .ZN(n940) );
  XOR2_X1 U1032 ( .A(G1341), .B(G19), .Z(n935) );
  XNOR2_X1 U1033 ( .A(G20), .B(n932), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(n933), .B(KEYINPUT126), .ZN(n934) );
  NAND2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(G6), .B(G1981), .ZN(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(n938), .B(KEYINPUT127), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(KEYINPUT60), .B(n941), .ZN(n950) );
  XNOR2_X1 U1041 ( .A(G1966), .B(G21), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G1986), .B(G24), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(G1971), .B(G22), .ZN(n942) );
  NOR2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n945) );
  XOR2_X1 U1045 ( .A(G1976), .B(G23), .Z(n944) );
  NAND2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1047 ( .A(KEYINPUT58), .B(n946), .ZN(n947) );
  NOR2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(G5), .B(G1961), .ZN(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1052 ( .A(KEYINPUT61), .B(n953), .Z(n955) );
  XOR2_X1 U1053 ( .A(G16), .B(KEYINPUT125), .Z(n954) );
  NOR2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n978) );
  INV_X1 U1055 ( .A(KEYINPUT55), .ZN(n1004) );
  XNOR2_X1 U1056 ( .A(G2090), .B(G35), .ZN(n969) );
  XNOR2_X1 U1057 ( .A(G1991), .B(G25), .ZN(n957) );
  XNOR2_X1 U1058 ( .A(G32), .B(G1996), .ZN(n956) );
  NOR2_X1 U1059 ( .A1(n957), .A2(n956), .ZN(n963) );
  XOR2_X1 U1060 ( .A(G2072), .B(G33), .Z(n958) );
  NAND2_X1 U1061 ( .A1(n958), .A2(G28), .ZN(n961) );
  XOR2_X1 U1062 ( .A(KEYINPUT121), .B(G2067), .Z(n959) );
  XNOR2_X1 U1063 ( .A(G26), .B(n959), .ZN(n960) );
  NOR2_X1 U1064 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1065 ( .A1(n963), .A2(n962), .ZN(n966) );
  XNOR2_X1 U1066 ( .A(G27), .B(n964), .ZN(n965) );
  NOR2_X1 U1067 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1068 ( .A(KEYINPUT53), .B(n967), .ZN(n968) );
  NOR2_X1 U1069 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1070 ( .A(G2084), .B(G34), .Z(n970) );
  XNOR2_X1 U1071 ( .A(KEYINPUT54), .B(n970), .ZN(n971) );
  NAND2_X1 U1072 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1073 ( .A(n1004), .B(n973), .ZN(n975) );
  INV_X1 U1074 ( .A(G29), .ZN(n974) );
  NAND2_X1 U1075 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1076 ( .A1(G11), .A2(n976), .ZN(n977) );
  NOR2_X1 U1077 ( .A1(n978), .A2(n977), .ZN(n1008) );
  XOR2_X1 U1078 ( .A(G2090), .B(G162), .Z(n979) );
  NOR2_X1 U1079 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1080 ( .A(KEYINPUT51), .B(n981), .ZN(n982) );
  XNOR2_X1 U1081 ( .A(n982), .B(KEYINPUT119), .ZN(n995) );
  NOR2_X1 U1082 ( .A1(n984), .A2(n983), .ZN(n986) );
  NAND2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(G160), .B(G2084), .ZN(n988) );
  NAND2_X1 U1085 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1086 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1087 ( .A(KEYINPUT118), .B(n991), .Z(n992) );
  NOR2_X1 U1088 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1089 ( .A1(n995), .A2(n994), .ZN(n1002) );
  XOR2_X1 U1090 ( .A(G2072), .B(n996), .Z(n998) );
  XOR2_X1 U1091 ( .A(G164), .B(G2078), .Z(n997) );
  NOR2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1093 ( .A(KEYINPUT50), .B(n999), .Z(n1000) );
  XNOR2_X1 U1094 ( .A(KEYINPUT120), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1096 ( .A(KEYINPUT52), .B(n1003), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1006), .A2(G29), .ZN(n1007) );
  NAND2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1037) );
  XOR2_X1 U1100 ( .A(KEYINPUT56), .B(G16), .Z(n1035) );
  XNOR2_X1 U1101 ( .A(n1009), .B(G1956), .ZN(n1011) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(G1348), .B(KEYINPUT122), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(n1015), .B(n1014), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1032) );
  XOR2_X1 U1107 ( .A(G168), .B(G1966), .Z(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1109 ( .A(KEYINPUT57), .B(n1020), .Z(n1030) );
  XOR2_X1 U1110 ( .A(G171), .B(G1961), .Z(n1022) );
  XOR2_X1 U1111 ( .A(G166), .B(G1971), .Z(n1021) );
  NOR2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  NAND2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1028) );
  XOR2_X1 U1114 ( .A(G1341), .B(n1025), .Z(n1026) );
  XNOR2_X1 U1115 ( .A(KEYINPUT123), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1118 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1119 ( .A(KEYINPUT124), .B(n1033), .ZN(n1034) );
  NOR2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NOR2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XNOR2_X1 U1122 ( .A(n1038), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

