//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XOR2_X1   g001(.A(G78gat), .B(G106gat), .Z(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT31), .B(G50gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G141gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G148gat), .ZN(new_n207));
  INV_X1    g006(.A(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G141gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n211));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n210), .A2(new_n211), .B1(KEYINPUT2), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G141gat), .B(G148gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT79), .ZN(new_n215));
  INV_X1    g014(.A(new_n212), .ZN(new_n216));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT78), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n217), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT78), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(new_n212), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n213), .A2(new_n215), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT80), .B(G148gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n207), .B1(new_n223), .B2(new_n206), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n212), .B1(new_n219), .B2(KEYINPUT2), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT29), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(G211gat), .B(G218gat), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT76), .ZN(new_n231));
  XNOR2_X1  g030(.A(G197gat), .B(G204gat), .ZN(new_n232));
  INV_X1    g031(.A(G211gat), .ZN(new_n233));
  INV_X1    g032(.A(G218gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n232), .B1(KEYINPUT22), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n231), .B(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT85), .B1(new_n229), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G228gat), .ZN(new_n240));
  INV_X1    g039(.A(G233gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT85), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n221), .A2(new_n218), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n212), .A2(KEYINPUT2), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n214), .B2(KEYINPUT79), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n210), .A2(new_n211), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n244), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n224), .A2(new_n225), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n243), .B(new_n237), .C1(new_n251), .C2(KEYINPUT29), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n228), .B1(new_n237), .B2(KEYINPUT29), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT81), .B1(new_n248), .B2(new_n249), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n248), .A2(KEYINPUT81), .A3(new_n249), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n239), .A2(new_n242), .A3(new_n252), .A4(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n229), .A2(new_n238), .ZN(new_n258));
  INV_X1    g057(.A(new_n230), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT29), .B1(new_n236), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n259), .B2(new_n236), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n227), .B1(new_n228), .B2(new_n261), .ZN(new_n262));
  OAI22_X1  g061(.A1(new_n258), .A2(new_n262), .B1(new_n240), .B2(new_n241), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G22gat), .ZN(new_n265));
  INV_X1    g064(.A(G22gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n257), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n265), .A2(KEYINPUT86), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT86), .B1(new_n265), .B2(new_n267), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n205), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n269), .A2(new_n205), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR3_X1   g075(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n277));
  OAI211_X1 g076(.A(KEYINPUT69), .B(new_n273), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT26), .ZN(new_n280));
  INV_X1    g079(.A(G169gat), .ZN(new_n281));
  INV_X1    g080(.A(G176gat), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(new_n275), .A3(new_n274), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT69), .B1(new_n284), .B2(new_n273), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n287));
  INV_X1    g086(.A(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT65), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G190gat), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n287), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT27), .B(G183gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(KEYINPUT68), .A3(new_n293), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT27), .ZN(new_n301));
  INV_X1    g100(.A(G183gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n301), .B1(new_n302), .B2(KEYINPUT66), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n304), .A2(KEYINPUT64), .A3(KEYINPUT27), .A4(G183gat), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n303), .B(new_n305), .C1(KEYINPUT64), .C2(G183gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n300), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n286), .B1(new_n298), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n273), .B(KEYINPUT24), .ZN(new_n310));
  INV_X1    g109(.A(new_n307), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT64), .B(G183gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n281), .A2(new_n282), .A3(KEYINPUT23), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n315), .B1(G169gat), .B2(G176gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n316), .A3(new_n275), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n288), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n317), .A2(KEYINPUT25), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n319), .A2(KEYINPUT25), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n309), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT72), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT70), .ZN(new_n326));
  INV_X1    g125(.A(G127gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(G134gat), .ZN(new_n328));
  INV_X1    g127(.A(G134gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n328), .B(new_n330), .C1(G127gat), .C2(new_n329), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT1), .ZN(new_n332));
  INV_X1    g131(.A(G113gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(G120gat), .ZN(new_n334));
  INV_X1    g133(.A(G120gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(G113gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n332), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT71), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n333), .B2(G120gat), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n333), .A2(G120gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n335), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n332), .B1(new_n329), .B2(G127gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n327), .A2(G134gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n331), .A2(new_n337), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT72), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n309), .A2(new_n323), .A3(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n325), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(G227gat), .A2(G233gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n324), .A2(KEYINPUT72), .A3(new_n346), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT32), .ZN(new_n355));
  XOR2_X1   g154(.A(G15gat), .B(G43gat), .Z(new_n356));
  XNOR2_X1  g155(.A(G71gat), .B(G99gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n355), .B1(KEYINPUT33), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT33), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT73), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT73), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n354), .A2(new_n363), .A3(new_n360), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n355), .A2(new_n358), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n359), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n351), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT34), .B1(new_n352), .B2(KEYINPUT74), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n372), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n366), .B1(new_n362), .B2(new_n364), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n374), .B1(new_n375), .B2(new_n359), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT77), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n273), .B1(new_n276), .B2(new_n277), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT69), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n278), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n292), .A2(KEYINPUT68), .A3(new_n293), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT68), .B1(new_n292), .B2(new_n293), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n306), .A2(new_n307), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n299), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n381), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n322), .A2(new_n321), .ZN(new_n388));
  INV_X1    g187(.A(new_n312), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n307), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n317), .B1(new_n390), .B2(new_n310), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT25), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n377), .B1(new_n387), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n309), .A2(new_n323), .A3(KEYINPUT77), .ZN(new_n395));
  INV_X1    g194(.A(G226gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(new_n241), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(KEYINPUT29), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n387), .A2(new_n393), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n397), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n238), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n387), .A2(new_n393), .A3(new_n377), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT77), .B1(new_n309), .B2(new_n323), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n397), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n324), .A2(new_n398), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(new_n237), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G8gat), .B(G36gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(G64gat), .B(G92gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n412), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n403), .A2(new_n408), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n415), .A3(KEYINPUT30), .ZN(new_n416));
  OR3_X1    g215(.A1(new_n409), .A2(KEYINPUT30), .A3(new_n412), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n272), .A2(new_n373), .A3(new_n376), .A4(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n248), .A2(new_n346), .A3(new_n249), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT4), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n248), .A2(new_n346), .A3(new_n249), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n222), .B2(new_n226), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n248), .A2(KEYINPUT81), .A3(new_n249), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n228), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n347), .B1(new_n250), .B2(KEYINPUT3), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n421), .B(new_n426), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(new_n421), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n346), .B1(new_n428), .B2(new_n429), .ZN(new_n434));
  INV_X1    g233(.A(new_n422), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n432), .A2(KEYINPUT5), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT82), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT5), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n347), .B1(new_n255), .B2(new_n254), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n422), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n440), .B1(new_n442), .B2(new_n433), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(KEYINPUT82), .A3(new_n432), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT83), .B1(new_n432), .B2(KEYINPUT5), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT3), .B1(new_n255), .B2(new_n254), .ZN(new_n446));
  INV_X1    g245(.A(new_n431), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n446), .A2(new_n447), .B1(new_n423), .B2(new_n425), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT83), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n440), .A4(new_n421), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n439), .A2(new_n444), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G1gat), .B(G29gat), .ZN(new_n452));
  INV_X1    g251(.A(G85gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT0), .B(G57gat), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n454), .B(new_n455), .Z(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n420), .B1(new_n451), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n450), .A2(new_n445), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT82), .B1(new_n443), .B2(new_n432), .ZN(new_n460));
  AND4_X1   g259(.A1(KEYINPUT82), .A2(new_n432), .A3(KEYINPUT5), .A4(new_n436), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n459), .B(new_n457), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT88), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT6), .B1(new_n465), .B2(new_n456), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT88), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(new_n462), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n451), .A2(new_n420), .A3(new_n457), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n464), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n202), .B1(new_n419), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT40), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n448), .A2(new_n421), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT39), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n456), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n441), .A2(new_n421), .A3(new_n422), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT39), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT87), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT87), .B1(new_n478), .B2(KEYINPUT39), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n481), .A2(new_n482), .A3(new_n474), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n473), .B1(new_n477), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n456), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n477), .A2(new_n483), .A3(new_n473), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n418), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n403), .A2(new_n489), .A3(new_n408), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT90), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n403), .A2(new_n492), .A3(new_n408), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n414), .A2(KEYINPUT38), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n399), .A2(new_n237), .A3(new_n401), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT89), .ZN(new_n497));
  INV_X1    g296(.A(new_n397), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n498), .B1(new_n394), .B2(new_n395), .ZN(new_n499));
  INV_X1    g298(.A(new_n407), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n238), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n399), .A2(new_n502), .A3(new_n237), .A4(new_n401), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n497), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n495), .B1(new_n504), .B2(KEYINPUT37), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n494), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n415), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n489), .B1(new_n403), .B2(new_n408), .ZN(new_n508));
  OR3_X1    g307(.A1(new_n508), .A2(KEYINPUT91), .A3(new_n414), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT91), .B1(new_n508), .B2(new_n414), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n509), .A2(new_n494), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n507), .B1(KEYINPUT38), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n488), .B1(new_n512), .B2(new_n471), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT75), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n374), .B1(new_n368), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(KEYINPUT75), .B(new_n372), .C1(new_n375), .C2(new_n359), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(KEYINPUT36), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n373), .A2(new_n376), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n272), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n472), .B1(new_n513), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT84), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n469), .B1(new_n462), .B2(new_n466), .ZN(new_n523));
  INV_X1    g322(.A(new_n418), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n466), .A2(new_n462), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n470), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(KEYINPUT84), .A3(new_n418), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n272), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n517), .A2(new_n530), .A3(new_n519), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(KEYINPUT35), .A3(new_n272), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n529), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n521), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G85gat), .A2(G92gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g336(.A1(G99gat), .A2(G106gat), .ZN(new_n538));
  INV_X1    g337(.A(G92gat), .ZN(new_n539));
  AOI22_X1  g338(.A1(KEYINPUT8), .A2(new_n538), .B1(new_n453), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(G99gat), .B(G106gat), .Z(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n543), .A2(KEYINPUT97), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(KEYINPUT97), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n541), .A2(new_n542), .ZN(new_n546));
  NOR3_X1   g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OR3_X1    g346(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n549));
  AOI22_X1  g348(.A1(new_n548), .A2(new_n549), .B1(G29gat), .B2(G36gat), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n551));
  XNOR2_X1  g350(.A(G43gat), .B(G50gat), .ZN(new_n552));
  OR2_X1    g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n552), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n547), .B1(KEYINPUT17), .B2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n556), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n558), .A2(new_n547), .B1(KEYINPUT41), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G134gat), .B(G162gat), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n562), .A2(KEYINPUT41), .ZN(new_n567));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n566), .A2(new_n570), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G57gat), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n575), .A2(G64gat), .ZN(new_n576));
  AND2_X1   g375(.A1(KEYINPUT94), .A2(G64gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(KEYINPUT94), .A2(G64gat), .ZN(new_n578));
  OAI21_X1  g377(.A(G57gat), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n576), .B1(new_n579), .B2(KEYINPUT95), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(KEYINPUT95), .B2(new_n579), .ZN(new_n581));
  INV_X1    g380(.A(G71gat), .ZN(new_n582));
  INV_X1    g381(.A(G78gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT9), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n581), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT93), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n584), .B1(new_n589), .B2(new_n585), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n575), .A2(G64gat), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT9), .B1(new_n576), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n590), .B(new_n592), .C1(new_n589), .C2(new_n585), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G127gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G155gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(new_n302), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(new_n233), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n598), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G15gat), .B(G22gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT16), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(new_n604), .B2(G1gat), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(G1gat), .B2(new_n603), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G8gat), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n607), .B1(new_n594), .B2(KEYINPUT21), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n602), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n602), .A2(new_n610), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n574), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n535), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n547), .A2(new_n594), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n542), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n541), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n615), .B1(new_n594), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT10), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n547), .A2(new_n594), .A3(KEYINPUT10), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G230gat), .A2(G233gat), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n619), .A2(new_n624), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G176gat), .B(G204gat), .Z(new_n628));
  XNOR2_X1  g427(.A(G120gat), .B(G148gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(KEYINPUT99), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT99), .B1(new_n627), .B2(new_n630), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n630), .B(KEYINPUT100), .Z(new_n634));
  OAI22_X1  g433(.A1(new_n632), .A2(new_n633), .B1(new_n627), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n607), .B1(new_n556), .B2(KEYINPUT17), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n560), .A2(new_n636), .B1(new_n607), .B2(new_n558), .ZN(new_n637));
  NAND2_X1  g436(.A1(G229gat), .A2(G233gat), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n639), .A2(KEYINPUT18), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(KEYINPUT18), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n556), .B(new_n607), .Z(new_n642));
  XOR2_X1   g441(.A(new_n638), .B(KEYINPUT13), .Z(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n640), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G113gat), .B(G141gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G197gat), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT11), .B(G169gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT12), .Z(new_n650));
  OR2_X1    g449(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n645), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n635), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n614), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n527), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT101), .B(G1gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1324gat));
  NOR2_X1   g458(.A1(new_n656), .A2(new_n418), .ZN(new_n660));
  INV_X1    g459(.A(G8gat), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT42), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT16), .B(G8gat), .Z(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  MUX2_X1   g463(.A(KEYINPUT42), .B(new_n662), .S(new_n664), .Z(G1325gat));
  INV_X1    g464(.A(G15gat), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n517), .A2(new_n519), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n656), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n373), .A2(new_n376), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n656), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n669), .B1(new_n666), .B2(new_n671), .ZN(G1326gat));
  NOR2_X1   g471(.A1(new_n656), .A2(new_n272), .ZN(new_n673));
  XOR2_X1   g472(.A(KEYINPUT43), .B(G22gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  NAND2_X1  g474(.A1(new_n611), .A2(new_n612), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n676), .A2(new_n635), .A3(new_n654), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n535), .A2(new_n574), .A3(new_n677), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n678), .A2(G29gat), .A3(new_n527), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT45), .Z(new_n680));
  OAI21_X1  g479(.A(new_n574), .B1(new_n521), .B2(new_n534), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT44), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n683), .B(new_n574), .C1(new_n521), .C2(new_n534), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n676), .B(KEYINPUT102), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n655), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT103), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n690));
  AOI211_X1 g489(.A(new_n690), .B(new_n687), .C1(new_n682), .C2(new_n684), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n692), .B2(new_n527), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n680), .A2(new_n693), .ZN(G1328gat));
  OAI21_X1  g493(.A(G36gat), .B1(new_n692), .B2(new_n418), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n418), .A2(G36gat), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n678), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT104), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n698), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT105), .B1(new_n698), .B2(KEYINPUT46), .ZN(new_n700));
  OAI221_X1 g499(.A(new_n695), .B1(KEYINPUT46), .B2(new_n698), .C1(new_n699), .C2(new_n700), .ZN(G1329gat));
  INV_X1    g500(.A(G43gat), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n687), .B1(new_n682), .B2(new_n684), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n702), .B1(new_n703), .B2(new_n667), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n670), .A2(G43gat), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT47), .B1(new_n678), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(KEYINPUT107), .B1(new_n704), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n707), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710));
  AOI211_X1 g509(.A(new_n668), .B(new_n687), .C1(new_n682), .C2(new_n684), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n709), .B(new_n710), .C1(new_n711), .C2(new_n702), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n678), .A2(KEYINPUT106), .A3(new_n706), .ZN(new_n714));
  OAI21_X1  g513(.A(KEYINPUT106), .B1(new_n678), .B2(new_n706), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n667), .B1(new_n689), .B2(new_n691), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(G43gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n713), .B1(new_n718), .B2(KEYINPUT47), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(KEYINPUT108), .B(new_n713), .C1(new_n718), .C2(KEYINPUT47), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1330gat));
  NOR2_X1   g522(.A1(new_n272), .A2(G50gat), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n678), .B2(KEYINPUT109), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(KEYINPUT109), .B2(new_n678), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n530), .B1(new_n689), .B2(new_n691), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(G50gat), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(G50gat), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n703), .B2(new_n530), .ZN(new_n732));
  OAI22_X1  g531(.A1(KEYINPUT48), .A2(new_n728), .B1(new_n730), .B2(new_n732), .ZN(G1331gat));
  NOR2_X1   g532(.A1(new_n627), .A2(new_n634), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n627), .A2(new_n630), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT99), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n734), .B1(new_n737), .B2(new_n631), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n653), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n535), .A2(new_n613), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n527), .ZN(new_n741));
  XNOR2_X1  g540(.A(KEYINPUT110), .B(G57gat), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1332gat));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n740), .B(new_n744), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n745), .A2(new_n524), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  AND2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n746), .B2(new_n747), .ZN(G1333gat));
  OR3_X1    g549(.A1(new_n740), .A2(KEYINPUT113), .A3(new_n670), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT113), .B1(new_n740), .B2(new_n670), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(new_n582), .A3(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n668), .A2(new_n582), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n745), .A2(KEYINPUT112), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(KEYINPUT112), .B1(new_n745), .B2(new_n754), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n753), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g557(.A1(new_n745), .A2(new_n530), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G78gat), .ZN(G1335gat));
  INV_X1    g559(.A(new_n681), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n676), .A2(new_n653), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT51), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n761), .A2(KEYINPUT51), .A3(new_n762), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(KEYINPUT114), .A3(new_n766), .ZN(new_n767));
  OR3_X1    g566(.A1(new_n763), .A2(KEYINPUT114), .A3(new_n764), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n635), .A2(new_n453), .A3(new_n523), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n676), .A2(new_n738), .A3(new_n653), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n685), .A2(new_n523), .A3(new_n771), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n769), .A2(new_n770), .B1(new_n453), .B2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT115), .ZN(G1336gat));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n765), .A2(new_n775), .A3(new_n766), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n738), .A2(G92gat), .A3(new_n418), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n763), .A2(KEYINPUT116), .A3(new_n764), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n685), .A2(new_n524), .A3(new_n771), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G92gat), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT52), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n767), .A2(new_n768), .A3(new_n777), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n783), .A2(new_n786), .ZN(G1337gat));
  NAND3_X1  g586(.A1(new_n685), .A2(new_n667), .A3(new_n771), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G99gat), .ZN(new_n789));
  OR3_X1    g588(.A1(new_n738), .A2(G99gat), .A3(new_n670), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n769), .B2(new_n790), .ZN(G1338gat));
  NOR3_X1   g590(.A1(new_n738), .A2(G106gat), .A3(new_n272), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n776), .A2(new_n778), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n685), .A2(new_n530), .A3(new_n771), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G106gat), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT53), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n767), .A2(new_n768), .A3(new_n792), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n799), .A3(new_n795), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n797), .A2(new_n800), .ZN(G1339gat));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n738), .A2(new_n654), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n802), .B1(new_n804), .B2(new_n613), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n676), .A2(new_n573), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n806), .A2(new_n803), .A3(KEYINPUT118), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n637), .A2(new_n638), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n642), .A2(new_n643), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n649), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n651), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n635), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n737), .A2(new_n631), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n630), .B1(new_n625), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g616(.A1(new_n623), .A2(new_n624), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n623), .A2(new_n624), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(KEYINPUT54), .A3(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT55), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n817), .A2(new_n820), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n815), .A2(new_n822), .A3(new_n653), .A4(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n574), .B1(new_n814), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n815), .A2(new_n822), .ZN(new_n828));
  INV_X1    g627(.A(new_n825), .ZN(new_n829));
  NOR4_X1   g628(.A1(new_n828), .A2(new_n573), .A3(new_n829), .A4(new_n812), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n686), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n530), .B(new_n670), .C1(new_n808), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n527), .A2(new_n524), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n654), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n532), .A2(new_n272), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n808), .B2(new_n831), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(new_n833), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n333), .A3(new_n653), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n835), .A2(new_n839), .ZN(G1340gat));
  OAI21_X1  g639(.A(G120gat), .B1(new_n834), .B2(new_n738), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n838), .A2(new_n335), .A3(new_n635), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1341gat));
  NOR3_X1   g642(.A1(new_n834), .A2(new_n327), .A3(new_n686), .ZN(new_n844));
  AOI21_X1  g643(.A(G127gat), .B1(new_n838), .B2(new_n676), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(G1342gat));
  OAI21_X1  g645(.A(G134gat), .B1(new_n834), .B2(new_n573), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n527), .B1(new_n808), .B2(new_n831), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n530), .B1(new_n516), .B2(new_n515), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n573), .A2(new_n524), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n848), .A2(new_n329), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT56), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(new_n851), .B2(KEYINPUT56), .ZN(new_n854));
  OAI221_X1 g653(.A(new_n847), .B1(KEYINPUT56), .B2(new_n851), .C1(new_n853), .C2(new_n854), .ZN(G1343gat));
  NAND2_X1  g654(.A1(KEYINPUT123), .A2(KEYINPUT58), .ZN(new_n856));
  INV_X1    g655(.A(new_n531), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n848), .A2(new_n857), .A3(new_n418), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n653), .A2(new_n206), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT121), .B1(new_n738), .B2(new_n812), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n823), .A2(KEYINPUT122), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n823), .A2(KEYINPUT122), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT55), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n815), .A2(new_n822), .A3(new_n653), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n814), .A2(KEYINPUT121), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n573), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n830), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n676), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n808), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n530), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT57), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n272), .B1(new_n808), .B2(new_n831), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT57), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n668), .A2(new_n833), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT120), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n873), .A2(new_n653), .A3(new_n876), .A4(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n860), .B1(new_n879), .B2(G141gat), .ZN(new_n880));
  NOR2_X1   g679(.A1(KEYINPUT123), .A2(KEYINPUT58), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n880), .B(new_n881), .ZN(G1344gat));
  OR3_X1    g681(.A1(new_n858), .A2(new_n223), .A3(new_n738), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n874), .A2(new_n875), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n806), .A2(new_n803), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n875), .B(new_n530), .C1(new_n870), .C2(new_n886), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n635), .A3(new_n878), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n884), .B1(new_n889), .B2(G148gat), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n223), .A2(new_n884), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n873), .A2(new_n876), .A3(new_n878), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n635), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n883), .B1(new_n890), .B2(new_n893), .ZN(G1345gat));
  NAND2_X1  g693(.A1(new_n848), .A2(new_n857), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n895), .A2(new_n524), .ZN(new_n896));
  AOI21_X1  g695(.A(G155gat), .B1(new_n896), .B2(new_n676), .ZN(new_n897));
  INV_X1    g696(.A(G155gat), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n686), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n897), .B1(new_n892), .B2(new_n899), .ZN(G1346gat));
  AND2_X1   g699(.A1(new_n892), .A2(new_n574), .ZN(new_n901));
  INV_X1    g700(.A(G162gat), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n850), .A2(new_n902), .ZN(new_n903));
  OAI22_X1  g702(.A1(new_n901), .A2(new_n902), .B1(new_n895), .B2(new_n903), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n523), .A2(new_n418), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n832), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G169gat), .B1(new_n906), .B2(new_n654), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n837), .A2(new_n905), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n653), .A2(new_n281), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(G1348gat));
  NOR3_X1   g709(.A1(new_n906), .A2(new_n282), .A3(new_n738), .ZN(new_n911));
  INV_X1    g710(.A(new_n908), .ZN(new_n912));
  AOI21_X1  g711(.A(G176gat), .B1(new_n912), .B2(new_n635), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n911), .A2(new_n913), .ZN(G1349gat));
  OAI21_X1  g713(.A(new_n312), .B1(new_n906), .B2(new_n686), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n912), .A2(new_n676), .A3(new_n293), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(KEYINPUT124), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n912), .A2(new_n574), .A3(new_n307), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT125), .ZN(new_n920));
  OAI21_X1  g719(.A(G190gat), .B1(new_n906), .B2(new_n573), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT61), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(KEYINPUT61), .B2(new_n921), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n922), .B1(new_n921), .B2(KEYINPUT61), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(G1351gat));
  NAND2_X1  g725(.A1(new_n668), .A2(new_n905), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n888), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n653), .ZN(new_n930));
  XOR2_X1   g729(.A(KEYINPUT127), .B(G197gat), .Z(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n874), .A2(new_n928), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n654), .A2(new_n931), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n932), .A2(new_n935), .ZN(G1352gat));
  INV_X1    g735(.A(G204gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n937), .A3(new_n635), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT62), .Z(new_n939));
  AND3_X1   g738(.A1(new_n888), .A2(new_n635), .A3(new_n928), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n937), .B2(new_n940), .ZN(G1353gat));
  NAND3_X1  g740(.A1(new_n933), .A2(new_n233), .A3(new_n676), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n888), .A2(new_n676), .A3(new_n928), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n943), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT63), .B1(new_n943), .B2(G211gat), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1354gat));
  AOI21_X1  g745(.A(G218gat), .B1(new_n933), .B2(new_n574), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n573), .A2(new_n234), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n929), .B2(new_n948), .ZN(G1355gat));
endmodule


