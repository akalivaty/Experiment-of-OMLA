//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n626, new_n627, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(G104), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT71), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G953), .ZN(new_n193));
  INV_X1    g007(.A(G237), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n191), .A2(new_n193), .A3(G214), .A4(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(G143), .A2(G214), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n191), .A2(new_n193), .A3(new_n198), .A4(new_n194), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT18), .A2(G131), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n197), .A2(KEYINPUT18), .A3(G131), .A4(new_n199), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  INV_X1    g019(.A(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G140), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT76), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT75), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n205), .A2(new_n207), .A3(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n206), .A2(KEYINPUT75), .A3(G140), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(G146), .A3(new_n214), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n202), .A2(new_n203), .B1(new_n211), .B2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n200), .A2(KEYINPUT17), .A3(G131), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(KEYINPUT16), .A3(new_n214), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n205), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n208), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n208), .A3(new_n220), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n217), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT86), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n195), .A2(new_n196), .ZN(new_n226));
  INV_X1    g040(.A(G131), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n199), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n225), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n200), .A2(G131), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT17), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n197), .A2(KEYINPUT86), .A3(new_n227), .A4(new_n199), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n229), .A2(new_n230), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  AOI211_X1 g047(.A(new_n189), .B(new_n216), .C1(new_n224), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n189), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n229), .A2(new_n230), .A3(new_n232), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n213), .A2(KEYINPUT19), .A3(new_n214), .ZN(new_n237));
  XNOR2_X1  g051(.A(G125), .B(G140), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT19), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT87), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AND4_X1   g054(.A1(KEYINPUT87), .A2(new_n205), .A3(new_n207), .A4(new_n239), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n237), .B(new_n208), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT88), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT87), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n205), .A2(new_n207), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(KEYINPUT19), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n238), .A2(KEYINPUT87), .A3(new_n239), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT88), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n248), .A2(new_n249), .A3(new_n208), .A4(new_n237), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n236), .A2(new_n222), .A3(new_n243), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n216), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n235), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n187), .B1(new_n234), .B2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(G475), .A2(G902), .ZN(new_n255));
  INV_X1    g069(.A(new_n233), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n217), .A2(new_n222), .A3(new_n223), .ZN(new_n257));
  OAI211_X1 g071(.A(new_n235), .B(new_n252), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n243), .A2(new_n222), .A3(new_n250), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n216), .B1(new_n259), .B2(new_n236), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n258), .B(KEYINPUT89), .C1(new_n260), .C2(new_n235), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n254), .A2(new_n255), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT20), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT90), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT90), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n265), .A3(KEYINPUT20), .ZN(new_n266));
  NOR3_X1   g080(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n234), .B2(new_n253), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G475), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n252), .B1(new_n256), .B2(new_n257), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n189), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n258), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G107), .ZN(new_n277));
  INV_X1    g091(.A(G116), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n278), .A2(G122), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n279), .B2(KEYINPUT14), .ZN(new_n280));
  XNOR2_X1  g094(.A(G116), .B(G122), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G128), .B(G143), .ZN(new_n283));
  XOR2_X1   g097(.A(new_n283), .B(KEYINPUT91), .Z(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(G134), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n283), .B(KEYINPUT91), .ZN(new_n286));
  INV_X1    g100(.A(G134), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n282), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n283), .A2(KEYINPUT13), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n196), .A2(G128), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n290), .B(G134), .C1(KEYINPUT13), .C2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n281), .B(new_n277), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n292), .B(new_n293), .C1(new_n284), .C2(G134), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT9), .B(G234), .ZN(new_n295));
  INV_X1    g109(.A(G217), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n295), .A2(new_n296), .A3(G953), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n289), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n289), .B2(new_n294), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n274), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G478), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n301), .A2(KEYINPUT15), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OAI221_X1 g117(.A(new_n274), .B1(KEYINPUT15), .B2(new_n301), .C1(new_n298), .C2(new_n299), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G952), .ZN(new_n306));
  AOI211_X1 g120(.A(G953), .B(new_n306), .C1(G234), .C2(G237), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n191), .A2(new_n193), .ZN(new_n308));
  AOI211_X1 g122(.A(new_n274), .B(new_n308), .C1(G234), .C2(G237), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT21), .B(G898), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n269), .A2(new_n276), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT92), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT92), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n269), .A2(new_n312), .A3(new_n315), .A4(new_n276), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT68), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n318), .B1(new_n278), .B2(G119), .ZN(new_n319));
  INV_X1    g133(.A(G119), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT68), .A3(G116), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n278), .A2(G119), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G113), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT2), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT2), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G113), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(new_n327), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n330), .A2(new_n319), .A3(new_n321), .A4(new_n322), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n329), .A2(new_n331), .A3(KEYINPUT69), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT69), .B1(new_n329), .B2(new_n331), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n196), .A2(G146), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT64), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n208), .B2(G143), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n196), .A2(KEYINPUT64), .A3(G146), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n335), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(KEYINPUT0), .A2(G128), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OR2_X1    g155(.A1(KEYINPUT0), .A2(G128), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n342), .A2(new_n340), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n208), .A2(G143), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n196), .A2(G146), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n339), .A2(new_n341), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT65), .ZN(new_n350));
  INV_X1    g164(.A(G137), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G134), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT11), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n351), .A2(KEYINPUT11), .A3(G134), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n287), .A2(G137), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT11), .B1(new_n351), .B2(G134), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n350), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n349), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n355), .B(new_n356), .C1(new_n359), .C2(new_n350), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n353), .B1(new_n287), .B2(G137), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(KEYINPUT65), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n362), .A2(new_n348), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n347), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n337), .A2(new_n338), .ZN(new_n367));
  INV_X1    g181(.A(G128), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(KEYINPUT1), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n344), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G128), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n346), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n375));
  XNOR2_X1  g189(.A(G134), .B(G137), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(new_n227), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n352), .A2(new_n356), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(KEYINPUT67), .A3(G131), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n357), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n363), .A2(KEYINPUT65), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n381), .A2(new_n360), .A3(new_n382), .A4(new_n227), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n374), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n334), .A2(new_n366), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(KEYINPUT28), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT70), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n329), .A2(new_n331), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n374), .A2(new_n380), .A3(new_n383), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n196), .A2(KEYINPUT64), .A3(G146), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT64), .B1(new_n196), .B2(G146), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n341), .B(new_n344), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n346), .A2(new_n340), .A3(new_n342), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n348), .B1(new_n362), .B2(new_n364), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n381), .A2(new_n360), .A3(new_n382), .A4(new_n349), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n390), .B1(new_n391), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT73), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n334), .A2(new_n366), .A3(KEYINPUT70), .A4(new_n384), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT73), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n403), .B(new_n390), .C1(new_n391), .C2(new_n399), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n389), .A2(new_n401), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n406));
  AOI211_X1 g220(.A(KEYINPUT29), .B(new_n387), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n408));
  OAI22_X1  g222(.A1(new_n391), .A2(new_n399), .B1(new_n333), .B2(new_n332), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n389), .A2(new_n402), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT28), .ZN(new_n411));
  INV_X1    g225(.A(new_n387), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n308), .A2(G210), .A3(new_n194), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT27), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT26), .B(G101), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n407), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n389), .A2(new_n402), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n391), .A2(new_n399), .A3(KEYINPUT30), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT30), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n366), .B2(new_n384), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n390), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(new_n418), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n274), .B1(new_n425), .B2(KEYINPUT29), .ZN(new_n426));
  OAI21_X1  g240(.A(G472), .B1(new_n419), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G472), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n424), .A2(new_n389), .A3(new_n402), .A4(new_n417), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT31), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT31), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n420), .A2(new_n431), .A3(new_n417), .A4(new_n424), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n405), .A2(new_n406), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n417), .B1(new_n434), .B2(new_n412), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n428), .B(new_n274), .C1(new_n433), .C2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT32), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n387), .B1(new_n405), .B2(new_n406), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n430), .B(new_n432), .C1(new_n439), .C2(new_n417), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n440), .A2(KEYINPUT32), .A3(new_n428), .A4(new_n274), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n427), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n308), .A2(G221), .A3(G234), .ZN(new_n443));
  XOR2_X1   g257(.A(KEYINPUT22), .B(G137), .Z(new_n444));
  XNOR2_X1  g258(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n445), .B(new_n446), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT24), .B(G110), .Z(new_n448));
  XNOR2_X1  g262(.A(G119), .B(G128), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT74), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT23), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n320), .B2(G128), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n368), .A2(KEYINPUT23), .A3(G119), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n453), .B(new_n454), .C1(G119), .C2(new_n368), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G110), .ZN(new_n456));
  INV_X1    g270(.A(new_n223), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n451), .B(new_n456), .C1(new_n457), .C2(new_n221), .ZN(new_n458));
  OAI22_X1  g272(.A1(new_n455), .A2(G110), .B1(new_n449), .B2(new_n448), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n222), .A2(new_n211), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n447), .B(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n296), .B1(G234), .B2(new_n274), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(G902), .ZN(new_n464));
  AND2_X1   g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT79), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT25), .ZN(new_n467));
  AOI21_X1  g281(.A(G902), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n466), .A2(new_n467), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n463), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n462), .A2(new_n468), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n473), .B1(new_n474), .B2(new_n470), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n465), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n442), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G221), .B1(new_n295), .B2(G902), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G469), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(new_n274), .ZN(new_n481));
  AOI22_X1  g295(.A1(new_n339), .A2(new_n369), .B1(new_n372), .B2(new_n346), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT10), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT80), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n277), .A3(G104), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT3), .ZN(new_n487));
  INV_X1    g301(.A(G101), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT3), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n485), .A2(new_n489), .A3(new_n277), .A4(G104), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n277), .A2(G104), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n487), .A2(new_n488), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n494));
  INV_X1    g308(.A(G104), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(G107), .ZN(new_n496));
  OAI21_X1  g310(.A(G101), .B1(new_n496), .B2(new_n491), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n493), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n494), .B1(new_n493), .B2(new_n497), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n484), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n367), .A2(new_n344), .A3(new_n369), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n367), .A2(new_n344), .B1(G128), .B2(new_n371), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n493), .A2(new_n497), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n483), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n491), .B1(new_n486), .B2(KEYINPUT3), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n490), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT4), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(G101), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n488), .B1(new_n506), .B2(new_n490), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n509), .B(new_n347), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n361), .A2(new_n365), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n500), .A2(new_n505), .A3(new_n512), .A4(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n500), .A2(new_n505), .A3(new_n512), .ZN(new_n515));
  INV_X1    g329(.A(new_n513), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n515), .A2(KEYINPUT84), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT84), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n308), .A2(G227), .ZN(new_n520));
  XOR2_X1   g334(.A(G110), .B(G140), .Z(new_n521));
  XOR2_X1   g335(.A(new_n520), .B(new_n521), .Z(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n493), .B(new_n497), .C1(new_n501), .C2(new_n502), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n504), .A2(new_n482), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OR2_X1    g341(.A1(KEYINPUT83), .A2(KEYINPUT12), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT82), .B1(new_n525), .B2(new_n526), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n529), .B(new_n516), .C1(KEYINPUT83), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n516), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT12), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n514), .A2(new_n522), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(G902), .B1(new_n524), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n481), .B1(new_n537), .B2(new_n480), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n531), .A2(new_n533), .A3(new_n514), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n523), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n535), .B1(new_n517), .B2(new_n518), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(G469), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n479), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(G214), .B1(G237), .B2(G902), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n374), .A2(G125), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(G125), .B2(new_n396), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n190), .A2(G224), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(KEYINPUT7), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT85), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n546), .A2(new_n550), .B1(KEYINPUT7), .B2(new_n548), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n396), .A2(G125), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n552), .B(KEYINPUT85), .C1(G125), .C2(new_n374), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n278), .A2(G119), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT5), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n324), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n557), .B1(new_n323), .B2(new_n556), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n331), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n504), .ZN(new_n561));
  XNOR2_X1  g375(.A(G110), .B(G122), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n559), .A2(new_n493), .A3(new_n497), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AND3_X1   g379(.A1(new_n549), .A2(new_n554), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n560), .B1(new_n498), .B2(new_n499), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n510), .A2(new_n511), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n509), .A2(new_n390), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n567), .B(new_n562), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(G902), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n562), .ZN(new_n572));
  INV_X1    g386(.A(new_n567), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n569), .A2(new_n568), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(KEYINPUT6), .A3(new_n570), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT6), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n577), .B(new_n572), .C1(new_n573), .C2(new_n574), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n547), .B(new_n548), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n571), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G210), .B1(G237), .B2(G902), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n571), .A2(new_n580), .A3(new_n582), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n545), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n543), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n317), .A2(new_n477), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  NAND2_X1  g403(.A1(new_n472), .A2(new_n475), .ZN(new_n590));
  INV_X1    g404(.A(new_n465), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n436), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n428), .B1(new_n440), .B2(new_n274), .ZN(new_n594));
  NOR4_X1   g408(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n311), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n298), .A2(new_n299), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT33), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G478), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n300), .A2(G478), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n301), .A2(new_n274), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n269), .B2(new_n276), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n587), .A2(new_n595), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT34), .B(G104), .Z(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(G6));
  NAND2_X1  g420(.A1(new_n254), .A2(new_n261), .ZN(new_n607));
  INV_X1    g421(.A(new_n267), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n264), .B(new_n266), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n276), .ZN(new_n610));
  INV_X1    g424(.A(new_n305), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n587), .A3(new_n595), .ZN(new_n613));
  XOR2_X1   g427(.A(KEYINPUT35), .B(G107), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G9));
  INV_X1    g429(.A(KEYINPUT36), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n447), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n617), .B(new_n461), .Z(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n464), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n590), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n621), .A2(new_n594), .A3(new_n593), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n317), .A2(new_n587), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT37), .B(G110), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G12));
  AND4_X1   g439(.A1(new_n442), .A2(new_n586), .A3(new_n543), .A4(new_n620), .ZN(new_n626));
  INV_X1    g440(.A(G900), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n307), .B1(new_n309), .B2(new_n627), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n610), .A2(new_n611), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G128), .ZN(G30));
  NAND2_X1  g445(.A1(new_n524), .A2(new_n536), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n480), .A3(new_n274), .ZN(new_n633));
  INV_X1    g447(.A(new_n481), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(new_n542), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(new_n628), .B(KEYINPUT39), .Z(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n478), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n543), .A2(KEYINPUT40), .A3(new_n636), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT94), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT94), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n639), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n571), .A2(new_n582), .A3(new_n580), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n582), .B1(new_n571), .B2(new_n580), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT93), .B(KEYINPUT38), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n420), .A2(new_n424), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n417), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n653), .B(new_n274), .C1(new_n410), .C2(new_n417), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G472), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n438), .A2(new_n441), .A3(new_n655), .ZN(new_n656));
  AND4_X1   g470(.A1(new_n544), .A2(new_n651), .A3(new_n621), .A4(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n611), .B1(new_n269), .B2(new_n276), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n642), .A2(new_n644), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G143), .ZN(G45));
  INV_X1    g474(.A(KEYINPUT95), .ZN(new_n661));
  INV_X1    g475(.A(new_n628), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n603), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n602), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n262), .A2(new_n265), .A3(KEYINPUT20), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n265), .B1(new_n262), .B2(KEYINPUT20), .ZN(new_n666));
  INV_X1    g480(.A(new_n268), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n665), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n664), .B(new_n662), .C1(new_n668), .C2(new_n275), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT95), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n626), .A2(new_n663), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G146), .ZN(G48));
  AOI22_X1  g486(.A1(new_n519), .A2(new_n523), .B1(new_n534), .B2(new_n535), .ZN(new_n673));
  OAI21_X1  g487(.A(G469), .B1(new_n673), .B2(G902), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n633), .A2(new_n674), .A3(new_n478), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n442), .A2(new_n476), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT96), .ZN(new_n677));
  INV_X1    g491(.A(new_n311), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n678), .B(new_n544), .C1(new_n645), .C2(new_n646), .ZN(new_n679));
  AOI211_X1 g493(.A(new_n602), .B(new_n679), .C1(new_n269), .C2(new_n276), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n676), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n442), .A2(new_n476), .A3(new_n675), .ZN(new_n682));
  INV_X1    g496(.A(new_n679), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n603), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT96), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n681), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT97), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n686), .B(new_n688), .ZN(G15));
  NAND4_X1  g503(.A1(new_n609), .A2(new_n683), .A3(new_n276), .A4(new_n305), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n682), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n278), .ZN(G18));
  AND2_X1   g506(.A1(new_n442), .A2(new_n620), .ZN(new_n693));
  AND4_X1   g507(.A1(new_n586), .A2(new_n478), .A3(new_n633), .A4(new_n674), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n317), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  NAND2_X1  g510(.A1(new_n269), .A2(new_n276), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n697), .A2(new_n305), .A3(new_n586), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n440), .A2(new_n274), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G472), .ZN(new_n700));
  NOR2_X1   g514(.A1(G472), .A2(G902), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n417), .B1(new_n411), .B2(new_n412), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n701), .B1(new_n433), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT98), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT98), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n705), .B(new_n701), .C1(new_n433), .C2(new_n702), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n700), .A2(new_n704), .A3(new_n476), .A4(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n633), .A2(new_n674), .A3(new_n678), .A4(new_n478), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n698), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT99), .B(G122), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G24));
  NAND4_X1  g526(.A1(new_n620), .A2(new_n700), .A3(new_n704), .A4(new_n706), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n670), .A2(new_n663), .A3(new_n694), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  NOR2_X1   g530(.A1(new_n479), .A2(new_n545), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n584), .A2(new_n585), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n515), .A2(new_n516), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT84), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n515), .A2(KEYINPUT84), .A3(new_n516), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n723), .A2(new_n535), .B1(new_n539), .B2(new_n523), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT100), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n725), .A3(G469), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n542), .A2(KEYINPUT100), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n718), .B1(new_n728), .B2(new_n538), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n442), .A2(new_n476), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n670), .A3(new_n663), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n436), .A2(KEYINPUT101), .A3(new_n437), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n427), .A3(new_n441), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT101), .B1(new_n436), .B2(new_n437), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n476), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n633), .A2(new_n634), .A3(new_n727), .A4(new_n726), .ZN(new_n739));
  INV_X1    g553(.A(new_n718), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n738), .A2(new_n663), .A3(new_n670), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n733), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  NAND2_X1  g558(.A1(new_n730), .A2(new_n629), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G134), .ZN(G36));
  NOR2_X1   g560(.A1(new_n697), .A2(new_n602), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT43), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n697), .B2(new_n602), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(KEYINPUT102), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n621), .B1(new_n436), .B2(new_n700), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT102), .B1(new_n748), .B2(new_n750), .ZN(new_n755));
  OR3_X1    g569(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n754), .B1(new_n753), .B2(new_n755), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n724), .A2(KEYINPUT45), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n724), .A2(KEYINPUT45), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(G469), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n758), .B1(new_n762), .B2(new_n481), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n634), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n763), .A2(new_n633), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n478), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n647), .A2(new_n544), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n767), .A2(new_n636), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n756), .A2(new_n757), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  XOR2_X1   g586(.A(new_n766), .B(KEYINPUT47), .Z(new_n773));
  AND2_X1   g587(.A1(new_n670), .A2(new_n663), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n442), .A2(new_n476), .A3(new_n768), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G140), .ZN(G42));
  INV_X1    g592(.A(new_n307), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n779), .B(new_n707), .C1(new_n748), .C2(new_n750), .ZN(new_n780));
  INV_X1    g594(.A(new_n675), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n651), .A2(new_n781), .A3(new_n544), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT50), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n780), .A2(KEYINPUT50), .A3(new_n782), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n781), .A2(new_n768), .ZN(new_n788));
  INV_X1    g602(.A(new_n656), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n592), .A2(new_n779), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n792), .A2(new_n269), .A3(new_n276), .A4(new_n602), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n748), .A2(new_n750), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n307), .A3(new_n788), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n793), .B1(new_n795), .B2(new_n713), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n787), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT107), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT107), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n787), .B2(new_n796), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n766), .B(KEYINPUT47), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n633), .A2(new_n674), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(KEYINPUT106), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(KEYINPUT106), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n479), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n780), .A2(new_n769), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n801), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n798), .A2(new_n800), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT108), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n798), .A2(KEYINPUT108), .A3(new_n800), .A4(new_n809), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n795), .A2(new_n737), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n814), .A2(KEYINPUT109), .A3(KEYINPUT48), .ZN(new_n815));
  INV_X1    g629(.A(new_n603), .ZN(new_n816));
  OAI211_X1 g630(.A(G952), .B(new_n190), .C1(new_n791), .C2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n817), .B1(new_n694), .B2(new_n780), .ZN(new_n818));
  XNOR2_X1  g632(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n815), .B(new_n818), .C1(new_n814), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n807), .A2(new_n808), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n797), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n820), .B1(new_n822), .B2(new_n801), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n812), .A2(new_n813), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT105), .ZN(new_n825));
  INV_X1    g639(.A(new_n709), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n658), .A2(new_n586), .ZN(new_n827));
  OAI22_X1  g641(.A1(new_n826), .A2(new_n827), .B1(new_n682), .B2(new_n690), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n694), .A2(new_n442), .A3(new_n620), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n316), .B2(new_n314), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n303), .A2(new_n304), .A3(new_n662), .ZN(new_n832));
  NOR4_X1   g646(.A1(new_n645), .A2(new_n646), .A3(new_n832), .A4(new_n545), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n635), .A3(new_n478), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n610), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n730), .A2(new_n629), .B1(new_n693), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n743), .A2(new_n686), .A3(new_n831), .A4(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n697), .A2(new_n611), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n587), .B(new_n595), .C1(new_n838), .C2(new_n603), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n588), .A2(new_n623), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n739), .A2(new_n740), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n713), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n670), .A2(new_n842), .A3(new_n663), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT104), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT104), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n670), .A2(new_n663), .A3(new_n842), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n825), .B1(new_n837), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n588), .A2(new_n623), .A3(new_n839), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n844), .B2(new_n846), .ZN(new_n851));
  INV_X1    g665(.A(new_n690), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n676), .A2(new_n852), .B1(new_n698), .B2(new_n709), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n686), .A2(new_n695), .A3(new_n853), .A4(new_n836), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n851), .A2(new_n854), .A3(KEYINPUT105), .A4(new_n743), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n739), .A2(new_n478), .A3(new_n662), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n698), .A2(new_n621), .A3(new_n656), .A4(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n671), .A2(new_n715), .A3(new_n630), .A4(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT52), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT53), .B1(new_n856), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n715), .A2(new_n630), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT53), .B1(new_n863), .B2(KEYINPUT52), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n864), .B(new_n860), .C1(new_n849), .C2(new_n855), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT54), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n837), .A2(new_n848), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n869), .B1(new_n863), .B2(KEYINPUT52), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n861), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n860), .B1(new_n849), .B2(new_n855), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n867), .B(new_n871), .C1(new_n872), .C2(KEYINPUT53), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  OAI22_X1  g688(.A1(new_n824), .A2(new_n874), .B1(G952), .B2(G953), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n476), .A2(new_n717), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT103), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n651), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n803), .B(KEYINPUT49), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n789), .A3(new_n747), .A4(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n875), .A2(new_n880), .ZN(G75));
  NOR2_X1   g695(.A1(new_n308), .A2(G952), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n871), .B1(new_n872), .B2(KEYINPUT53), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(G210), .A2(G902), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n576), .A2(new_n578), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(new_n579), .ZN(new_n889));
  XNOR2_X1  g703(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n889), .B(new_n890), .Z(new_n891));
  XOR2_X1   g705(.A(KEYINPUT112), .B(KEYINPUT56), .Z(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n883), .B1(new_n887), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n886), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT56), .B1(new_n884), .B2(new_n895), .ZN(new_n896));
  OR3_X1    g710(.A1(new_n896), .A2(KEYINPUT111), .A3(new_n891), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT111), .B1(new_n896), .B2(new_n891), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(G51));
  XNOR2_X1  g713(.A(KEYINPUT113), .B(KEYINPUT57), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n481), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n686), .A2(new_n695), .A3(new_n853), .A4(new_n836), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n741), .B(new_n476), .C1(new_n735), .C2(new_n736), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  AOI22_X1  g718(.A1(new_n774), .A2(new_n904), .B1(new_n731), .B2(new_n732), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT105), .B1(new_n906), .B2(new_n851), .ZN(new_n907));
  NOR4_X1   g721(.A1(new_n848), .A2(new_n902), .A3(new_n825), .A4(new_n905), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n861), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n869), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n867), .B1(new_n910), .B2(new_n871), .ZN(new_n911));
  INV_X1    g725(.A(new_n873), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n901), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n632), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n884), .A2(G902), .A3(new_n762), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n882), .B1(new_n914), .B2(new_n915), .ZN(G54));
  INV_X1    g730(.A(KEYINPUT58), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n270), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n884), .A2(G902), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(new_n607), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n607), .A2(new_n917), .A3(new_n270), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n884), .A2(G902), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n883), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT114), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(new_n607), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT114), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n925), .A2(new_n926), .A3(new_n883), .A4(new_n922), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(new_n927), .ZN(G60));
  XOR2_X1   g742(.A(new_n597), .B(KEYINPUT115), .Z(new_n929));
  XOR2_X1   g743(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n600), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n929), .B(new_n931), .C1(new_n911), .C2(new_n912), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n883), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n874), .B2(new_n931), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(G63));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT60), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n884), .A2(new_n618), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n937), .B1(new_n910), .B2(new_n871), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n883), .B(new_n939), .C1(new_n940), .C2(new_n462), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n447), .A2(new_n461), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n447), .A2(new_n461), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n944), .B(new_n945), .C1(new_n885), .C2(new_n937), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n946), .A2(KEYINPUT61), .A3(new_n883), .A4(new_n939), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n947), .ZN(G66));
  INV_X1    g762(.A(G224), .ZN(new_n949));
  OAI21_X1  g763(.A(G953), .B1(new_n310), .B2(new_n949), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT117), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n840), .A2(new_n686), .A3(new_n831), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n308), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n888), .B1(G898), .B2(new_n308), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  NAND2_X1  g771(.A1(new_n743), .A2(new_n745), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT121), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n767), .A2(new_n636), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n737), .A2(new_n827), .ZN(new_n961));
  AOI22_X1  g775(.A1(new_n773), .A2(new_n776), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n671), .A2(new_n715), .A3(new_n630), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n959), .A2(new_n962), .A3(new_n771), .A4(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n965), .A2(new_n954), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n421), .A2(new_n423), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n248), .A2(new_n237), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(new_n627), .B2(new_n308), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n308), .B1(G227), .B2(G900), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT120), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  INV_X1    g789(.A(new_n659), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n975), .B1(new_n976), .B2(new_n963), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n964), .A2(KEYINPUT62), .A3(new_n659), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n838), .A2(new_n603), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n442), .A2(new_n476), .ZN(new_n981));
  NOR4_X1   g795(.A1(new_n980), .A2(new_n981), .A3(new_n637), .A4(new_n768), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n773), .B2(new_n776), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n979), .A2(new_n983), .A3(new_n771), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(KEYINPUT118), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT118), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n979), .A2(new_n983), .A3(new_n771), .A4(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n954), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n988), .A2(new_n969), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(KEYINPUT119), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT119), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(new_n988), .B2(new_n969), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n974), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n972), .B1(new_n989), .B2(new_n971), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(G72));
  NAND3_X1  g809(.A1(new_n985), .A2(new_n953), .A3(new_n987), .ZN(new_n996));
  XOR2_X1   g810(.A(KEYINPUT122), .B(KEYINPUT63), .Z(new_n997));
  NOR2_X1   g811(.A1(new_n428), .A2(new_n274), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT123), .Z(new_n1000));
  NAND2_X1  g814(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n653), .ZN(new_n1002));
  AOI21_X1  g816(.A(KEYINPUT124), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT124), .ZN(new_n1004));
  AOI211_X1 g818(.A(new_n1004), .B(new_n653), .C1(new_n996), .C2(new_n1000), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1000), .B1(new_n965), .B2(new_n952), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n425), .B(KEYINPUT125), .Z(new_n1008));
  AOI21_X1  g822(.A(new_n882), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n864), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n872), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n910), .A2(new_n1011), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n653), .A2(new_n425), .A3(new_n999), .ZN(new_n1013));
  AOI21_X1  g827(.A(KEYINPUT126), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g828(.A(KEYINPUT126), .B(new_n1013), .C1(new_n862), .C2(new_n865), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1009), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1006), .A2(new_n1017), .ZN(G57));
endmodule


