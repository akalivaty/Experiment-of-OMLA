//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n549, new_n550, new_n551, new_n552, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n562, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g033(.A(G261), .ZN(G325));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  OR2_X1    g035(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(G567), .ZN(new_n463));
  OR3_X1    g038(.A1(new_n456), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n462), .B1(new_n456), .B2(new_n463), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n461), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(KEYINPUT68), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2104), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n477), .A2(new_n479), .A3(KEYINPUT3), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  NAND4_X1  g056(.A1(new_n480), .A2(G137), .A3(new_n481), .A4(new_n470), .ZN(new_n482));
  XNOR2_X1  g057(.A(KEYINPUT68), .B(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G101), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n476), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G160));
  NAND2_X1  g062(.A1(new_n480), .A2(new_n470), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(new_n481), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n481), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n488), .A2(G2105), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(G136), .B2(new_n494), .ZN(G162));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n470), .A2(new_n472), .A3(new_n481), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT4), .A2(G138), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n480), .A2(new_n481), .A3(new_n470), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n480), .A2(new_n470), .A3(new_n503), .ZN(new_n504));
  OR2_X1    g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(G2104), .C1(G114), .C2(new_n481), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n504), .A2(KEYINPUT69), .A3(new_n506), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n502), .B1(new_n509), .B2(new_n510), .ZN(G164));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n516), .A2(KEYINPUT73), .B1(G75), .B2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n512), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G50), .ZN(new_n520));
  AOI21_X1  g095(.A(KEYINPUT70), .B1(KEYINPUT71), .B2(G651), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT6), .B1(new_n523), .B2(new_n512), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n521), .A2(KEYINPUT6), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n525), .A2(G543), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n525), .A2(new_n515), .A3(new_n526), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT72), .B(G88), .Z(new_n529));
  OAI22_X1  g104(.A1(new_n520), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n519), .A2(new_n530), .ZN(G166));
  XNOR2_X1  g106(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n532));
  AND3_X1   g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n515), .A2(new_n535), .A3(G63), .A4(G651), .ZN(new_n536));
  INV_X1    g111(.A(new_n515), .ZN(new_n537));
  NAND2_X1  g112(.A1(G63), .A2(G651), .ZN(new_n538));
  OAI21_X1  g113(.A(KEYINPUT74), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n534), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n528), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G89), .ZN(new_n542));
  INV_X1    g117(.A(new_n527), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G51), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n540), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(KEYINPUT76), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(KEYINPUT76), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(G168));
  NAND2_X1  g123(.A1(new_n543), .A2(G52), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n541), .A2(G90), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(new_n512), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(new_n550), .A3(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  NAND2_X1  g129(.A1(new_n543), .A2(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n541), .A2(G81), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n512), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  INV_X1    g141(.A(KEYINPUT6), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(KEYINPUT70), .B2(G651), .ZN(new_n568));
  MUX2_X1   g143(.A(new_n568), .B(new_n567), .S(new_n521), .Z(new_n569));
  NAND3_X1  g144(.A1(new_n569), .A2(G91), .A3(new_n515), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT79), .ZN(new_n571));
  XOR2_X1   g146(.A(KEYINPUT78), .B(KEYINPUT9), .Z(new_n572));
  NAND3_X1  g147(.A1(new_n543), .A2(G53), .A3(new_n572), .ZN(new_n573));
  NOR2_X1   g148(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n527), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n573), .B(new_n576), .C1(new_n512), .C2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n571), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G299));
  INV_X1    g155(.A(G168), .ZN(G286));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND4_X1  g157(.A1(new_n525), .A2(G49), .A3(G543), .A4(new_n526), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT80), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n569), .A2(new_n586), .A3(G87), .A4(new_n515), .ZN(new_n587));
  INV_X1    g162(.A(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT80), .B1(new_n528), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n585), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G288));
  NAND4_X1  g166(.A1(new_n525), .A2(G48), .A3(G543), .A4(new_n526), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n525), .A2(G86), .A3(new_n515), .A4(new_n526), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n513), .B2(new_n514), .ZN(new_n595));
  AND2_X1   g170(.A1(G73), .A2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n592), .A2(new_n593), .A3(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n543), .A2(G47), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n541), .A2(G85), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n601), .A2(new_n512), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT81), .B1(new_n528), .B2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  NOR3_X1   g184(.A1(new_n528), .A2(KEYINPUT81), .A3(new_n607), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n606), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n610), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n608), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n537), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n543), .A2(G54), .B1(new_n616), .B2(G651), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n611), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n605), .B1(new_n619), .B2(G868), .ZN(G284));
  XOR2_X1   g195(.A(G284), .B(KEYINPUT82), .Z(G321));
  NOR2_X1   g196(.A1(G299), .A2(G868), .ZN(new_n622));
  AOI21_X1  g197(.A(new_n622), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g198(.A(new_n622), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n619), .B1(new_n625), .B2(G860), .ZN(G148));
  NOR2_X1   g201(.A1(new_n560), .A2(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n625), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT83), .Z(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g206(.A1(new_n497), .A2(new_n483), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n494), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n489), .A2(G123), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT84), .ZN(new_n639));
  INV_X1    g214(.A(G111), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n638), .A2(new_n639), .B1(new_n640), .B2(G2105), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n639), .B2(new_n638), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n636), .A2(new_n637), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n635), .A2(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT85), .B(G2438), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(KEYINPUT14), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT86), .Z(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT16), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n655), .B(new_n656), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n653), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n661), .A3(G14), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G401));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT87), .Z(new_n666));
  NOR2_X1   g241(.A1(G2072), .A2(G2078), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n444), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n664), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(KEYINPUT17), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n669), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n664), .B(new_n665), .C1(new_n444), .C2(new_n667), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT18), .Z(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n666), .A3(new_n664), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2100), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT88), .B(G2096), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(G227));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1961), .B(G1966), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n681), .A2(new_n682), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n683), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT20), .Z(new_n687));
  AOI211_X1 g262(.A(new_n685), .B(new_n687), .C1(new_n680), .C2(new_n684), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G4), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(new_n619), .B2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G1348), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G32), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n494), .A2(G141), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n489), .A2(G129), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT26), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n484), .A2(G105), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n702), .A2(new_n703), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n701), .B1(new_n714), .B2(new_n700), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT27), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G1996), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n699), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G29), .A2(G35), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G162), .B2(G29), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G2090), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT90), .B(G16), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n727), .A2(G19), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n560), .B2(new_n727), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT93), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(G1341), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(G1341), .ZN(new_n732));
  NOR3_X1   g307(.A1(new_n725), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g308(.A1(G168), .A2(new_n695), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n695), .B2(G21), .ZN(new_n735));
  INV_X1    g310(.A(G1966), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT30), .B(G28), .ZN(new_n738));
  OR2_X1    g313(.A1(KEYINPUT31), .A2(G11), .ZN(new_n739));
  NAND2_X1  g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n738), .A2(new_n700), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G34), .ZN(new_n742));
  AOI21_X1  g317(.A(G29), .B1(new_n742), .B2(KEYINPUT24), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(KEYINPUT24), .B2(new_n742), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n486), .B2(new_n700), .ZN(new_n745));
  INV_X1    g320(.A(G2084), .ZN(new_n746));
  OAI221_X1 g321(.A(new_n741), .B1(new_n643), .B2(new_n700), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n695), .A2(G5), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G171), .B2(new_n695), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G1961), .ZN(new_n750));
  AOI211_X1 g325(.A(new_n747), .B(new_n750), .C1(new_n746), .C2(new_n745), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n735), .A2(new_n736), .B1(new_n724), .B2(new_n723), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n733), .A2(new_n737), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n716), .A2(G1996), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n700), .A2(G26), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT28), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n494), .A2(G140), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n489), .A2(G128), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G116), .C2(new_n481), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n756), .B1(new_n761), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2067), .ZN(new_n763));
  NOR2_X1   g338(.A1(G29), .A2(G33), .ZN(new_n764));
  XOR2_X1   g339(.A(new_n764), .B(KEYINPUT94), .Z(new_n765));
  NAND2_X1  g340(.A1(new_n494), .A2(G139), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT95), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(G115), .A2(G2104), .ZN(new_n769));
  INV_X1    g344(.A(G127), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n473), .B2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT25), .ZN(new_n772));
  NAND2_X1  g347(.A1(G103), .A2(G2104), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(G2105), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n481), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n771), .A2(G2105), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n768), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n765), .B1(new_n777), .B2(new_n700), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n763), .B1(new_n778), .B2(new_n442), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n442), .B2(new_n778), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n726), .A2(G20), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT23), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n579), .B2(new_n695), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1956), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n700), .A2(G27), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G164), .B2(new_n700), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT97), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(new_n443), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n780), .A2(new_n784), .A3(new_n788), .ZN(new_n789));
  NOR4_X1   g364(.A1(new_n719), .A2(new_n753), .A3(new_n754), .A4(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G6), .B(G305), .S(G16), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT91), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT32), .B(G1981), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n590), .A2(new_n695), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n695), .B2(G23), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT33), .B(G1976), .Z(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n727), .A2(G22), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G166), .B2(new_n727), .ZN(new_n801));
  INV_X1    g376(.A(G1971), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n796), .A2(new_n798), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n799), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  OR3_X1    g380(.A1(new_n794), .A2(new_n805), .A3(KEYINPUT34), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT34), .B1(new_n794), .B2(new_n805), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n727), .A2(G24), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n603), .B2(new_n727), .ZN(new_n809));
  INV_X1    g384(.A(G1986), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(G25), .A2(G29), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n494), .A2(G131), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n489), .A2(G119), .ZN(new_n814));
  OR2_X1    g389(.A1(G95), .A2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n815), .B(G2104), .C1(G107), .C2(new_n481), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n812), .B1(new_n818), .B2(G29), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT35), .B(G1991), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT89), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n811), .A2(new_n822), .A3(KEYINPUT92), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n806), .A2(new_n807), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n790), .A2(new_n825), .A3(new_n826), .ZN(G150));
  INV_X1    g402(.A(G150), .ZN(G311));
  NAND2_X1  g403(.A1(new_n619), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n543), .A2(G55), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n541), .A2(G93), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n831), .B(new_n832), .C1(new_n512), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n560), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n830), .B(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n837), .A2(new_n838), .A3(G860), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n834), .A2(G860), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT37), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n839), .A2(new_n841), .ZN(G145));
  NAND2_X1  g417(.A1(new_n489), .A2(G130), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT99), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n494), .A2(G142), .ZN(new_n845));
  OR2_X1    g420(.A1(G106), .A2(G2105), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(G2104), .C1(G118), .C2(new_n481), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n761), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n711), .A2(new_n712), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n850), .B1(new_n711), .B2(new_n712), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  INV_X1    g430(.A(new_n849), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n855), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n817), .B(new_n633), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n858), .B1(new_n854), .B2(new_n857), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n502), .A2(new_n507), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n854), .A2(new_n857), .ZN(new_n865));
  INV_X1    g440(.A(new_n858), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n864), .B1(new_n867), .B2(new_n859), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n777), .B1(new_n863), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n862), .B1(new_n860), .B2(new_n861), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n864), .A3(new_n859), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n870), .A2(new_n768), .A3(new_n776), .A4(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n643), .B(new_n486), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(G162), .Z(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G37), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n874), .B1(new_n869), .B2(new_n872), .ZN(new_n878));
  OAI21_X1  g453(.A(KEYINPUT100), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n880), .A2(new_n881), .A3(new_n875), .A4(new_n876), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g459(.A1(new_n579), .A2(new_n618), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT101), .ZN(new_n886));
  NAND2_X1  g461(.A1(G299), .A2(new_n619), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n579), .A2(new_n618), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT102), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n890), .A2(new_n894), .A3(new_n891), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n891), .B1(G299), .B2(new_n619), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(new_n885), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n835), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n628), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n887), .A2(new_n885), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n902), .B(new_n904), .C1(new_n905), .C2(KEYINPUT42), .ZN(new_n906));
  XOR2_X1   g481(.A(G166), .B(G305), .Z(new_n907));
  XNOR2_X1  g482(.A(new_n603), .B(new_n590), .ZN(new_n908));
  XOR2_X1   g483(.A(new_n907), .B(new_n908), .Z(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n910), .B1(new_n905), .B2(KEYINPUT42), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n905), .A2(KEYINPUT42), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n892), .A2(KEYINPUT102), .B1(new_n885), .B2(new_n896), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n900), .B1(new_n913), .B2(new_n895), .ZN(new_n914));
  INV_X1    g489(.A(new_n904), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n906), .A2(new_n911), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n911), .B1(new_n906), .B2(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G868), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n834), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(G295));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n919), .A2(new_n923), .A3(new_n921), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n923), .B1(new_n919), .B2(new_n921), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(G331));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  XNOR2_X1  g502(.A(G301), .B(KEYINPUT105), .ZN(new_n928));
  OR2_X1    g503(.A1(G168), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G168), .A2(new_n928), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n835), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n932), .A2(new_n903), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n899), .A3(new_n930), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n929), .A2(KEYINPUT107), .A3(new_n899), .A4(new_n930), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n933), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n932), .A2(new_n934), .ZN(new_n939));
  AND3_X1   g514(.A1(new_n898), .A2(KEYINPUT106), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT106), .B1(new_n898), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G37), .B1(new_n942), .B2(new_n909), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  OAI211_X1 g519(.A(new_n910), .B(new_n938), .C1(new_n940), .C2(new_n941), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n936), .A2(new_n932), .A3(new_n937), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT108), .B1(new_n903), .B2(new_n891), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n903), .A2(KEYINPUT108), .A3(new_n891), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n896), .A2(new_n886), .A3(new_n889), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n947), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n933), .A2(new_n934), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G37), .B1(new_n954), .B2(new_n909), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n945), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n927), .B1(new_n946), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n944), .B1(new_n943), .B2(new_n945), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n955), .A2(new_n945), .A3(new_n944), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n958), .B1(new_n961), .B2(new_n927), .ZN(G397));
  INV_X1    g537(.A(KEYINPUT123), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n476), .A2(G40), .A3(new_n485), .A4(new_n482), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n502), .B2(new_n507), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n499), .A2(new_n501), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n504), .A2(KEYINPUT69), .A3(new_n506), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT69), .B1(new_n504), .B2(new_n506), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(new_n965), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n968), .B1(new_n973), .B2(new_n967), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n736), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n976), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n977));
  INV_X1    g552(.A(new_n964), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(new_n972), .B2(new_n965), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n979), .B(new_n965), .C1(new_n502), .C2(new_n507), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n976), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n977), .B(new_n978), .C1(new_n980), .C2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n975), .B1(new_n984), .B2(G2084), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT122), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(new_n986), .A3(G8), .ZN(new_n987));
  AOI21_X1  g562(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G8), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n509), .A2(new_n510), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n991), .B2(new_n969), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n982), .B1(new_n992), .B2(new_n979), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n993), .A2(new_n746), .A3(new_n978), .A4(new_n977), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n990), .B1(new_n994), .B2(new_n975), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(new_n986), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n963), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n985), .A2(G8), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT122), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n999), .A2(KEYINPUT123), .A3(new_n987), .A4(new_n988), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT51), .B(G8), .C1(new_n985), .C2(G286), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT62), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n985), .A2(G8), .A3(G286), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n590), .B2(G1976), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(KEYINPUT115), .B(new_n1006), .C1(new_n590), .C2(G1976), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n966), .A2(new_n964), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(new_n990), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n590), .A2(G1976), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1011), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1015), .A2(new_n1013), .A3(G8), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT52), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G305), .A2(G1981), .ZN(new_n1018));
  INV_X1    g593(.A(G1981), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n592), .A2(new_n593), .A3(new_n1019), .A4(new_n597), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1018), .A2(KEYINPUT49), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT49), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n1012), .ZN(new_n1024));
  AND4_X1   g599(.A1(KEYINPUT117), .A2(new_n1014), .A3(new_n1017), .A4(new_n1024), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1023), .A2(new_n1012), .B1(new_n1016), .B2(KEYINPUT52), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT117), .B1(new_n1026), .B2(new_n1014), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n978), .B1(new_n966), .B2(new_n967), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT112), .B1(new_n973), .B2(new_n967), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n1032));
  AOI211_X1 g607(.A(new_n1032), .B(KEYINPUT45), .C1(new_n972), .C2(new_n965), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1030), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1032), .B1(new_n992), .B2(KEYINPUT45), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n973), .A2(KEYINPUT112), .A3(new_n967), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(KEYINPUT113), .A3(new_n1030), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1040), .A3(new_n802), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n984), .A2(G2090), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n990), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G303), .A2(G8), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT55), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1028), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n964), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n973), .B2(KEYINPUT50), .ZN(new_n1049));
  OR2_X1    g624(.A1(new_n1049), .A2(G2090), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1041), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(G8), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n1045), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT113), .B1(new_n1039), .B2(new_n1030), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n1035), .B(new_n1029), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n443), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OR3_X1    g633(.A1(new_n974), .A2(new_n1057), .A3(G2078), .ZN(new_n1059));
  INV_X1    g634(.A(G1961), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n984), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(G301), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1047), .A2(new_n1053), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1005), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT125), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT125), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1005), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT126), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1067), .A2(new_n1069), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1046), .B1(new_n1051), .B2(G8), .ZN(new_n1076));
  AOI211_X1 g651(.A(new_n990), .B(new_n1045), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1077));
  NOR3_X1   g652(.A1(new_n1076), .A2(new_n1077), .A3(new_n1028), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n966), .A2(KEYINPUT109), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT45), .B1(new_n966), .B2(KEYINPUT109), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(KEYINPUT53), .A3(new_n1030), .A4(new_n443), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1061), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(G2078), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1085));
  OAI211_X1 g660(.A(G301), .B(new_n1084), .C1(new_n1085), .C2(KEYINPUT53), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1062), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(G301), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1058), .A2(G301), .A3(new_n1063), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1083), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1091), .B(KEYINPUT54), .C1(new_n1092), .C2(G301), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1070), .A2(new_n1078), .A3(new_n1090), .A4(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1063), .B1(new_n1085), .B2(KEYINPUT53), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G171), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT54), .B1(new_n1098), .B2(new_n1086), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1047), .A2(new_n1053), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1101), .A2(KEYINPUT124), .A3(new_n1070), .A4(new_n1093), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT58), .B(G1341), .ZN(new_n1103));
  OAI22_X1  g678(.A1(new_n1034), .A2(G1996), .B1(new_n1011), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n560), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n1108));
  INV_X1    g683(.A(G2067), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n984), .A2(new_n698), .B1(new_n1109), .B2(new_n1011), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1110), .A2(new_n618), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n618), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1108), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1110), .A2(new_n1108), .A3(new_n619), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1107), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT56), .B(G2072), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1039), .A2(new_n1030), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g696(.A(KEYINPUT119), .B(G1956), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1049), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1126));
  XOR2_X1   g701(.A(new_n579), .B(new_n1126), .Z(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1127), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1121), .A2(new_n1129), .A3(new_n1124), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(KEYINPUT61), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1129), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n1123), .B(new_n1127), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1115), .A2(new_n1131), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1111), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1133), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1096), .A2(new_n1102), .A3(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G288), .A2(G1976), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT116), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1020), .B1(new_n1142), .B2(new_n1023), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1012), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1077), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1026), .A2(new_n1014), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1144), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n995), .A2(G168), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT118), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1078), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1077), .A2(new_n1151), .A3(new_n1146), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1153), .B(new_n1149), .C1(new_n1046), .C2(new_n1043), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1147), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1075), .A2(new_n1140), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1081), .A2(new_n964), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n603), .A2(new_n810), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT110), .Z(new_n1160));
  NAND2_X1  g735(.A1(G290), .A2(G1986), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1158), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT111), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n761), .B(new_n1109), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n714), .A2(G1996), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n713), .A2(new_n718), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n817), .B(new_n821), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1158), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1163), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1156), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1157), .A2(new_n718), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT46), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n714), .A2(new_n1164), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1174), .B1(new_n1158), .B2(new_n1175), .ZN(new_n1176));
  XOR2_X1   g751(.A(new_n1176), .B(KEYINPUT47), .Z(new_n1177));
  NOR2_X1   g752(.A1(new_n1160), .A2(new_n1158), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT127), .Z(new_n1179));
  INV_X1    g754(.A(KEYINPUT48), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1181), .A2(new_n1182), .A3(new_n1170), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n818), .A2(new_n821), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1167), .A2(new_n1184), .B1(G2067), .B2(new_n761), .ZN(new_n1185));
  AOI211_X1 g760(.A(new_n1177), .B(new_n1183), .C1(new_n1157), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1172), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g762(.A1(G229), .A2(new_n466), .A3(G401), .A4(G227), .ZN(new_n1189));
  OAI211_X1 g763(.A(new_n883), .B(new_n1189), .C1(new_n959), .C2(new_n960), .ZN(G225));
  INV_X1    g764(.A(G225), .ZN(G308));
endmodule


