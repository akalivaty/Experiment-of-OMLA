//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  OR2_X1    g000(.A1(KEYINPUT64), .A2(G143), .ZN(new_n187));
  NAND2_X1  g001(.A1(KEYINPUT64), .A2(G143), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(G146), .A3(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT65), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT65), .A2(G146), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(G143), .A3(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n189), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT69), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT69), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n189), .A2(new_n194), .A3(new_n199), .A4(new_n196), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(G146), .B1(new_n187), .B2(new_n188), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n203));
  OAI21_X1  g017(.A(G128), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n189), .A2(new_n194), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n208), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OR2_X1    g028(.A1(new_n214), .A2(G101), .ZN(new_n215));
  INV_X1    g029(.A(new_n213), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n208), .A2(G107), .ZN(new_n217));
  OAI21_X1  g031(.A(G101), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n207), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n214), .A2(G101), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n215), .A2(new_n223), .A3(KEYINPUT4), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n214), .A2(new_n225), .A3(G101), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT0), .B(G128), .Z(new_n228));
  AOI21_X1  g042(.A(G143), .B1(new_n192), .B2(new_n193), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n202), .B2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n189), .A2(new_n194), .A3(KEYINPUT0), .A4(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n221), .A2(new_n222), .B1(new_n227), .B2(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n202), .A2(new_n229), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G128), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n201), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT10), .A4(new_n220), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n198), .A2(new_n200), .B1(new_n235), .B2(new_n237), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n215), .A2(KEYINPUT10), .A3(new_n218), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT82), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G137), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(G134), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT11), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n248), .A2(KEYINPUT66), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(G134), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G134), .ZN(new_n252));
  OAI22_X1  g066(.A1(KEYINPUT66), .A2(new_n248), .B1(new_n252), .B2(G137), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n248), .A2(KEYINPUT66), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n251), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G131), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n251), .A2(new_n255), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n234), .A2(new_n245), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT83), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT83), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n234), .A2(new_n245), .A3(new_n264), .A4(new_n261), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n233), .A2(new_n224), .A3(new_n226), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n219), .B1(new_n201), .B2(new_n206), .ZN(new_n268));
  INV_X1    g082(.A(new_n222), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n270), .B1(new_n244), .B2(new_n241), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(new_n261), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  INV_X1    g089(.A(G227), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G953), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n275), .B(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n239), .A2(new_n220), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n260), .B1(new_n280), .B2(new_n268), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT12), .ZN(new_n282));
  OR2_X1    g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n281), .A2(new_n282), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n266), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT84), .ZN(new_n287));
  AOI22_X1  g101(.A1(new_n263), .A2(new_n265), .B1(new_n283), .B2(new_n284), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT84), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n279), .B1(new_n291), .B2(new_n278), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G469), .ZN(new_n293));
  INV_X1    g107(.A(G469), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT85), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n274), .A2(new_n278), .ZN(new_n297));
  INV_X1    g111(.A(new_n278), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n266), .A2(new_n298), .A3(new_n285), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n296), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT85), .B1(new_n288), .B2(new_n298), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n294), .B(new_n295), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n294), .A2(new_n295), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n293), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G221), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT9), .B(G234), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n306), .B1(new_n308), .B2(new_n295), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT70), .B(G237), .ZN(new_n311));
  INV_X1    g125(.A(G953), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(G214), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G143), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n187), .A2(new_n188), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n313), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n258), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT17), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n315), .A2(new_n258), .A3(new_n317), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT93), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n319), .A2(KEYINPUT93), .A3(new_n320), .A4(new_n321), .ZN(new_n325));
  XNOR2_X1  g139(.A(G125), .B(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT16), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  OR3_X1    g142(.A1(new_n328), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n191), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n327), .A2(G146), .A3(new_n329), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g147(.A(new_n333), .B(KEYINPUT92), .Z(new_n334));
  NAND2_X1  g148(.A1(new_n318), .A2(KEYINPUT17), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n324), .A2(new_n325), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(KEYINPUT18), .A2(G131), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(KEYINPUT90), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n315), .A2(new_n317), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT91), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n193), .ZN(new_n342));
  NOR2_X1   g156(.A1(KEYINPUT65), .A2(G146), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n344), .A2(new_n326), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  OR2_X1    g160(.A1(new_n326), .A2(new_n191), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n318), .A2(KEYINPUT18), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n336), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G113), .B(G122), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n351), .B(new_n208), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT95), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n336), .A2(new_n352), .A3(new_n349), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n352), .B1(new_n336), .B2(new_n349), .ZN(new_n358));
  AOI21_X1  g172(.A(G902), .B1(new_n358), .B2(KEYINPUT95), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G475), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n314), .A2(G128), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n362), .B1(new_n316), .B2(G128), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n363), .A2(new_n252), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n252), .ZN(new_n365));
  INV_X1    g179(.A(G116), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(G122), .ZN(new_n367));
  INV_X1    g181(.A(G122), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G116), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n364), .A2(new_n365), .B1(new_n211), .B2(new_n370), .ZN(new_n371));
  OR3_X1    g185(.A1(new_n368), .A2(KEYINPUT14), .A3(G116), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT14), .B1(new_n368), .B2(G116), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n372), .B(new_n373), .C1(new_n366), .C2(G122), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G107), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(KEYINPUT97), .ZN(new_n376));
  XOR2_X1   g190(.A(KEYINPUT96), .B(KEYINPUT13), .Z(new_n377));
  NAND3_X1  g191(.A1(new_n363), .A2(KEYINPUT13), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n316), .A2(G128), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n378), .B(G134), .C1(new_n379), .C2(new_n377), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n370), .A2(new_n211), .ZN(new_n381));
  OAI21_X1  g195(.A(G107), .B1(new_n367), .B2(new_n369), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n363), .A2(new_n252), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n371), .A2(new_n376), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G217), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n307), .A2(new_n385), .A3(G953), .ZN(new_n386));
  OR3_X1    g200(.A1(new_n384), .A2(KEYINPUT98), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT98), .B1(new_n384), .B2(new_n386), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(new_n386), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n295), .ZN(new_n391));
  INV_X1    g205(.A(G478), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(KEYINPUT15), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n393), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n390), .B2(new_n295), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n319), .A2(new_n321), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n326), .B(KEYINPUT19), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n344), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n332), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n349), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n353), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n356), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(G475), .A2(G902), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT94), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT20), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n409));
  AOI211_X1 g223(.A(new_n409), .B(new_n406), .C1(new_n356), .C2(new_n403), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(G234), .A2(G237), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n412), .A2(G902), .A3(G953), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT21), .B(G898), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n412), .A2(G952), .A3(new_n312), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n361), .A2(new_n397), .A3(new_n411), .A4(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G210), .B1(G237), .B2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G110), .B(G122), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT8), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n366), .A2(KEYINPUT5), .A3(G119), .ZN(new_n424));
  INV_X1    g238(.A(G113), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G116), .B(G119), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT5), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT2), .B(G113), .Z(new_n429));
  AOI22_X1  g243(.A1(new_n426), .A2(new_n428), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n220), .A2(KEYINPUT87), .A3(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n220), .B2(new_n430), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT87), .B1(new_n220), .B2(new_n430), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n423), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n242), .A2(new_n328), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n312), .A2(G224), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n436), .B(KEYINPUT86), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n232), .A2(G125), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT7), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n220), .A2(new_n430), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n429), .B(new_n427), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n224), .A2(new_n442), .A3(new_n226), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n441), .A2(new_n443), .A3(new_n422), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n435), .A2(new_n438), .ZN(new_n445));
  OR2_X1    g259(.A1(KEYINPUT88), .A2(KEYINPUT7), .ZN(new_n446));
  NAND2_X1  g260(.A1(KEYINPUT88), .A2(KEYINPUT7), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n437), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n434), .A2(new_n440), .A3(new_n444), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n295), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n441), .A2(new_n443), .ZN(new_n452));
  INV_X1    g266(.A(new_n422), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT6), .A3(new_n444), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(new_n456), .A3(new_n453), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n435), .A2(new_n438), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n437), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n455), .B(new_n457), .C1(new_n459), .C2(new_n439), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n421), .B1(new_n451), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n460), .A2(new_n450), .A3(new_n295), .A4(new_n420), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G214), .B1(G237), .B2(G902), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n450), .A2(new_n295), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n467), .A2(KEYINPUT89), .A3(new_n420), .A4(new_n460), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n419), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n305), .A2(new_n310), .A3(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(KEYINPUT76), .B(KEYINPUT23), .C1(new_n195), .C2(G119), .ZN(new_n472));
  INV_X1    g286(.A(G119), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(G128), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n472), .B(new_n474), .C1(KEYINPUT76), .C2(KEYINPUT23), .ZN(new_n476));
  AOI21_X1  g290(.A(G110), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT24), .B(G110), .Z(new_n478));
  XNOR2_X1  g292(.A(G119), .B(G128), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n332), .B(new_n346), .C1(new_n477), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n479), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n475), .A2(new_n476), .ZN(new_n483));
  INV_X1    g297(.A(G110), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n486), .A2(KEYINPUT77), .A3(new_n333), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT77), .B1(new_n486), .B2(new_n333), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n481), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT22), .B(G137), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n312), .A2(G221), .A3(G234), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n490), .B(new_n491), .Z(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n481), .B(new_n492), .C1(new_n487), .C2(new_n488), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n385), .B1(G234), .B2(new_n295), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(G902), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT78), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n494), .A2(new_n495), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT25), .B1(new_n501), .B2(G902), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT25), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n494), .A2(new_n503), .A3(new_n295), .A4(new_n495), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n504), .A3(new_n496), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT79), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT79), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n500), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n247), .A2(KEYINPUT68), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n252), .A2(KEYINPUT68), .A3(G137), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n250), .ZN(new_n514));
  OAI21_X1  g328(.A(G131), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n259), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n516), .B1(new_n201), .B2(new_n238), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n232), .B1(new_n259), .B2(new_n257), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT73), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n442), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n251), .A2(new_n255), .A3(new_n258), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n258), .B1(new_n251), .B2(new_n255), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n231), .B(new_n230), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT73), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n523), .B(new_n524), .C1(new_n242), .C2(new_n516), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n519), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT28), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n523), .B(new_n520), .C1(new_n242), .C2(new_n516), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT67), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n523), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n233), .A2(new_n260), .A3(KEYINPUT67), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n517), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n531), .B1(new_n535), .B2(new_n520), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT28), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n526), .A2(KEYINPUT74), .A3(new_n527), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n530), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n311), .A2(G210), .A3(new_n312), .ZN(new_n540));
  XOR2_X1   g354(.A(KEYINPUT26), .B(G101), .Z(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n542), .A2(new_n543), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n523), .B(KEYINPUT30), .C1(new_n242), .C2(new_n516), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n442), .B(new_n549), .C1(new_n535), .C2(KEYINPUT30), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n547), .A2(KEYINPUT72), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n550), .A2(new_n551), .A3(new_n531), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n547), .A2(KEYINPUT31), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT31), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n554), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n557), .A2(new_n531), .A3(new_n550), .A4(new_n551), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n548), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT75), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n548), .A2(KEYINPUT75), .A3(new_n559), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(G472), .A2(G902), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT32), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n565), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT32), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n548), .A2(KEYINPUT75), .A3(new_n559), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT75), .B1(new_n548), .B2(new_n559), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT29), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n530), .A2(new_n537), .A3(new_n573), .A4(new_n538), .ZN(new_n574));
  INV_X1    g388(.A(new_n538), .ZN(new_n575));
  AOI21_X1  g389(.A(KEYINPUT74), .B1(new_n526), .B2(new_n527), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n442), .B1(new_n517), .B2(new_n518), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n527), .B1(new_n577), .B2(new_n531), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n546), .B(new_n574), .C1(new_n579), .C2(new_n573), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n550), .A2(new_n531), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(new_n546), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n582), .B2(new_n573), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(G472), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n572), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n511), .B1(new_n566), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT80), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n567), .B1(new_n562), .B2(new_n563), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n572), .B(new_n585), .C1(new_n590), .C2(KEYINPUT32), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(KEYINPUT80), .A3(new_n511), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n471), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT99), .B(G101), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G3));
  AOI21_X1  g409(.A(new_n303), .B1(new_n292), .B2(G469), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n309), .B1(new_n596), .B2(new_n302), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n295), .B1(new_n570), .B2(new_n571), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT100), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n564), .A2(KEYINPUT100), .A3(new_n295), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n601), .A3(G472), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n510), .A2(new_n590), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n597), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT101), .ZN(new_n605));
  INV_X1    g419(.A(new_n466), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n464), .A2(KEYINPUT102), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n607), .A2(new_n462), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n467), .A2(new_n609), .A3(new_n420), .A4(new_n460), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n606), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n418), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n361), .A2(new_n411), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n391), .A2(new_n392), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n390), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n615), .B1(new_n384), .B2(new_n386), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n617), .B1(new_n384), .B2(new_n386), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n392), .A2(G902), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n614), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n613), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n612), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n605), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT34), .B(G104), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  INV_X1    g441(.A(new_n397), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n628), .A2(new_n361), .A3(new_n411), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n612), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n605), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  INV_X1    g447(.A(new_n471), .ZN(new_n634));
  INV_X1    g448(.A(G472), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n598), .B2(new_n599), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n590), .B1(new_n636), .B2(new_n601), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n493), .A2(KEYINPUT36), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n489), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n497), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n505), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n634), .A2(new_n637), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT37), .B(G110), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G12));
  NAND3_X1  g458(.A1(new_n305), .A2(new_n310), .A3(new_n611), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n566), .A2(new_n586), .ZN(new_n646));
  INV_X1    g460(.A(new_n641), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT103), .B(G900), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n416), .B1(new_n649), .B2(new_n413), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n629), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  XOR2_X1   g467(.A(new_n650), .B(KEYINPUT39), .Z(new_n654));
  NAND2_X1  g468(.A1(new_n597), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(KEYINPUT40), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n570), .A2(new_n571), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n568), .B1(new_n659), .B2(new_n567), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n581), .A2(new_n546), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n577), .A2(new_n531), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(G902), .B1(new_n663), .B2(new_n547), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n660), .B(new_n572), .C1(new_n635), .C2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n465), .A2(new_n468), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n613), .A2(new_n628), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n670), .A2(new_n606), .A3(new_n641), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n666), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n658), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT106), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n658), .A2(new_n675), .A3(new_n672), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n316), .ZN(G45));
  INV_X1    g493(.A(new_n650), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n408), .A2(new_n410), .ZN(new_n681));
  INV_X1    g495(.A(G475), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n357), .B2(new_n359), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n622), .B(new_n680), .C1(new_n681), .C2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n648), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  AOI21_X1  g501(.A(new_n272), .B1(new_n265), .B2(new_n263), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n299), .B1(new_n688), .B2(new_n298), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n301), .B1(new_n689), .B2(KEYINPUT85), .ZN(new_n690));
  OAI21_X1  g504(.A(G469), .B1(new_n690), .B2(G902), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n302), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n309), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n694), .A2(new_n587), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n624), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n630), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  INV_X1    g514(.A(new_n419), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n646), .A2(new_n647), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n691), .A2(new_n302), .A3(new_n611), .A4(new_n310), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n701), .B(new_n702), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  NOR2_X1   g522(.A1(new_n612), .A2(new_n670), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n559), .B1(new_n546), .B2(new_n579), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n565), .B(KEYINPUT109), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n598), .A2(G472), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n713));
  INV_X1    g527(.A(new_n506), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n693), .B(new_n709), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G122), .ZN(G24));
  AND3_X1   g532(.A1(new_n712), .A2(new_n641), .A3(new_n685), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n705), .B2(new_n706), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G125), .ZN(G27));
  AOI22_X1  g535(.A1(new_n564), .A2(new_n569), .B1(G472), .B2(new_n584), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n510), .B1(new_n722), .B2(new_n660), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n606), .B1(new_n465), .B2(new_n468), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(new_n597), .A3(new_n685), .A4(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n684), .A2(new_n726), .ZN(new_n727));
  AND4_X1   g541(.A1(new_n310), .A2(new_n727), .A3(new_n305), .A4(new_n724), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n646), .A2(new_n506), .ZN(new_n729));
  AOI22_X1  g543(.A1(new_n725), .A2(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n258), .ZN(G33));
  AND4_X1   g545(.A1(new_n723), .A2(new_n597), .A3(new_n651), .A4(new_n724), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n252), .ZN(G36));
  INV_X1    g547(.A(new_n724), .ZN(new_n734));
  INV_X1    g548(.A(new_n613), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n622), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT43), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n637), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n738), .A2(new_n739), .A3(new_n641), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n734), .B1(new_n740), .B2(KEYINPUT44), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT112), .ZN(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n292), .B2(KEYINPUT45), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n743), .B1(KEYINPUT45), .B2(new_n292), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n303), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT111), .ZN(new_n746));
  OR3_X1    g560(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT46), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n746), .B1(new_n745), .B2(KEYINPUT46), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(KEYINPUT46), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n747), .A2(new_n302), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n310), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n740), .A2(KEYINPUT44), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n742), .A2(new_n654), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G137), .ZN(G39));
  NOR4_X1   g569(.A1(new_n591), .A2(new_n511), .A3(new_n684), .A4(new_n734), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n750), .A2(KEYINPUT47), .A3(new_n310), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT47), .B1(new_n750), .B2(new_n310), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT113), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n761), .B(new_n756), .C1(new_n757), .C2(new_n758), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G140), .ZN(G42));
  OR4_X1    g578(.A1(new_n506), .A2(new_n736), .A3(new_n309), .A4(new_n606), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n692), .B(KEYINPUT49), .ZN(new_n766));
  OR4_X1    g580(.A1(new_n666), .A2(new_n765), .A3(new_n766), .A4(new_n669), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n694), .A2(new_n734), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n769), .A2(new_n510), .A3(new_n417), .A4(new_n666), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n613), .A2(new_n622), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n738), .A2(new_n416), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT116), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n715), .A2(new_n716), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n694), .A2(new_n466), .A3(new_n669), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n779));
  AOI22_X1  g593(.A1(new_n776), .A2(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n777), .A2(new_n775), .A3(new_n778), .A4(new_n779), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n768), .A2(new_n641), .A3(new_n712), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n772), .B(new_n780), .C1(new_n774), .C2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n692), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n309), .B1(new_n785), .B2(KEYINPUT117), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(KEYINPUT117), .B2(new_n785), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n757), .A2(new_n758), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n776), .A2(new_n724), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n784), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n465), .A2(new_n466), .A3(new_n468), .A4(new_n418), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n623), .B2(new_n629), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n597), .A2(new_n602), .A3(new_n603), .A4(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n305), .A2(new_n470), .A3(new_n310), .A4(new_n641), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n798), .B1(new_n739), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n795), .B1(new_n800), .B2(new_n593), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n591), .A2(KEYINPUT80), .A3(new_n511), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT80), .B1(new_n591), .B2(new_n511), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n634), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n642), .A3(KEYINPUT114), .A4(new_n798), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  OAI211_X1 g620(.A(new_n723), .B(new_n693), .C1(new_n624), .C2(new_n630), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n707), .A2(new_n717), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n597), .A2(new_n641), .A3(new_n724), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n712), .A2(new_n685), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n591), .A2(new_n397), .A3(new_n735), .A4(new_n680), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n730), .A2(new_n813), .A3(new_n732), .ZN(new_n814));
  AND4_X1   g628(.A1(new_n794), .A2(new_n806), .A3(new_n809), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n808), .B1(new_n801), .B2(new_n805), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n794), .B1(new_n816), .B2(new_n814), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n645), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n819), .B(new_n702), .C1(new_n651), .C2(new_n685), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n611), .A2(new_n628), .A3(new_n613), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n821), .A2(new_n641), .A3(new_n650), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(new_n597), .A3(new_n666), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(new_n720), .A3(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n820), .A2(new_n720), .A3(KEYINPUT52), .A4(new_n823), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT53), .B1(new_n818), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(KEYINPUT53), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n815), .A2(new_n817), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT54), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n816), .A2(new_n814), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(KEYINPUT115), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n816), .A2(new_n794), .A3(new_n814), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n828), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n830), .A2(new_n833), .ZN(new_n840));
  INV_X1    g654(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n838), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n832), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n774), .A2(new_n729), .A3(new_n768), .ZN(new_n844));
  XOR2_X1   g658(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n845));
  OR2_X1    g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n776), .B1(new_n705), .B2(new_n706), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n844), .A2(new_n845), .ZN(new_n848));
  INV_X1    g662(.A(G952), .ZN(new_n849));
  INV_X1    g663(.A(new_n623), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n849), .B(G953), .C1(new_n770), .C2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n846), .A2(new_n847), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n792), .A2(new_n793), .A3(new_n843), .A4(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(G952), .A2(G953), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n767), .B1(new_n853), .B2(new_n854), .ZN(G75));
  NOR2_X1   g669(.A1(new_n829), .A2(new_n840), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n295), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT56), .B1(new_n857), .B2(G210), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n459), .A2(new_n439), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n455), .A2(new_n457), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n460), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT55), .Z(new_n863));
  AND2_X1   g677(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n858), .A2(new_n863), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n849), .A2(G953), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT120), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n864), .A2(new_n865), .A3(new_n868), .ZN(G51));
  OAI21_X1  g683(.A(KEYINPUT54), .B1(new_n829), .B2(new_n840), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n842), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n303), .B(KEYINPUT57), .Z(new_n873));
  OAI22_X1  g687(.A1(new_n872), .A2(new_n873), .B1(new_n300), .B2(new_n301), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n857), .A2(new_n744), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n868), .B1(new_n874), .B2(new_n875), .ZN(G54));
  NAND3_X1  g690(.A1(new_n857), .A2(KEYINPUT58), .A3(G475), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n877), .A2(new_n404), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n404), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n868), .B1(new_n878), .B2(new_n879), .ZN(G60));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n881));
  XNOR2_X1  g695(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n392), .A2(new_n295), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n882), .B(new_n883), .Z(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n832), .B2(new_n842), .ZN(new_n885));
  INV_X1    g699(.A(new_n619), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n881), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n884), .ZN(new_n888));
  INV_X1    g702(.A(new_n831), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n839), .B1(new_n889), .B2(new_n838), .ZN(new_n890));
  AOI211_X1 g704(.A(KEYINPUT54), .B(new_n840), .C1(new_n836), .C2(new_n837), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(KEYINPUT122), .A3(new_n619), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n619), .A2(new_n884), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n868), .B1(new_n871), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n887), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n887), .A2(new_n893), .A3(KEYINPUT123), .A4(new_n895), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(G63));
  NAND2_X1  g714(.A1(G217), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT124), .Z(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT60), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n856), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(new_n639), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n501), .B1(new_n856), .B2(new_n903), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n867), .A3(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(G66));
  INV_X1    g723(.A(G224), .ZN(new_n910));
  OAI21_X1  g724(.A(G953), .B1(new_n414), .B2(new_n910), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT125), .Z(new_n912));
  INV_X1    g726(.A(new_n816), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(new_n312), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n860), .B1(G898), .B2(new_n312), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n914), .B(new_n915), .Z(G69));
  OAI21_X1  g730(.A(new_n549), .B1(new_n535), .B2(KEYINPUT30), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(new_n399), .Z(new_n918));
  INV_X1    g732(.A(G900), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n919), .B2(new_n312), .ZN(new_n920));
  INV_X1    g734(.A(new_n754), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n760), .B2(new_n762), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n646), .A2(new_n506), .A3(new_n821), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n752), .A2(new_n654), .A3(new_n923), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n820), .A2(new_n720), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n730), .A2(new_n732), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n920), .B1(new_n928), .B2(new_n312), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n674), .A2(new_n676), .A3(new_n925), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT62), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n674), .A2(KEYINPUT62), .A3(new_n676), .A4(new_n925), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n589), .A2(new_n592), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n623), .A2(new_n629), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n657), .A2(new_n935), .A3(new_n724), .A4(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n934), .A2(new_n922), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n918), .B1(new_n938), .B2(new_n312), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n312), .B1(G227), .B2(G900), .ZN(new_n940));
  OR3_X1    g754(.A1(new_n929), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n929), .B2(new_n939), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(G72));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n934), .A2(new_n922), .A3(new_n816), .A4(new_n937), .ZN(new_n945));
  NAND2_X1  g759(.A1(G472), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT63), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n661), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI211_X1 g764(.A(KEYINPUT126), .B(new_n661), .C1(new_n945), .C2(new_n947), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n889), .A2(new_n838), .ZN(new_n953));
  INV_X1    g767(.A(new_n947), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n949), .A2(new_n582), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n868), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n763), .A2(new_n754), .A3(new_n816), .A4(new_n927), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n947), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n582), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n958), .A2(new_n959), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n956), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n952), .A2(new_n963), .ZN(G57));
endmodule


