//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n202));
  AND2_X1   g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  OR3_X1    g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT26), .ZN(new_n205));
  AOI22_X1  g004(.A1(new_n204), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n207));
  AOI21_X1  g006(.A(G190gat), .B1(new_n207), .B2(KEYINPUT27), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT27), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT28), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT27), .ZN(new_n214));
  INV_X1    g013(.A(G190gat), .ZN(new_n215));
  AND4_X1   g014(.A1(KEYINPUT28), .A2(new_n212), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n205), .B(new_n206), .C1(new_n211), .C2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G190gat), .ZN(new_n220));
  NOR2_X1   g019(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n218), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT23), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT25), .ZN(new_n230));
  NOR4_X1   g029(.A1(new_n222), .A2(new_n229), .A3(KEYINPUT65), .A4(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n219), .A2(G190gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n215), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n233));
  OR2_X1    g032(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n225), .A2(new_n227), .A3(KEYINPUT65), .A4(new_n228), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n235), .A2(new_n236), .B1(new_n237), .B2(KEYINPUT25), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n217), .B1(new_n231), .B2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(G127gat), .B(G134gat), .Z(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(KEYINPUT1), .B2(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(G113gat), .B(G120gat), .Z(new_n243));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n244));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n239), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n242), .A2(new_n246), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n249), .B(new_n217), .C1(new_n231), .C2(new_n238), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G227gat), .A2(G233gat), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n252), .B(KEYINPUT64), .Z(new_n253));
  AOI21_X1  g052(.A(new_n202), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  AOI211_X1 g054(.A(KEYINPUT67), .B(new_n255), .C1(new_n248), .C2(new_n250), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT32), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G15gat), .B(G43gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(G71gat), .B(G99gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  OR2_X1    g060(.A1(new_n261), .A2(KEYINPUT69), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(KEYINPUT69), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n262), .A2(KEYINPUT33), .A3(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT68), .ZN(new_n267));
  INV_X1    g066(.A(new_n250), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n223), .A2(new_n224), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n203), .B1(new_n269), .B2(new_n226), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n234), .A2(G190gat), .A3(new_n219), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n270), .A2(new_n271), .A3(new_n225), .A4(new_n218), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n237), .A2(KEYINPUT25), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT25), .A4(new_n237), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n249), .B1(new_n276), .B2(new_n217), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n253), .B1(new_n268), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT67), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n251), .A2(new_n202), .A3(new_n253), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n260), .B1(new_n281), .B2(KEYINPUT32), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT33), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(new_n254), .B2(new_n256), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n267), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AND4_X1   g084(.A1(new_n267), .A2(new_n257), .A3(new_n284), .A4(new_n261), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n266), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT34), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n248), .A2(new_n288), .A3(new_n250), .A4(new_n255), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n251), .B1(G227gat), .B2(G233gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(new_n288), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G155gat), .ZN(new_n293));
  INV_X1    g092(.A(G162gat), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT2), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G141gat), .ZN(new_n296));
  INV_X1    g095(.A(G148gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n295), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G155gat), .B(G162gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT75), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n298), .A2(new_n303), .A3(new_n299), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(G141gat), .B(G148gat), .Z(new_n306));
  OAI211_X1 g105(.A(new_n306), .B(new_n295), .C1(new_n303), .C2(new_n301), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(G211gat), .B(G218gat), .Z(new_n312));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n313));
  AND2_X1   g112(.A1(G197gat), .A2(G204gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(G197gat), .A2(G204gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n313), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G197gat), .ZN(new_n319));
  INV_X1    g118(.A(G204gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G197gat), .A2(G204gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n317), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(KEYINPUT70), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n312), .B1(new_n318), .B2(new_n325), .ZN(new_n326));
  NOR3_X1   g125(.A1(new_n316), .A2(new_n313), .A3(new_n317), .ZN(new_n327));
  INV_X1    g126(.A(new_n312), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n311), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G228gat), .ZN(new_n332));
  INV_X1    g131(.A(G233gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n305), .A2(new_n307), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n326), .B2(new_n329), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n337), .B1(new_n339), .B2(new_n308), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT79), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT70), .B1(new_n323), .B2(new_n324), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n328), .B1(new_n327), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n312), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT29), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n336), .B1(new_n345), .B2(KEYINPUT3), .ZN(new_n346));
  INV_X1    g145(.A(new_n334), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(new_n311), .B2(new_n330), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n343), .A2(new_n344), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT3), .B1(new_n351), .B2(new_n310), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n331), .B1(new_n352), .B2(new_n337), .ZN(new_n353));
  AOI22_X1  g152(.A1(new_n341), .A2(new_n350), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G22gat), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT81), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n347), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n335), .A2(new_n340), .A3(KEYINPUT79), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n349), .B1(new_n346), .B2(new_n348), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n361), .A3(G22gat), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n355), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n341), .A2(new_n350), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n366), .A2(KEYINPUT80), .A3(new_n355), .A4(new_n357), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n356), .A2(new_n362), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G78gat), .B(G106gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(KEYINPUT31), .B(G50gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n369), .B(new_n370), .Z(new_n371));
  NAND2_X1  g170(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n354), .A2(new_n355), .ZN(new_n373));
  INV_X1    g172(.A(new_n363), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n373), .A2(new_n374), .A3(new_n371), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n257), .A2(new_n284), .A3(new_n261), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT68), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n282), .A2(new_n267), .A3(new_n284), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n291), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n382), .A3(new_n266), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n292), .A2(new_n377), .A3(KEYINPUT88), .A4(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT35), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT73), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT71), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n239), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n276), .A2(KEYINPUT71), .A3(new_n217), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n310), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n392), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n239), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n387), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT73), .B1(new_n391), .B2(new_n392), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n330), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n389), .A2(new_n390), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n394), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n239), .A2(new_n338), .A3(new_n392), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n351), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT74), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT74), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n398), .A2(new_n406), .A3(new_n403), .ZN(new_n407));
  XNOR2_X1  g206(.A(G8gat), .B(G36gat), .ZN(new_n408));
  XNOR2_X1  g207(.A(G64gat), .B(G92gat), .ZN(new_n409));
  XOR2_X1   g208(.A(new_n408), .B(new_n409), .Z(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n405), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n398), .A2(new_n403), .A3(new_n410), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n413), .A2(new_n414), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n412), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n382), .B1(new_n381), .B2(new_n266), .ZN(new_n419));
  AOI211_X1 g218(.A(new_n291), .B(new_n265), .C1(new_n379), .C2(new_n380), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n309), .A2(new_n247), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n336), .A2(KEYINPUT3), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT77), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n249), .A2(new_n426), .A3(new_n307), .A4(new_n305), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT77), .B1(new_n336), .B2(new_n247), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT4), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n336), .A2(new_n247), .ZN(new_n430));
  XOR2_X1   g229(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n422), .B(new_n425), .C1(new_n429), .C2(new_n432), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n427), .B(new_n428), .C1(new_n249), .C2(new_n337), .ZN(new_n434));
  INV_X1    g233(.A(new_n422), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(KEYINPUT5), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n427), .A2(new_n428), .A3(KEYINPUT4), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n430), .A2(new_n431), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n438), .A2(new_n439), .B1(new_n424), .B2(new_n423), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n435), .A2(KEYINPUT5), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n440), .A2(KEYINPUT78), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT78), .B1(new_n440), .B2(new_n441), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n437), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G1gat), .B(G29gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT0), .ZN(new_n446));
  XNOR2_X1  g245(.A(G57gat), .B(G85gat), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n446), .B(new_n447), .Z(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n437), .B(new_n448), .C1(new_n442), .C2(new_n443), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n444), .A2(KEYINPUT6), .A3(new_n449), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n418), .A2(new_n421), .A3(new_n455), .A4(new_n377), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n386), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n292), .A2(new_n383), .A3(new_n377), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n452), .A2(new_n451), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n438), .A2(new_n439), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n460), .A2(new_n425), .A3(new_n441), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT78), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n440), .A2(KEYINPUT78), .A3(new_n441), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n448), .B1(new_n465), .B2(new_n437), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n459), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n454), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n458), .A2(new_n469), .A3(new_n417), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n384), .A2(new_n385), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n474));
  NAND3_X1  g273(.A1(new_n398), .A2(new_n403), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n351), .B1(new_n396), .B2(new_n397), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n402), .A2(new_n330), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(KEYINPUT37), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT38), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n475), .A2(new_n478), .A3(new_n479), .A4(new_n411), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n453), .A2(new_n454), .A3(new_n413), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT86), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n469), .A2(new_n484), .A3(new_n413), .A4(new_n480), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n405), .A2(KEYINPUT37), .A3(new_n407), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n411), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT87), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n487), .A2(KEYINPUT87), .A3(new_n411), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n491), .A3(new_n475), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n486), .B1(new_n492), .B2(KEYINPUT38), .ZN(new_n493));
  OR3_X1    g292(.A1(new_n440), .A2(KEYINPUT39), .A3(new_n422), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n440), .A2(new_n422), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT39), .B1(new_n434), .B2(new_n435), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n494), .B(new_n448), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT40), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n466), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n497), .A2(new_n498), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n500), .A2(KEYINPUT84), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(KEYINPUT84), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n377), .B1(new_n418), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n493), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n455), .A2(new_n412), .A3(new_n415), .A4(new_n416), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n377), .A2(KEYINPUT82), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n375), .B1(new_n368), .B2(new_n371), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT82), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT36), .B1(new_n419), .B2(new_n420), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n292), .A2(new_n514), .A3(new_n383), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n506), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n507), .A2(new_n508), .A3(new_n511), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n518), .A2(KEYINPUT83), .A3(new_n513), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n473), .B1(new_n505), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT97), .B(G85gat), .ZN(new_n522));
  INV_X1    g321(.A(G92gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n522), .A2(new_n523), .B1(KEYINPUT8), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(G85gat), .A2(G92gat), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(KEYINPUT96), .B2(KEYINPUT7), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT7), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n528), .A2(new_n529), .A3(G85gat), .A4(G92gat), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n527), .B(new_n530), .C1(new_n528), .C2(new_n529), .ZN(new_n531));
  XNOR2_X1  g330(.A(G99gat), .B(G106gat), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n525), .B(new_n531), .C1(KEYINPUT98), .C2(new_n532), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n532), .A2(KEYINPUT98), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(KEYINPUT99), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G29gat), .A2(G36gat), .ZN(new_n538));
  NOR3_X1   g337(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT90), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n542), .B1(new_n539), .B2(new_n540), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n538), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G43gat), .B(G50gat), .Z(new_n545));
  INV_X1    g344(.A(KEYINPUT89), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G43gat), .B(G50gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT89), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n544), .A2(KEYINPUT15), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n547), .A2(KEYINPUT15), .A3(new_n549), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n539), .A2(KEYINPUT91), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n539), .A2(KEYINPUT91), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n542), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT15), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n545), .A2(new_n555), .B1(G29gat), .B2(G36gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n551), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT17), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n537), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n536), .A2(new_n558), .ZN(new_n561));
  NAND3_X1  g360(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n562));
  AND3_X1   g361(.A1(new_n561), .A2(KEYINPUT100), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT100), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G190gat), .B(G218gat), .Z(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n565), .A2(new_n566), .ZN(new_n569));
  XNOR2_X1  g368(.A(G134gat), .B(G162gat), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n570), .B(new_n571), .Z(new_n572));
  AOI22_X1  g371(.A1(new_n568), .A2(new_n569), .B1(KEYINPUT101), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n572), .B(KEYINPUT101), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n568), .A2(new_n569), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(G71gat), .A2(G78gat), .ZN(new_n578));
  NOR2_X1   g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(G57gat), .B(G64gat), .Z(new_n581));
  AOI21_X1  g380(.A(new_n580), .B1(new_n581), .B2(KEYINPUT94), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(KEYINPUT9), .B2(new_n578), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(G127gat), .ZN(new_n588));
  XOR2_X1   g387(.A(G183gat), .B(G211gat), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(G8gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(G15gat), .B(G22gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT16), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n592), .B1(new_n593), .B2(G1gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT92), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n591), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n594), .B1(G1gat), .B2(new_n592), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n600), .B1(KEYINPUT21), .B2(new_n584), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT95), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(new_n293), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n602), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n590), .B(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n577), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n535), .B(new_n584), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT10), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n536), .A2(KEYINPUT10), .A3(new_n584), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT102), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n608), .A2(new_n613), .ZN(new_n616));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n617), .B(new_n618), .Z(new_n619));
  NAND3_X1  g418(.A1(new_n615), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT103), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n615), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n611), .A2(KEYINPUT103), .A3(new_n614), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n622), .A2(new_n623), .B1(new_n613), .B2(new_n608), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n620), .B1(new_n624), .B2(new_n619), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n600), .A2(new_n558), .ZN(new_n628));
  INV_X1    g427(.A(new_n600), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n628), .B1(new_n559), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G229gat), .A2(G233gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n633));
  OR2_X1    g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n600), .B(new_n558), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n631), .B(KEYINPUT13), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n634), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G113gat), .B(G141gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G197gat), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT11), .B(G169gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT12), .Z(new_n644));
  NAND2_X1  g443(.A1(new_n639), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n634), .A2(new_n646), .A3(new_n635), .A4(new_n638), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n627), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n521), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n469), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g453(.A(new_n591), .B1(new_n652), .B2(new_n417), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G8gat), .ZN(new_n657));
  NOR3_X1   g456(.A1(new_n651), .A2(new_n418), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT42), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(KEYINPUT42), .B2(new_n658), .ZN(G1325gat));
  INV_X1    g459(.A(new_n421), .ZN(new_n661));
  OR3_X1    g460(.A1(new_n651), .A2(G15gat), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n516), .ZN(new_n663));
  OAI21_X1  g462(.A(G15gat), .B1(new_n651), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT105), .ZN(G1326gat));
  AND2_X1   g465(.A1(new_n508), .A2(new_n511), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n651), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT43), .B(G22gat), .Z(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  AND2_X1   g470(.A1(new_n521), .A2(new_n577), .ZN(new_n672));
  INV_X1    g471(.A(new_n606), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n625), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n649), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NOR3_X1   g476(.A1(new_n677), .A2(G29gat), .A3(new_n455), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT45), .Z(new_n679));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n648), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT107), .B1(new_n457), .B2(new_n472), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n512), .A2(new_n516), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n493), .B2(new_n504), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n386), .A2(new_n456), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n470), .A2(new_n471), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n684), .A2(new_n686), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT108), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n684), .A2(new_n686), .A3(new_n693), .A4(new_n690), .ZN(new_n694));
  INV_X1    g493(.A(new_n577), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n695), .A2(KEYINPUT44), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n692), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n521), .A2(new_n577), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT44), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n683), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(G29gat), .B1(new_n701), .B2(new_n455), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n679), .A2(new_n702), .ZN(G1328gat));
  NOR2_X1   g502(.A1(new_n418), .A2(G36gat), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT109), .B1(new_n677), .B2(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n698), .A2(new_n649), .A3(new_n675), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n707), .A2(new_n708), .A3(new_n704), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n706), .B(new_n709), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(KEYINPUT110), .B2(KEYINPUT46), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n706), .A2(new_n709), .A3(new_n710), .A4(new_n711), .ZN(new_n714));
  OAI21_X1  g513(.A(G36gat), .B1(new_n701), .B2(new_n418), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(G1329gat));
  NOR3_X1   g515(.A1(new_n677), .A2(G43gat), .A3(new_n661), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n663), .B(new_n683), .C1(new_n697), .C2(new_n699), .ZN(new_n720));
  OAI21_X1  g519(.A(G43gat), .B1(new_n720), .B2(KEYINPUT111), .ZN(new_n721));
  AND3_X1   g520(.A1(new_n700), .A2(KEYINPUT111), .A3(new_n516), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(G43gat), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n718), .B1(new_n725), .B2(new_n717), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(G1330gat));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728));
  INV_X1    g527(.A(G50gat), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n729), .B1(new_n700), .B2(new_n667), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n668), .A2(G50gat), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n672), .A2(new_n676), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n728), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n697), .A2(new_n699), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n509), .A3(new_n682), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G50gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n732), .A2(KEYINPUT48), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n735), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  AOI211_X1 g540(.A(KEYINPUT112), .B(new_n739), .C1(new_n737), .C2(G50gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n734), .B1(new_n741), .B2(new_n742), .ZN(G1331gat));
  AND2_X1   g542(.A1(new_n692), .A2(new_n694), .ZN(new_n744));
  INV_X1    g543(.A(new_n607), .ZN(new_n745));
  INV_X1    g544(.A(new_n681), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n745), .A2(new_n626), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n744), .A2(new_n469), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G57gat), .ZN(G1332gat));
  NAND3_X1  g548(.A1(new_n744), .A2(new_n417), .A3(new_n747), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT49), .B(G64gat), .Z(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n750), .B2(new_n752), .ZN(G1333gat));
  NAND3_X1  g552(.A1(new_n744), .A2(new_n516), .A3(new_n747), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G71gat), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n661), .A2(G71gat), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n744), .A2(new_n747), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1334gat));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n667), .A3(new_n747), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g561(.A1(new_n681), .A2(new_n606), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n625), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n736), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT113), .B1(new_n767), .B2(new_n455), .ZN(new_n768));
  INV_X1    g567(.A(new_n522), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n767), .A2(KEYINPUT113), .A3(new_n455), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n577), .B1(KEYINPUT114), .B2(KEYINPUT51), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n772), .A2(new_n763), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n691), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n625), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n469), .A2(new_n522), .ZN(new_n778));
  OAI22_X1  g577(.A1(new_n770), .A2(new_n771), .B1(new_n777), .B2(new_n778), .ZN(G1336gat));
  OAI21_X1  g578(.A(G92gat), .B1(new_n767), .B2(new_n418), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n417), .A2(new_n523), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n780), .B(new_n781), .C1(new_n777), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n777), .A2(new_n782), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n765), .B1(new_n697), .B2(new_n699), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n523), .B1(new_n785), .B2(new_n417), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT52), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n783), .A2(new_n787), .ZN(G1337gat));
  OAI21_X1  g587(.A(G99gat), .B1(new_n767), .B2(new_n663), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n626), .A2(new_n661), .A3(G99gat), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT115), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(G1338gat));
  INV_X1    g592(.A(new_n777), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n377), .A2(G106gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n785), .A2(new_n667), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n794), .A2(new_n795), .B1(new_n796), .B2(G106gat), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  INV_X1    g597(.A(G106gat), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n785), .B2(new_n509), .ZN(new_n800));
  INV_X1    g599(.A(new_n795), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n798), .B1(new_n777), .B2(new_n801), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n797), .A2(new_n798), .B1(new_n800), .B2(new_n802), .ZN(G1339gat));
  NAND3_X1  g602(.A1(new_n607), .A2(new_n626), .A3(new_n681), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n630), .A2(new_n631), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n636), .A2(new_n637), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n643), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n647), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  INV_X1    g610(.A(new_n576), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n573), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT103), .B1(new_n611), .B2(new_n614), .ZN(new_n815));
  AOI211_X1 g614(.A(new_n621), .B(new_n613), .C1(new_n609), .C2(new_n610), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n815), .A2(new_n816), .A3(KEYINPUT54), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n609), .A2(new_n613), .A3(new_n610), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n615), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n619), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n814), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n622), .A2(new_n823), .A3(new_n623), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n824), .A2(KEYINPUT55), .A3(new_n820), .A4(new_n819), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n620), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n813), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n625), .A2(new_n808), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n681), .B2(new_n826), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n577), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(KEYINPUT117), .B(new_n828), .C1(new_n681), .C2(new_n826), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n827), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n804), .B1(new_n833), .B2(new_n673), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n458), .A2(new_n417), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n469), .A3(new_n835), .ZN(new_n836));
  OR3_X1    g635(.A1(new_n836), .A2(G113gat), .A3(new_n681), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n667), .A2(new_n661), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n417), .A2(new_n455), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n648), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n842));
  AND3_X1   g641(.A1(new_n841), .A2(new_n842), .A3(G113gat), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n841), .B2(G113gat), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n837), .B1(new_n843), .B2(new_n844), .ZN(G1340gat));
  NAND2_X1  g644(.A1(new_n839), .A2(new_n840), .ZN(new_n846));
  INV_X1    g645(.A(G120gat), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n846), .A2(new_n847), .A3(new_n626), .ZN(new_n848));
  INV_X1    g647(.A(new_n836), .ZN(new_n849));
  AOI21_X1  g648(.A(G120gat), .B1(new_n849), .B2(new_n625), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n848), .A2(new_n850), .ZN(G1341gat));
  OAI21_X1  g650(.A(G127gat), .B1(new_n846), .B2(new_n606), .ZN(new_n852));
  OR3_X1    g651(.A1(new_n836), .A2(G127gat), .A3(new_n606), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1342gat));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n695), .A2(G134gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n849), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n856), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT119), .B1(new_n836), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n834), .A2(new_n577), .A3(new_n840), .A4(new_n838), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(G134gat), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT120), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n857), .A2(KEYINPUT56), .A3(new_n859), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n862), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n834), .A2(new_n868), .A3(new_n509), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n663), .A2(new_n840), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n813), .A2(new_n826), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n822), .A2(new_n825), .A3(new_n648), .A4(new_n620), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n828), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n695), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n673), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n804), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n667), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n870), .B1(new_n877), .B2(KEYINPUT57), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n869), .A2(new_n648), .A3(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n869), .A2(KEYINPUT121), .A3(new_n878), .A4(new_n648), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(G141gat), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n834), .A2(new_n469), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n516), .A2(new_n377), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(new_n417), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n884), .A2(new_n296), .A3(new_n648), .A4(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n883), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n869), .A2(new_n878), .ZN(new_n892));
  OAI21_X1  g691(.A(G141gat), .B1(new_n892), .B2(new_n681), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n888), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(KEYINPUT58), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n891), .A2(new_n895), .ZN(G1344gat));
  XOR2_X1   g695(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n297), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n887), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n901), .B2(new_n625), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n892), .A2(new_n626), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n829), .A2(new_n830), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n695), .A3(new_n832), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n673), .B1(new_n905), .B2(new_n871), .ZN(new_n906));
  OAI211_X1 g705(.A(KEYINPUT57), .B(new_n509), .C1(new_n906), .C2(new_n876), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n607), .A2(new_n649), .A3(new_n626), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n667), .B1(new_n875), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n911), .A3(new_n868), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n577), .B1(new_n872), .B2(new_n828), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n606), .B1(new_n913), .B2(new_n827), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n668), .B1(new_n914), .B2(new_n908), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT123), .B1(new_n915), .B2(KEYINPUT57), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n907), .A2(new_n912), .A3(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n663), .A2(new_n625), .A3(new_n840), .A4(new_n898), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n903), .A2(KEYINPUT59), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n902), .B1(new_n920), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g720(.A(G155gat), .B1(new_n892), .B2(new_n606), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n673), .A2(new_n293), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n900), .B2(new_n923), .ZN(G1346gat));
  NAND4_X1  g723(.A1(new_n884), .A2(new_n294), .A3(new_n577), .A4(new_n887), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT124), .ZN(new_n926));
  OAI21_X1  g725(.A(G162gat), .B1(new_n892), .B2(new_n695), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n418), .A2(new_n469), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n834), .A2(new_n648), .A3(new_n838), .A4(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(G169gat), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n834), .A2(new_n455), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n418), .A2(new_n458), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n746), .A2(new_n223), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(G1348gat));
  NAND3_X1  g737(.A1(new_n839), .A2(new_n625), .A3(new_n929), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(G176gat), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n625), .A2(new_n224), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n934), .B2(new_n941), .ZN(G1349gat));
  NAND3_X1  g741(.A1(new_n839), .A2(new_n673), .A3(new_n929), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(G183gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n673), .A2(new_n212), .A3(new_n214), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n934), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT60), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n943), .A2(G183gat), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n948), .B(new_n949), .C1(new_n934), .C2(new_n945), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n947), .A2(new_n950), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n839), .A2(new_n577), .A3(new_n929), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n952), .A2(new_n953), .A3(G190gat), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n953), .B1(new_n952), .B2(G190gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n577), .A2(new_n215), .ZN(new_n956));
  OAI22_X1  g755(.A1(new_n954), .A2(new_n955), .B1(new_n934), .B2(new_n956), .ZN(G1351gat));
  NOR3_X1   g756(.A1(new_n516), .A2(new_n469), .A3(new_n418), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n917), .A2(new_n648), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT127), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n917), .A2(new_n961), .A3(new_n648), .A4(new_n958), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n960), .A2(G197gat), .A3(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n886), .A2(new_n418), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n932), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n932), .A2(new_n967), .A3(new_n964), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n966), .A2(new_n319), .A3(new_n746), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n963), .A2(new_n969), .ZN(G1352gat));
  NAND4_X1  g769(.A1(new_n932), .A2(new_n320), .A3(new_n625), .A4(new_n964), .ZN(new_n971));
  OR2_X1    g770(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n917), .A2(new_n625), .A3(new_n958), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n972), .B(new_n973), .C1(new_n320), .C2(new_n974), .ZN(G1353gat));
  NAND3_X1  g774(.A1(new_n917), .A2(new_n673), .A3(new_n958), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n976), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  AOI21_X1  g776(.A(KEYINPUT63), .B1(new_n976), .B2(G211gat), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n966), .A2(new_n968), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n606), .A2(G211gat), .ZN(new_n980));
  OAI22_X1  g779(.A1(new_n977), .A2(new_n978), .B1(new_n979), .B2(new_n980), .ZN(G1354gat));
  NAND3_X1  g780(.A1(new_n917), .A2(new_n577), .A3(new_n958), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G218gat), .ZN(new_n983));
  OR2_X1    g782(.A1(new_n695), .A2(G218gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n979), .B2(new_n984), .ZN(G1355gat));
endmodule


