

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777;

  AND2_X1 U367 ( .A1(n382), .A2(n381), .ZN(n380) );
  NOR2_X1 U368 ( .A1(n408), .A2(KEYINPUT48), .ZN(n407) );
  NOR2_X1 U369 ( .A1(n561), .A2(n560), .ZN(n562) );
  INV_X1 U370 ( .A(n611), .ZN(n616) );
  INV_X1 U371 ( .A(G472), .ZN(n346) );
  INV_X2 U372 ( .A(G953), .ZN(n769) );
  NOR2_X2 U373 ( .A1(n581), .A2(n563), .ZN(n750) );
  XNOR2_X2 U374 ( .A(n347), .B(n346), .ZN(n620) );
  OR2_X2 U375 ( .A1(n697), .A2(G902), .ZN(n347) );
  XNOR2_X1 U376 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n455) );
  AND2_X2 U377 ( .A1(n375), .A2(n363), .ZN(n354) );
  OR2_X2 U378 ( .A1(n549), .A2(n564), .ZN(n464) );
  XNOR2_X1 U379 ( .A(n422), .B(n421), .ZN(n684) );
  XNOR2_X2 U380 ( .A(n600), .B(n599), .ZN(n619) );
  NOR2_X2 U381 ( .A1(n673), .A2(n613), .ZN(n424) );
  NOR2_X2 U382 ( .A1(n576), .A2(n556), .ZN(n522) );
  AND2_X1 U383 ( .A1(n554), .A2(n659), .ZN(n448) );
  NOR2_X2 U384 ( .A1(n552), .A2(n595), .ZN(n659) );
  XNOR2_X1 U385 ( .A(n761), .B(n507), .ZN(n516) );
  AND2_X1 U386 ( .A1(n439), .A2(KEYINPUT87), .ZN(n438) );
  NOR2_X1 U387 ( .A1(n392), .A2(n358), .ZN(n443) );
  AND2_X1 U388 ( .A1(n394), .A2(n428), .ZN(n379) );
  NOR2_X1 U389 ( .A1(n361), .A2(n368), .ZN(n364) );
  OR2_X1 U390 ( .A1(n630), .A2(KEYINPUT91), .ZN(n428) );
  XNOR2_X1 U391 ( .A(n623), .B(n622), .ZN(n747) );
  NAND2_X1 U392 ( .A1(n411), .A2(n409), .ZN(n447) );
  XOR2_X1 U393 ( .A(n565), .B(KEYINPUT38), .Z(n556) );
  BUF_X1 U394 ( .A(n559), .Z(n554) );
  XNOR2_X1 U395 ( .A(n469), .B(n459), .ZN(n697) );
  XNOR2_X1 U396 ( .A(n516), .B(n515), .ZN(n719) );
  XNOR2_X1 U397 ( .A(n455), .B(KEYINPUT3), .ZN(n385) );
  XNOR2_X1 U398 ( .A(KEYINPUT69), .B(G469), .ZN(n470) );
  XNOR2_X2 U399 ( .A(n656), .B(KEYINPUT6), .ZN(n611) );
  INV_X1 U400 ( .A(KEYINPUT74), .ZN(n445) );
  XNOR2_X1 U401 ( .A(G125), .B(G146), .ZN(n509) );
  AND2_X1 U402 ( .A1(n629), .A2(n628), .ZN(n630) );
  INV_X1 U403 ( .A(KEYINPUT46), .ZN(n376) );
  NAND2_X1 U404 ( .A1(n437), .A2(n436), .ZN(n417) );
  NAND2_X1 U405 ( .A1(n520), .A2(n688), .ZN(n436) );
  AND2_X1 U406 ( .A1(n402), .A2(n586), .ZN(n401) );
  NOR2_X1 U407 ( .A1(G953), .A2(G237), .ZN(n536) );
  NAND2_X1 U408 ( .A1(n417), .A2(n567), .ZN(n391) );
  NAND2_X1 U409 ( .A1(n448), .A2(n500), .ZN(n501) );
  OR2_X1 U410 ( .A1(n719), .A2(n434), .ZN(n433) );
  NAND2_X1 U411 ( .A1(n435), .A2(n687), .ZN(n434) );
  INV_X1 U412 ( .A(n520), .ZN(n435) );
  INV_X1 U413 ( .A(n417), .ZN(n416) );
  XNOR2_X1 U414 ( .A(n620), .B(KEYINPUT104), .ZN(n549) );
  XNOR2_X1 U415 ( .A(G110), .B(G137), .ZN(n479) );
  INV_X1 U416 ( .A(KEYINPUT23), .ZN(n481) );
  XOR2_X1 U417 ( .A(KEYINPUT10), .B(G140), .Z(n476) );
  BUF_X1 U418 ( .A(n549), .Z(n605) );
  NOR2_X1 U419 ( .A1(n769), .A2(G952), .ZN(n722) );
  NAND2_X1 U420 ( .A1(n367), .A2(n366), .ZN(n365) );
  NOR2_X1 U421 ( .A1(n568), .A2(n371), .ZN(n366) );
  NAND2_X1 U422 ( .A1(n370), .A2(n369), .ZN(n368) );
  NAND2_X1 U423 ( .A1(n568), .A2(n371), .ZN(n369) );
  NAND2_X1 U424 ( .A1(n674), .A2(n371), .ZN(n370) );
  NAND2_X1 U425 ( .A1(n365), .A2(n374), .ZN(n361) );
  AND2_X1 U426 ( .A1(n575), .A2(n446), .ZN(n431) );
  NAND2_X1 U427 ( .A1(G237), .A2(G234), .ZN(n494) );
  XOR2_X1 U428 ( .A(KEYINPUT14), .B(KEYINPUT93), .Z(n495) );
  NOR2_X1 U429 ( .A1(G902), .A2(G237), .ZN(n461) );
  AND2_X1 U430 ( .A1(n426), .A2(KEYINPUT44), .ZN(n425) );
  INV_X1 U431 ( .A(KEYINPUT28), .ZN(n415) );
  NAND2_X1 U432 ( .A1(n561), .A2(n415), .ZN(n414) );
  XNOR2_X1 U433 ( .A(n384), .B(n383), .ZN(n760) );
  XNOR2_X1 U434 ( .A(G107), .B(G104), .ZN(n384) );
  XNOR2_X1 U435 ( .A(G107), .B(G116), .ZN(n523) );
  AND2_X1 U436 ( .A1(n403), .A2(n348), .ZN(n398) );
  XOR2_X1 U437 ( .A(G113), .B(G104), .Z(n542) );
  XNOR2_X1 U438 ( .A(G143), .B(G122), .ZN(n541) );
  XOR2_X1 U439 ( .A(KEYINPUT99), .B(KEYINPUT12), .Z(n538) );
  XOR2_X1 U440 ( .A(G101), .B(G140), .Z(n466) );
  XNOR2_X1 U441 ( .A(KEYINPUT16), .B(G122), .ZN(n504) );
  XNOR2_X1 U442 ( .A(KEYINPUT66), .B(KEYINPUT4), .ZN(n450) );
  XNOR2_X1 U443 ( .A(n760), .B(KEYINPUT72), .ZN(n507) );
  NAND2_X1 U444 ( .A1(n447), .A2(n555), .ZN(n568) );
  INV_X1 U445 ( .A(KEYINPUT42), .ZN(n371) );
  AND2_X1 U446 ( .A1(n391), .A2(n389), .ZN(n388) );
  NAND2_X1 U447 ( .A1(n416), .A2(n351), .ZN(n387) );
  NAND2_X1 U448 ( .A1(n390), .A2(n567), .ZN(n389) );
  NAND2_X1 U449 ( .A1(n410), .A2(n413), .ZN(n409) );
  AND2_X1 U450 ( .A1(n412), .A2(n414), .ZN(n411) );
  NOR2_X1 U451 ( .A1(n561), .A2(n415), .ZN(n413) );
  XNOR2_X1 U452 ( .A(n554), .B(KEYINPUT106), .ZN(n555) );
  XNOR2_X1 U453 ( .A(n501), .B(KEYINPUT77), .ZN(n502) );
  XNOR2_X1 U454 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U455 ( .A(n475), .B(n474), .ZN(n477) );
  NAND2_X1 U456 ( .A1(n373), .A2(n372), .ZN(n363) );
  NOR2_X1 U457 ( .A1(n744), .A2(n356), .ZN(n372) );
  INV_X1 U458 ( .A(KEYINPUT36), .ZN(n399) );
  NOR2_X1 U459 ( .A1(n582), .A2(n565), .ZN(n400) );
  INV_X1 U460 ( .A(KEYINPUT35), .ZN(n421) );
  NOR2_X1 U461 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U462 ( .A1(n693), .A2(n722), .ZN(n694) );
  INV_X1 U463 ( .A(KEYINPUT53), .ZN(n418) );
  INV_X1 U464 ( .A(n368), .ZN(n362) );
  XNOR2_X1 U465 ( .A(n609), .B(n383), .ZN(G12) );
  AND2_X1 U466 ( .A1(n401), .A2(n688), .ZN(n348) );
  AND2_X1 U467 ( .A1(n646), .A2(n570), .ZN(n349) );
  AND2_X1 U468 ( .A1(n592), .A2(n555), .ZN(n350) );
  NAND2_X1 U469 ( .A1(n416), .A2(n433), .ZN(n565) );
  AND2_X1 U470 ( .A1(n433), .A2(n432), .ZN(n351) );
  XOR2_X1 U471 ( .A(n614), .B(KEYINPUT80), .Z(n352) );
  NOR2_X1 U472 ( .A1(n601), .A2(n616), .ZN(n353) );
  AND2_X1 U473 ( .A1(n447), .A2(n350), .ZN(n355) );
  NAND2_X1 U474 ( .A1(n388), .A2(n387), .ZN(n592) );
  XNOR2_X1 U475 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n356) );
  AND2_X1 U476 ( .A1(n375), .A2(n374), .ZN(n357) );
  OR2_X1 U477 ( .A1(KEYINPUT87), .A2(n687), .ZN(n358) );
  NAND2_X1 U478 ( .A1(n688), .A2(KEYINPUT2), .ZN(n359) );
  INV_X1 U479 ( .A(G110), .ZN(n383) );
  NAND2_X1 U480 ( .A1(n431), .A2(n574), .ZN(n430) );
  XNOR2_X2 U481 ( .A(n360), .B(n612), .ZN(n673) );
  NAND2_X1 U482 ( .A1(n395), .A2(n396), .ZN(n360) );
  NAND2_X1 U483 ( .A1(n562), .A2(n740), .ZN(n582) );
  OR2_X1 U484 ( .A1(n753), .A2(n392), .ZN(n640) );
  NAND2_X1 U485 ( .A1(n362), .A2(n365), .ZN(n777) );
  NAND2_X1 U486 ( .A1(n357), .A2(n363), .ZN(n776) );
  NAND2_X1 U487 ( .A1(n364), .A2(n354), .ZN(n377) );
  INV_X1 U488 ( .A(n674), .ZN(n367) );
  INV_X1 U489 ( .A(n580), .ZN(n373) );
  NAND2_X1 U490 ( .A1(n744), .A2(n356), .ZN(n374) );
  NAND2_X1 U491 ( .A1(n580), .A2(n356), .ZN(n375) );
  XNOR2_X2 U492 ( .A(n377), .B(n376), .ZN(n406) );
  XNOR2_X2 U493 ( .A(n378), .B(n635), .ZN(n753) );
  NAND2_X2 U494 ( .A1(n380), .A2(n379), .ZN(n378) );
  NAND2_X1 U495 ( .A1(n633), .A2(n632), .ZN(n381) );
  NAND2_X1 U496 ( .A1(n429), .A2(n427), .ZN(n382) );
  XNOR2_X2 U497 ( .A(n506), .B(n505), .ZN(n761) );
  XNOR2_X2 U498 ( .A(n386), .B(n385), .ZN(n506) );
  XNOR2_X2 U499 ( .A(n456), .B(n457), .ZN(n386) );
  NAND2_X1 U500 ( .A1(n433), .A2(n642), .ZN(n390) );
  NAND2_X1 U501 ( .A1(n403), .A2(n401), .ZN(n392) );
  XNOR2_X1 U502 ( .A(n392), .B(n771), .ZN(n770) );
  NAND2_X1 U503 ( .A1(n393), .A2(KEYINPUT48), .ZN(n404) );
  INV_X1 U504 ( .A(n406), .ZN(n393) );
  XNOR2_X1 U505 ( .A(n430), .B(n445), .ZN(n444) );
  NOR2_X2 U506 ( .A1(n640), .A2(n639), .ZN(n689) );
  XNOR2_X2 U507 ( .A(G119), .B(G116), .ZN(n456) );
  XNOR2_X2 U508 ( .A(n594), .B(n593), .ZN(n626) );
  INV_X1 U509 ( .A(n753), .ZN(n442) );
  NAND2_X1 U510 ( .A1(n631), .A2(n425), .ZN(n394) );
  INV_X1 U511 ( .A(n621), .ZN(n395) );
  INV_X1 U512 ( .A(n611), .ZN(n396) );
  XNOR2_X1 U513 ( .A(n544), .B(G137), .ZN(n451) );
  XNOR2_X2 U514 ( .A(G131), .B(KEYINPUT67), .ZN(n544) );
  NAND2_X1 U515 ( .A1(n444), .A2(n397), .ZN(n408) );
  XNOR2_X1 U516 ( .A(n750), .B(KEYINPUT89), .ZN(n397) );
  NAND2_X1 U517 ( .A1(n398), .A2(n442), .ZN(n439) );
  NAND2_X1 U518 ( .A1(n407), .A2(n406), .ZN(n405) );
  AND2_X2 U519 ( .A1(n405), .A2(n404), .ZN(n403) );
  XNOR2_X1 U520 ( .A(n400), .B(n399), .ZN(n563) );
  NAND2_X1 U521 ( .A1(n408), .A2(KEYINPUT48), .ZN(n402) );
  INV_X1 U522 ( .A(n605), .ZN(n410) );
  NAND2_X1 U523 ( .A1(n605), .A2(n415), .ZN(n412) );
  NAND2_X1 U524 ( .A1(n355), .A2(n349), .ZN(n571) );
  XNOR2_X1 U525 ( .A(n419), .B(n418), .ZN(G75) );
  NAND2_X1 U526 ( .A1(n420), .A2(n769), .ZN(n419) );
  XNOR2_X1 U527 ( .A(n680), .B(KEYINPUT122), .ZN(n420) );
  NAND2_X1 U528 ( .A1(n423), .A2(n352), .ZN(n422) );
  XNOR2_X1 U529 ( .A(n424), .B(KEYINPUT34), .ZN(n423) );
  NAND2_X1 U530 ( .A1(n631), .A2(KEYINPUT44), .ZN(n429) );
  INV_X1 U531 ( .A(KEYINPUT91), .ZN(n426) );
  AND2_X1 U532 ( .A1(n630), .A2(KEYINPUT91), .ZN(n427) );
  NOR2_X1 U533 ( .A1(n564), .A2(n567), .ZN(n432) );
  NAND2_X1 U534 ( .A1(n719), .A2(n520), .ZN(n437) );
  NOR2_X1 U535 ( .A1(n438), .A2(n440), .ZN(n690) );
  NAND2_X1 U536 ( .A1(n441), .A2(n359), .ZN(n440) );
  NAND2_X1 U537 ( .A1(n443), .A2(n442), .ZN(n441) );
  INV_X1 U538 ( .A(n738), .ZN(n446) );
  NOR2_X1 U539 ( .A1(n710), .A2(n722), .ZN(n711) );
  NOR2_X1 U540 ( .A1(n723), .A2(n722), .ZN(n724) );
  INV_X1 U541 ( .A(KEYINPUT84), .ZN(n637) );
  INV_X1 U542 ( .A(KEYINPUT30), .ZN(n463) );
  BUF_X1 U543 ( .A(n620), .Z(n624) );
  NOR2_X1 U544 ( .A1(n700), .A2(n722), .ZN(n702) );
  BUF_X1 U545 ( .A(n684), .Z(n686) );
  XNOR2_X2 U546 ( .A(G143), .B(KEYINPUT64), .ZN(n449) );
  XNOR2_X2 U547 ( .A(n449), .B(G128), .ZN(n531) );
  XNOR2_X2 U548 ( .A(n531), .B(n450), .ZN(n514) );
  XNOR2_X1 U549 ( .A(n451), .B(G134), .ZN(n452) );
  XNOR2_X2 U550 ( .A(n514), .B(n452), .ZN(n768) );
  XNOR2_X2 U551 ( .A(n768), .B(G146), .ZN(n469) );
  XOR2_X1 U552 ( .A(KEYINPUT5), .B(KEYINPUT98), .Z(n454) );
  NAND2_X1 U553 ( .A1(n536), .A2(G210), .ZN(n453) );
  XNOR2_X1 U554 ( .A(n454), .B(n453), .ZN(n458) );
  XNOR2_X2 U555 ( .A(G113), .B(G101), .ZN(n457) );
  XOR2_X1 U556 ( .A(n458), .B(n506), .Z(n459) );
  XNOR2_X1 U557 ( .A(n461), .B(KEYINPUT76), .ZN(n518) );
  INV_X1 U558 ( .A(G214), .ZN(n462) );
  OR2_X1 U559 ( .A1(n518), .A2(n462), .ZN(n642) );
  XNOR2_X1 U560 ( .A(n464), .B(n463), .ZN(n503) );
  NAND2_X1 U561 ( .A1(G227), .A2(n769), .ZN(n465) );
  XNOR2_X1 U562 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U563 ( .A(n507), .B(n467), .ZN(n468) );
  XNOR2_X1 U564 ( .A(n469), .B(n468), .ZN(n713) );
  NOR2_X2 U565 ( .A1(G902), .A2(n713), .ZN(n471) );
  XNOR2_X2 U566 ( .A(n471), .B(n470), .ZN(n559) );
  XOR2_X1 U567 ( .A(KEYINPUT24), .B(KEYINPUT86), .Z(n473) );
  XNOR2_X1 U568 ( .A(G128), .B(G119), .ZN(n472) );
  XNOR2_X1 U569 ( .A(n473), .B(n472), .ZN(n475) );
  XOR2_X1 U570 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n474) );
  XNOR2_X1 U571 ( .A(n476), .B(n509), .ZN(n767) );
  XNOR2_X1 U572 ( .A(n477), .B(n767), .ZN(n484) );
  NAND2_X1 U573 ( .A1(G234), .A2(n769), .ZN(n478) );
  XOR2_X1 U574 ( .A(KEYINPUT8), .B(n478), .Z(n529) );
  NAND2_X1 U575 ( .A1(n529), .A2(G221), .ZN(n480) );
  XNOR2_X1 U576 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U577 ( .A(n484), .B(n483), .ZN(n704) );
  INV_X1 U578 ( .A(G902), .ZN(n534) );
  NAND2_X1 U579 ( .A1(n704), .A2(n534), .ZN(n491) );
  XOR2_X1 U580 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n487) );
  XNOR2_X1 U581 ( .A(KEYINPUT15), .B(G902), .ZN(n687) );
  NAND2_X1 U582 ( .A1(n687), .A2(G234), .ZN(n485) );
  XNOR2_X1 U583 ( .A(n485), .B(KEYINPUT20), .ZN(n492) );
  NAND2_X1 U584 ( .A1(n492), .A2(G217), .ZN(n486) );
  XNOR2_X1 U585 ( .A(n487), .B(n486), .ZN(n489) );
  INV_X1 U586 ( .A(KEYINPUT96), .ZN(n488) );
  XNOR2_X1 U587 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X2 U588 ( .A(n491), .B(n490), .ZN(n552) );
  NAND2_X1 U589 ( .A1(G221), .A2(n492), .ZN(n493) );
  XNOR2_X1 U590 ( .A(KEYINPUT21), .B(n493), .ZN(n653) );
  XOR2_X1 U591 ( .A(n653), .B(KEYINPUT97), .Z(n595) );
  XNOR2_X1 U592 ( .A(n495), .B(n494), .ZN(n496) );
  AND2_X1 U593 ( .A1(n496), .A2(G952), .ZN(n671) );
  AND2_X1 U594 ( .A1(n671), .A2(n769), .ZN(n587) );
  NAND2_X1 U595 ( .A1(G902), .A2(n496), .ZN(n588) );
  OR2_X1 U596 ( .A1(n769), .A2(n588), .ZN(n497) );
  NOR2_X1 U597 ( .A1(G900), .A2(n497), .ZN(n498) );
  NOR2_X1 U598 ( .A1(n587), .A2(n498), .ZN(n499) );
  XOR2_X1 U599 ( .A(KEYINPUT83), .B(n499), .Z(n550) );
  INV_X1 U600 ( .A(n550), .ZN(n500) );
  NAND2_X1 U601 ( .A1(n503), .A2(n502), .ZN(n576) );
  XNOR2_X1 U602 ( .A(n504), .B(KEYINPUT73), .ZN(n505) );
  XNOR2_X1 U603 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n508) );
  XNOR2_X1 U604 ( .A(n509), .B(n508), .ZN(n512) );
  NAND2_X1 U605 ( .A1(n769), .A2(G224), .ZN(n510) );
  XNOR2_X1 U606 ( .A(n510), .B(KEYINPUT79), .ZN(n511) );
  XNOR2_X1 U607 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U608 ( .A(n514), .B(n513), .ZN(n515) );
  INV_X1 U609 ( .A(n687), .ZN(n688) );
  INV_X1 U610 ( .A(G210), .ZN(n517) );
  OR2_X1 U611 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U612 ( .A(n519), .B(KEYINPUT82), .ZN(n520) );
  XNOR2_X1 U613 ( .A(KEYINPUT90), .B(KEYINPUT39), .ZN(n521) );
  XNOR2_X1 U614 ( .A(n522), .B(n521), .ZN(n580) );
  XOR2_X1 U615 ( .A(G134), .B(G122), .Z(n524) );
  XNOR2_X1 U616 ( .A(n524), .B(n523), .ZN(n528) );
  XOR2_X1 U617 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n526) );
  XNOR2_X1 U618 ( .A(KEYINPUT9), .B(KEYINPUT102), .ZN(n525) );
  XNOR2_X1 U619 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U620 ( .A(n528), .B(n527), .Z(n533) );
  AND2_X1 U621 ( .A1(G217), .A2(n529), .ZN(n530) );
  XNOR2_X1 U622 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U623 ( .A(n533), .B(n532), .ZN(n692) );
  NAND2_X1 U624 ( .A1(n692), .A2(n534), .ZN(n535) );
  XNOR2_X1 U625 ( .A(n535), .B(G478), .ZN(n577) );
  NAND2_X1 U626 ( .A1(n536), .A2(G214), .ZN(n537) );
  XNOR2_X1 U627 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U628 ( .A(KEYINPUT11), .B(n539), .ZN(n540) );
  XNOR2_X1 U629 ( .A(n540), .B(n767), .ZN(n546) );
  XNOR2_X1 U630 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U631 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U632 ( .A(n546), .B(n545), .ZN(n707) );
  NOR2_X1 U633 ( .A1(G902), .A2(n707), .ZN(n548) );
  XNOR2_X1 U634 ( .A(KEYINPUT13), .B(G475), .ZN(n547) );
  XNOR2_X1 U635 ( .A(n548), .B(n547), .ZN(n578) );
  XOR2_X1 U636 ( .A(n578), .B(KEYINPUT100), .Z(n569) );
  NOR2_X1 U637 ( .A1(n577), .A2(n569), .ZN(n740) );
  INV_X1 U638 ( .A(n740), .ZN(n744) );
  NOR2_X1 U639 ( .A1(n653), .A2(n550), .ZN(n551) );
  XNOR2_X1 U640 ( .A(KEYINPUT68), .B(n551), .ZN(n553) );
  NAND2_X1 U641 ( .A1(n553), .A2(n552), .ZN(n561) );
  INV_X1 U642 ( .A(n556), .ZN(n643) );
  NAND2_X1 U643 ( .A1(n643), .A2(n642), .ZN(n647) );
  OR2_X1 U644 ( .A1(n577), .A2(n578), .ZN(n645) );
  NOR2_X1 U645 ( .A1(n647), .A2(n645), .ZN(n558) );
  XNOR2_X1 U646 ( .A(KEYINPUT108), .B(KEYINPUT41), .ZN(n557) );
  XNOR2_X2 U647 ( .A(n558), .B(n557), .ZN(n674) );
  XNOR2_X1 U648 ( .A(n559), .B(KEYINPUT1), .ZN(n610) );
  INV_X1 U649 ( .A(n610), .ZN(n581) );
  INV_X1 U650 ( .A(n620), .ZN(n656) );
  NAND2_X1 U651 ( .A1(n616), .A2(n642), .ZN(n560) );
  INV_X1 U652 ( .A(n642), .ZN(n564) );
  INV_X1 U653 ( .A(KEYINPUT65), .ZN(n566) );
  XNOR2_X1 U654 ( .A(n566), .B(KEYINPUT19), .ZN(n567) );
  NAND2_X1 U655 ( .A1(n577), .A2(n569), .ZN(n748) );
  INV_X1 U656 ( .A(n748), .ZN(n733) );
  OR2_X1 U657 ( .A1(n740), .A2(n733), .ZN(n646) );
  INV_X1 U658 ( .A(KEYINPUT75), .ZN(n570) );
  NAND2_X1 U659 ( .A1(n571), .A2(KEYINPUT47), .ZN(n575) );
  XNOR2_X1 U660 ( .A(KEYINPUT75), .B(n646), .ZN(n572) );
  NOR2_X1 U661 ( .A1(KEYINPUT47), .A2(n572), .ZN(n573) );
  NAND2_X1 U662 ( .A1(n355), .A2(n573), .ZN(n574) );
  NAND2_X1 U663 ( .A1(n578), .A2(n577), .ZN(n614) );
  OR2_X1 U664 ( .A1(n614), .A2(n565), .ZN(n579) );
  NOR2_X1 U665 ( .A1(n576), .A2(n579), .ZN(n738) );
  NOR2_X1 U666 ( .A1(n580), .A2(n748), .ZN(n752) );
  XOR2_X1 U667 ( .A(KEYINPUT43), .B(KEYINPUT105), .Z(n584) );
  INV_X1 U668 ( .A(n581), .ZN(n658) );
  OR2_X1 U669 ( .A1(n582), .A2(n658), .ZN(n583) );
  XNOR2_X1 U670 ( .A(n584), .B(n583), .ZN(n585) );
  AND2_X1 U671 ( .A1(n585), .A2(n565), .ZN(n681) );
  NOR2_X1 U672 ( .A1(n752), .A2(n681), .ZN(n586) );
  INV_X1 U673 ( .A(n587), .ZN(n590) );
  INV_X1 U674 ( .A(G898), .ZN(n757) );
  NAND2_X1 U675 ( .A1(G953), .A2(n757), .ZN(n762) );
  OR2_X1 U676 ( .A1(n762), .A2(n588), .ZN(n589) );
  NAND2_X1 U677 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U678 ( .A1(n592), .A2(n591), .ZN(n594) );
  INV_X1 U679 ( .A(KEYINPUT0), .ZN(n593) );
  NOR2_X1 U680 ( .A1(n595), .A2(n645), .ZN(n597) );
  INV_X1 U681 ( .A(KEYINPUT103), .ZN(n596) );
  XNOR2_X1 U682 ( .A(n597), .B(n596), .ZN(n598) );
  NAND2_X1 U683 ( .A1(n626), .A2(n598), .ZN(n600) );
  INV_X1 U684 ( .A(KEYINPUT22), .ZN(n599) );
  NAND2_X1 U685 ( .A1(n658), .A2(n552), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n619), .A2(n353), .ZN(n603) );
  XNOR2_X1 U687 ( .A(KEYINPUT81), .B(KEYINPUT32), .ZN(n602) );
  XNOR2_X1 U688 ( .A(n603), .B(n602), .ZN(n683) );
  INV_X1 U689 ( .A(n619), .ZN(n608) );
  INV_X1 U690 ( .A(n552), .ZN(n604) );
  NOR2_X1 U691 ( .A1(n658), .A2(n604), .ZN(n606) );
  NAND2_X1 U692 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U693 ( .A1(n683), .A2(n609), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n610), .A2(n659), .ZN(n621) );
  INV_X1 U695 ( .A(KEYINPUT33), .ZN(n612) );
  INV_X1 U696 ( .A(n626), .ZN(n613) );
  NAND2_X1 U697 ( .A1(n615), .A2(n684), .ZN(n631) );
  OR2_X1 U698 ( .A1(n658), .A2(n552), .ZN(n617) );
  NOR2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n618) );
  AND2_X1 U700 ( .A1(n619), .A2(n618), .ZN(n725) );
  INV_X1 U701 ( .A(n725), .ZN(n629) );
  NOR2_X1 U702 ( .A1(n624), .A2(n621), .ZN(n664) );
  NAND2_X1 U703 ( .A1(n626), .A2(n664), .ZN(n623) );
  INV_X1 U704 ( .A(KEYINPUT31), .ZN(n622) );
  AND2_X1 U705 ( .A1(n448), .A2(n624), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n727) );
  NAND2_X1 U707 ( .A1(n747), .A2(n727), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n627), .A2(n646), .ZN(n628) );
  INV_X1 U709 ( .A(n631), .ZN(n633) );
  INV_X1 U710 ( .A(KEYINPUT44), .ZN(n632) );
  INV_X1 U711 ( .A(KEYINPUT88), .ZN(n634) );
  XNOR2_X1 U712 ( .A(n634), .B(KEYINPUT45), .ZN(n635) );
  XNOR2_X1 U713 ( .A(KEYINPUT2), .B(KEYINPUT85), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n640), .A2(n636), .ZN(n638) );
  XNOR2_X1 U715 ( .A(n638), .B(n637), .ZN(n641) );
  INV_X1 U716 ( .A(KEYINPUT2), .ZN(n639) );
  NOR2_X1 U717 ( .A1(n641), .A2(n689), .ZN(n679) );
  NOR2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n650) );
  INV_X1 U720 ( .A(n646), .ZN(n648) );
  NOR2_X1 U721 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U723 ( .A(KEYINPUT119), .B(n651), .Z(n652) );
  NOR2_X1 U724 ( .A1(n673), .A2(n652), .ZN(n668) );
  NAND2_X1 U725 ( .A1(n552), .A2(n653), .ZN(n654) );
  XNOR2_X1 U726 ( .A(KEYINPUT49), .B(n654), .ZN(n655) );
  NOR2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U728 ( .A(KEYINPUT118), .B(n657), .Z(n662) );
  NOR2_X1 U729 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U730 ( .A(KEYINPUT50), .B(n660), .ZN(n661) );
  NOR2_X1 U731 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U733 ( .A(KEYINPUT51), .B(n665), .Z(n666) );
  NOR2_X1 U734 ( .A1(n674), .A2(n666), .ZN(n667) );
  NOR2_X1 U735 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U736 ( .A(KEYINPUT52), .B(n669), .Z(n670) );
  XNOR2_X1 U737 ( .A(n670), .B(KEYINPUT120), .ZN(n672) );
  NAND2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n677) );
  NOR2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U740 ( .A(n675), .B(KEYINPUT121), .ZN(n676) );
  NAND2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U743 ( .A(n681), .B(G140), .Z(G42) );
  XNOR2_X1 U744 ( .A(G119), .B(KEYINPUT127), .ZN(n682) );
  XNOR2_X1 U745 ( .A(n683), .B(n682), .ZN(G21) );
  XNOR2_X1 U746 ( .A(G122), .B(KEYINPUT126), .ZN(n685) );
  XNOR2_X1 U747 ( .A(n686), .B(n685), .ZN(G24) );
  NOR2_X2 U748 ( .A1(n690), .A2(n689), .ZN(n695) );
  NAND2_X1 U749 ( .A1(n695), .A2(G478), .ZN(n691) );
  XOR2_X1 U750 ( .A(n692), .B(n691), .Z(n693) );
  XNOR2_X1 U751 ( .A(n694), .B(KEYINPUT124), .ZN(G63) );
  BUF_X2 U752 ( .A(n695), .Z(n717) );
  NAND2_X1 U753 ( .A1(n717), .A2(G472), .ZN(n699) );
  XOR2_X1 U754 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n696) );
  XNOR2_X1 U755 ( .A(n697), .B(n696), .ZN(n698) );
  XNOR2_X1 U756 ( .A(n699), .B(n698), .ZN(n700) );
  XOR2_X1 U757 ( .A(KEYINPUT92), .B(KEYINPUT63), .Z(n701) );
  XNOR2_X1 U758 ( .A(n702), .B(n701), .ZN(G57) );
  NAND2_X1 U759 ( .A1(n717), .A2(G217), .ZN(n703) );
  XOR2_X1 U760 ( .A(n704), .B(n703), .Z(n705) );
  NOR2_X1 U761 ( .A1(n705), .A2(n722), .ZN(G66) );
  NAND2_X1 U762 ( .A1(n717), .A2(G475), .ZN(n709) );
  XNOR2_X1 U763 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n706) );
  XNOR2_X1 U764 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U765 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U766 ( .A(n711), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U767 ( .A1(n717), .A2(G469), .ZN(n715) );
  XOR2_X1 U768 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n712) );
  XNOR2_X1 U769 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U770 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U771 ( .A1(n716), .A2(n722), .ZN(G54) );
  NAND2_X1 U772 ( .A1(n717), .A2(G210), .ZN(n721) );
  XOR2_X1 U773 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n718) );
  XNOR2_X1 U774 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U775 ( .A(n721), .B(n720), .ZN(n723) );
  XNOR2_X1 U776 ( .A(n724), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U777 ( .A(G101), .B(n725), .Z(G3) );
  NOR2_X1 U778 ( .A1(n744), .A2(n727), .ZN(n726) );
  XOR2_X1 U779 ( .A(G104), .B(n726), .Z(G6) );
  NOR2_X1 U780 ( .A1(n748), .A2(n727), .ZN(n732) );
  XOR2_X1 U781 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n729) );
  XNOR2_X1 U782 ( .A(G107), .B(KEYINPUT26), .ZN(n728) );
  XNOR2_X1 U783 ( .A(n729), .B(n728), .ZN(n730) );
  XNOR2_X1 U784 ( .A(KEYINPUT110), .B(n730), .ZN(n731) );
  XNOR2_X1 U785 ( .A(n732), .B(n731), .ZN(G9) );
  XOR2_X1 U786 ( .A(G128), .B(KEYINPUT112), .Z(n735) );
  NAND2_X1 U787 ( .A1(n355), .A2(n733), .ZN(n734) );
  XNOR2_X1 U788 ( .A(n735), .B(n734), .ZN(n737) );
  XOR2_X1 U789 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n736) );
  XNOR2_X1 U790 ( .A(n737), .B(n736), .ZN(G30) );
  XOR2_X1 U791 ( .A(n738), .B(G143), .Z(n739) );
  XNOR2_X1 U792 ( .A(KEYINPUT114), .B(n739), .ZN(G45) );
  XOR2_X1 U793 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n742) );
  NAND2_X1 U794 ( .A1(n355), .A2(n740), .ZN(n741) );
  XNOR2_X1 U795 ( .A(n742), .B(n741), .ZN(n743) );
  XNOR2_X1 U796 ( .A(G146), .B(n743), .ZN(G48) );
  NOR2_X1 U797 ( .A1(n744), .A2(n747), .ZN(n746) );
  XNOR2_X1 U798 ( .A(G113), .B(KEYINPUT117), .ZN(n745) );
  XNOR2_X1 U799 ( .A(n746), .B(n745), .ZN(G15) );
  NOR2_X1 U800 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U801 ( .A(G116), .B(n749), .Z(G18) );
  XNOR2_X1 U802 ( .A(G125), .B(n750), .ZN(n751) );
  XNOR2_X1 U803 ( .A(n751), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U804 ( .A(G134), .B(n752), .Z(G36) );
  BUF_X1 U805 ( .A(n753), .Z(n754) );
  NOR2_X1 U806 ( .A1(n754), .A2(G953), .ZN(n759) );
  NAND2_X1 U807 ( .A1(G953), .A2(G224), .ZN(n755) );
  XOR2_X1 U808 ( .A(KEYINPUT61), .B(n755), .Z(n756) );
  NOR2_X1 U809 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U810 ( .A1(n759), .A2(n758), .ZN(n766) );
  XNOR2_X1 U811 ( .A(n761), .B(n760), .ZN(n763) );
  NAND2_X1 U812 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U813 ( .A(KEYINPUT125), .B(n764), .Z(n765) );
  XNOR2_X1 U814 ( .A(n766), .B(n765), .ZN(G69) );
  XOR2_X1 U815 ( .A(n768), .B(n767), .Z(n771) );
  NAND2_X1 U816 ( .A1(n770), .A2(n769), .ZN(n775) );
  XNOR2_X1 U817 ( .A(G227), .B(n771), .ZN(n772) );
  NAND2_X1 U818 ( .A1(n772), .A2(G900), .ZN(n773) );
  NAND2_X1 U819 ( .A1(n773), .A2(G953), .ZN(n774) );
  NAND2_X1 U820 ( .A1(n775), .A2(n774), .ZN(G72) );
  XOR2_X1 U821 ( .A(n776), .B(G131), .Z(G33) );
  XOR2_X1 U822 ( .A(n777), .B(G137), .Z(G39) );
endmodule

