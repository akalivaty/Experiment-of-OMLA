//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1269, new_n1270, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1331, new_n1332;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  OR3_X1    g0010(.A1(new_n210), .A2(KEYINPUT64), .A3(G13), .ZN(new_n211));
  OAI21_X1  g0011(.A(KEYINPUT64), .B1(new_n210), .B2(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G264), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n209), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(G50), .B1(G58), .B2(G68), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(new_n217), .A2(KEYINPUT0), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n223), .B1(KEYINPUT0), .B2(new_n217), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n206), .C2(new_n216), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n229), .B1(new_n202), .B2(new_n230), .C1(new_n205), .C2(new_n215), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n210), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT1), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n224), .A2(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n230), .ZN(new_n236));
  XOR2_X1   g0036(.A(KEYINPUT2), .B(G226), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT68), .ZN(new_n250));
  OAI21_X1  g0050(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n219), .A2(G33), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n251), .B1(new_n252), .B2(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n218), .ZN(new_n259));
  INV_X1    g0059(.A(G13), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n260), .A2(new_n219), .A3(G1), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n257), .A2(new_n259), .B1(new_n201), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT9), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n261), .A2(new_n259), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT65), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n261), .A2(new_n259), .A3(KEYINPUT65), .ZN(new_n269));
  OAI211_X1 g0069(.A(G50), .B(new_n265), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n262), .A2(new_n263), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n263), .B1(new_n262), .B2(new_n270), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n279), .A3(G274), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n281), .B1(G226), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n287), .A2(new_n289), .A3(G222), .A4(new_n290), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n287), .A2(new_n289), .A3(G223), .A4(G1698), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT3), .B(G33), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n291), .B(new_n292), .C1(new_n226), .C2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n279), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n285), .A2(new_n296), .A3(G190), .ZN(new_n297));
  INV_X1    g0097(.A(G200), .ZN(new_n298));
  INV_X1    g0098(.A(G226), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n280), .B1(new_n299), .B2(new_n283), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(new_n295), .B2(new_n294), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n297), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n250), .B(KEYINPUT10), .C1(new_n274), .C2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n262), .A2(new_n270), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT9), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n302), .B1(new_n305), .B2(new_n271), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT68), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT67), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n272), .B2(new_n273), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n305), .A2(KEYINPUT67), .A3(new_n271), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n303), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n219), .A2(G33), .A3(G77), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n315), .B1(new_n219), .B2(G68), .C1(new_n254), .C2(new_n201), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n259), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT11), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(KEYINPUT69), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT69), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n316), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT11), .B1(new_n316), .B2(new_n259), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G68), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n261), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT12), .ZN(new_n328));
  INV_X1    g0128(.A(new_n259), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n260), .A2(G1), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G20), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n331), .A3(KEYINPUT66), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT66), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n261), .B2(new_n259), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(G68), .A3(new_n265), .ZN(new_n336));
  AND4_X1   g0136(.A1(new_n321), .A2(new_n325), .A3(new_n328), .A4(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G169), .ZN(new_n338));
  OR2_X1    g0138(.A1(new_n338), .A2(KEYINPUT70), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n293), .A2(G232), .A3(G1698), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n293), .A2(G226), .A3(new_n290), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n295), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n281), .B1(G238), .B2(new_n284), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n340), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(new_n346), .A3(new_n340), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n339), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n337), .B1(new_n350), .B2(KEYINPUT14), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n348), .A2(G179), .A3(new_n349), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT14), .ZN(new_n353));
  INV_X1    g0153(.A(new_n349), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(new_n347), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n352), .B(new_n353), .C1(new_n355), .C2(new_n339), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n325), .A2(new_n321), .A3(new_n328), .A4(new_n336), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n355), .B2(G190), .ZN(new_n358));
  OAI21_X1  g0158(.A(G200), .B1(new_n354), .B2(new_n347), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n351), .A2(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G179), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n301), .A2(new_n361), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n304), .B(new_n362), .C1(G169), .C2(new_n301), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n335), .A2(G77), .A3(new_n265), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G20), .A2(G77), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT15), .B(G87), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n365), .B1(new_n255), .B2(new_n254), .C1(new_n256), .C2(new_n366), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n259), .B1(new_n226), .B2(new_n261), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n293), .A2(G238), .A3(G1698), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n293), .A2(G232), .A3(new_n290), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n370), .B(new_n371), .C1(new_n206), .C2(new_n293), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n295), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n281), .B1(G244), .B2(new_n284), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n369), .B1(new_n376), .B2(G190), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n298), .B2(new_n376), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n361), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n375), .A2(new_n338), .B1(new_n364), .B2(new_n368), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n314), .A2(new_n360), .A3(new_n363), .A4(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n255), .B1(new_n264), .B2(G20), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n268), .B2(new_n269), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n255), .A2(new_n261), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AND2_X1   g0187(.A1(G58), .A2(G68), .ZN(new_n388));
  NOR2_X1   g0188(.A1(G58), .A2(G68), .ZN(new_n389));
  OAI21_X1  g0189(.A(G20), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n253), .A2(KEYINPUT72), .A3(G159), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT72), .B1(new_n253), .B2(G159), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(G20), .B1(new_n287), .B2(new_n289), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n326), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT7), .B1(new_n293), .B2(G20), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n329), .B1(new_n398), .B2(KEYINPUT16), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT16), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n219), .A2(KEYINPUT7), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n288), .A2(KEYINPUT73), .A3(G33), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n287), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT73), .B1(new_n288), .B2(G33), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n395), .B1(new_n293), .B2(G20), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n326), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n400), .B1(new_n407), .B2(new_n393), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n387), .B1(new_n399), .B2(new_n408), .ZN(new_n409));
  OR2_X1    g0209(.A1(G223), .A2(G1698), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n299), .A2(G1698), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n287), .A2(new_n410), .A3(new_n289), .A4(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n295), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n279), .A2(G232), .A3(new_n282), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n280), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n298), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n279), .B1(new_n412), .B2(new_n413), .ZN(new_n420));
  INV_X1    g0220(.A(G190), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n420), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT74), .B1(new_n409), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n396), .A2(new_n397), .ZN(new_n425));
  INV_X1    g0225(.A(new_n393), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT16), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n408), .A2(new_n259), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n387), .ZN(new_n429));
  AND4_X1   g0229(.A1(KEYINPUT74), .A2(new_n428), .A3(new_n429), .A4(new_n423), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT17), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n429), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n420), .A2(new_n417), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n434), .A2(new_n338), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n420), .A2(new_n417), .A3(new_n361), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n432), .B1(new_n433), .B2(new_n438), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n409), .A2(KEYINPUT18), .A3(new_n437), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT17), .B1(new_n409), .B2(new_n423), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n431), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(G20), .B1(G33), .B2(G283), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT75), .B(G97), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n445), .B1(new_n446), .B2(G33), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT84), .ZN(new_n448));
  INV_X1    g0248(.A(G116), .ZN(new_n449));
  AOI221_X4 g0249(.A(new_n448), .B1(new_n449), .B2(G20), .C1(new_n258), .C2(new_n218), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(G20), .ZN(new_n451));
  AOI21_X1  g0251(.A(KEYINPUT84), .B1(new_n259), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n447), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT20), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n447), .B(KEYINPUT20), .C1(new_n450), .C2(new_n452), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT76), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n286), .B2(G1), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n264), .A2(KEYINPUT76), .A3(G33), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n332), .A2(new_n334), .A3(G116), .A4(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT83), .B1(new_n331), .B2(G116), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT83), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n261), .A2(new_n464), .A3(new_n449), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n457), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n287), .A2(new_n289), .A3(G264), .A4(G1698), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n287), .A2(new_n289), .A3(G257), .A4(new_n290), .ZN(new_n470));
  INV_X1    g0270(.A(G303), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n469), .B(new_n470), .C1(new_n471), .C2(new_n293), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n295), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n275), .A2(KEYINPUT5), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n264), .B(G45), .C1(new_n275), .C2(KEYINPUT5), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT78), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n276), .A2(G1), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT5), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G41), .ZN(new_n480));
  AOI21_X1  g0280(.A(KEYINPUT78), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(G270), .B(new_n279), .C1(new_n477), .C2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n481), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(KEYINPUT78), .A3(new_n480), .ZN(new_n484));
  INV_X1    g0284(.A(G274), .ZN(new_n485));
  INV_X1    g0285(.A(new_n218), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(new_n278), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n483), .A2(new_n484), .A3(new_n487), .A4(new_n474), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n473), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT82), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n473), .A2(new_n482), .A3(KEYINPUT82), .A4(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n468), .B1(new_n493), .B2(G200), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(new_n421), .B2(new_n493), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n338), .B1(new_n457), .B2(new_n467), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n493), .A2(new_n496), .A3(KEYINPUT21), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n489), .A2(new_n361), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n468), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT21), .B1(new_n493), .B2(new_n496), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT85), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI211_X1 g0303(.A(KEYINPUT85), .B(KEYINPUT21), .C1(new_n493), .C2(new_n496), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n495), .B(new_n500), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n287), .A2(new_n289), .A3(G244), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G283), .ZN(new_n509));
  AND2_X1   g0309(.A1(KEYINPUT4), .A2(G244), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n287), .A2(new_n289), .A3(new_n510), .A4(new_n290), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n287), .A2(new_n289), .A3(G250), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n290), .B1(new_n513), .B2(KEYINPUT4), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n295), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT77), .ZN(new_n516));
  OAI211_X1 g0316(.A(G257), .B(new_n279), .C1(new_n477), .C2(new_n481), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n488), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT77), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n520), .B(new_n295), .C1(new_n512), .C2(new_n514), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n516), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G200), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n515), .A2(G190), .A3(new_n488), .A4(new_n517), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n446), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G97), .A2(G107), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT6), .B1(new_n207), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(G20), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n253), .A2(G77), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n206), .B1(new_n405), .B2(new_n406), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n259), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n266), .A2(new_n461), .ZN(new_n534));
  MUX2_X1   g0334(.A(new_n331), .B(new_n534), .S(G97), .Z(new_n535));
  AND3_X1   g0335(.A1(new_n524), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n519), .A2(new_n515), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n537), .A2(new_n338), .B1(new_n533), .B2(new_n535), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n517), .A2(new_n488), .A3(new_n361), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n516), .A2(new_n521), .A3(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n523), .A2(new_n536), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n266), .A2(G87), .A3(new_n461), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT81), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n266), .A2(KEYINPUT81), .A3(G87), .A4(new_n461), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT19), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(new_n446), .B2(new_n256), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n205), .A2(KEYINPUT75), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT75), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G97), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G87), .A2(G107), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n219), .B1(new_n343), .B2(new_n547), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n293), .A2(new_n219), .A3(G68), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n548), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(new_n259), .B1(new_n261), .B2(new_n366), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n546), .A2(new_n558), .ZN(new_n559));
  OR2_X1    g0359(.A1(G238), .A2(G1698), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n227), .A2(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n287), .A2(new_n560), .A3(new_n289), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G116), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n279), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n478), .A2(new_n485), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n209), .B1(new_n276), .B2(G1), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n279), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT79), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT79), .ZN(new_n570));
  INV_X1    g0370(.A(new_n563), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G238), .A2(G1698), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n227), .B2(G1698), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n571), .B1(new_n573), .B2(new_n293), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n570), .B(new_n567), .C1(new_n574), .C2(new_n279), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n569), .A2(new_n575), .A3(G190), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n569), .A2(new_n575), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n559), .B(new_n576), .C1(new_n298), .C2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n569), .A2(new_n575), .A3(new_n361), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT80), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n577), .A2(new_n338), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n569), .A2(new_n575), .A3(KEYINPUT80), .A4(new_n361), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n557), .A2(new_n259), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n366), .A2(new_n261), .ZN(new_n586));
  INV_X1    g0386(.A(new_n366), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n266), .A2(new_n587), .A3(new_n461), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n582), .A2(new_n583), .A3(new_n584), .A4(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n579), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(G264), .B(new_n279), .C1(new_n477), .C2(new_n481), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n287), .A2(new_n289), .A3(G257), .A4(G1698), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n287), .A2(new_n289), .A3(G250), .A4(new_n290), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT88), .ZN(new_n596));
  AND2_X1   g0396(.A1(KEYINPUT87), .A2(G294), .ZN(new_n597));
  NOR2_X1   g0397(.A1(KEYINPUT87), .A2(G294), .ZN(new_n598));
  OAI21_X1  g0398(.A(G33), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n594), .A2(new_n595), .A3(new_n596), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n279), .B1(new_n601), .B2(KEYINPUT88), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n593), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(G179), .A3(new_n488), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n601), .A2(KEYINPUT88), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n295), .A3(new_n600), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(new_n488), .A3(new_n592), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G169), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT23), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n219), .B2(G107), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n611), .A2(new_n612), .B1(new_n571), .B2(new_n219), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n287), .A2(new_n289), .A3(new_n219), .A4(G87), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT86), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT86), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n293), .A2(new_n616), .A3(new_n219), .A4(G87), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT22), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n615), .B2(new_n617), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n613), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT24), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT24), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n623), .B(new_n613), .C1(new_n619), .C2(new_n620), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n329), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n331), .A2(G107), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n626), .B(KEYINPUT25), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n266), .A2(G107), .A3(new_n461), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n609), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n615), .A2(new_n617), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT22), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n615), .A2(new_n617), .A3(new_n618), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n623), .B1(new_n634), .B2(new_n613), .ZN(new_n635));
  INV_X1    g0435(.A(new_n624), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n259), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n607), .A2(new_n298), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n606), .A2(new_n421), .A3(new_n488), .A4(new_n592), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n629), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n541), .A2(new_n591), .A3(new_n630), .A4(new_n642), .ZN(new_n643));
  NOR4_X1   g0443(.A1(new_n383), .A2(new_n444), .A3(new_n505), .A4(new_n643), .ZN(G372));
  NOR2_X1   g0444(.A1(new_n383), .A2(new_n444), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n536), .A2(new_n523), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n533), .A2(new_n535), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n648));
  INV_X1    g0448(.A(new_n514), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n279), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n338), .B1(new_n650), .B2(new_n518), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n540), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(G200), .B1(new_n564), .B2(new_n568), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n576), .A2(new_n558), .A3(new_n546), .A4(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n338), .B1(new_n564), .B2(new_n568), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n580), .A2(new_n589), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n646), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n637), .A2(new_n640), .A3(new_n641), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT89), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n500), .B(new_n630), .C1(new_n503), .C2(new_n504), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n540), .A2(new_n647), .A3(new_n651), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n654), .A2(new_n656), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT89), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(new_n642), .A4(new_n646), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n660), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n591), .B2(new_n662), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n657), .A2(new_n662), .A3(new_n668), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n656), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n645), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT90), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT17), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n428), .A2(new_n429), .A3(new_n423), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT74), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n409), .A2(KEYINPUT74), .A3(new_n423), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n358), .A2(new_n359), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(new_n379), .A3(new_n380), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n351), .A2(new_n356), .ZN(new_n684));
  AOI211_X1 g0484(.A(new_n442), .B(new_n681), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n441), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n314), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n687), .A2(new_n363), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n675), .A2(new_n688), .ZN(G369));
  NAND2_X1  g0489(.A1(new_n497), .A2(new_n499), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n493), .A2(new_n496), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT85), .B1(new_n691), .B2(KEYINPUT21), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n501), .A2(new_n502), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n330), .A2(new_n219), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(new_n697), .A3(G213), .ZN(new_n698));
  INV_X1    g0498(.A(G343), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n468), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n694), .A2(new_n495), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n694), .B2(new_n701), .ZN(new_n703));
  AND3_X1   g0503(.A1(new_n703), .A2(KEYINPUT91), .A3(G330), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT91), .B1(new_n703), .B2(G330), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n630), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n700), .ZN(new_n709));
  XOR2_X1   g0509(.A(new_n709), .B(KEYINPUT92), .Z(new_n710));
  OAI21_X1  g0510(.A(new_n700), .B1(new_n625), .B2(new_n629), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n630), .A2(new_n642), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n694), .A2(new_n700), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n700), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n708), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n714), .A2(new_n716), .A3(new_n718), .ZN(G399));
  NOR2_X1   g0519(.A1(new_n214), .A2(G41), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n553), .A2(G116), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR3_X1   g0522(.A1(new_n720), .A2(new_n264), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(new_n222), .B2(new_n720), .ZN(new_n724));
  XOR2_X1   g0524(.A(new_n724), .B(KEYINPUT28), .Z(new_n725));
  AOI211_X1 g0525(.A(KEYINPUT29), .B(new_n700), .C1(new_n667), .C2(new_n672), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n662), .A2(new_n668), .A3(new_n590), .A4(new_n579), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT26), .B1(new_n663), .B2(new_n652), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n656), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n658), .A2(new_n659), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n661), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n700), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G330), .ZN(new_n735));
  AND4_X1   g0535(.A1(new_n630), .A2(new_n541), .A3(new_n591), .A4(new_n642), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n694), .A3(new_n495), .A4(new_n717), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n650), .A2(new_n518), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n738), .A2(new_n498), .A3(new_n578), .A4(new_n603), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n577), .A2(new_n489), .A3(new_n361), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(KEYINPUT30), .A3(new_n603), .A4(new_n738), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n564), .A2(new_n568), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G179), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n493), .A2(new_n522), .A3(new_n607), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n741), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(KEYINPUT31), .A3(new_n700), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT31), .B1(new_n747), .B2(new_n700), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n735), .B1(new_n737), .B2(new_n751), .ZN(new_n752));
  OR3_X1    g0552(.A1(new_n726), .A2(new_n734), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT93), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n725), .B1(new_n754), .B2(G1), .ZN(G364));
  INV_X1    g0555(.A(new_n720), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n260), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n264), .B1(new_n757), .B2(G45), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT94), .Z(new_n763));
  OR2_X1    g0563(.A1(new_n703), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n763), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n218), .B1(G20), .B2(new_n338), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT95), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n214), .A2(new_n293), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n222), .A2(new_n276), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n769), .B(new_n770), .C1(new_n276), .C2(new_n245), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n287), .A2(new_n289), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n214), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n773), .A2(G355), .B1(new_n449), .B2(new_n214), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n768), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n219), .B1(new_n776), .B2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n597), .A2(new_n598), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n219), .A2(new_n421), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n298), .A2(G179), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n293), .B(new_n779), .C1(G303), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n361), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n219), .A2(G190), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n781), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n787), .A2(G322), .B1(new_n790), .B2(G283), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n785), .A2(new_n788), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n788), .A2(new_n776), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G311), .A2(new_n793), .B1(new_n795), .B2(G329), .ZN(new_n796));
  NAND3_X1  g0596(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G190), .ZN(new_n798));
  XNOR2_X1  g0598(.A(KEYINPUT33), .B(G317), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n797), .A2(new_n421), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n798), .A2(new_n799), .B1(new_n800), .B2(G326), .ZN(new_n801));
  NAND4_X1  g0601(.A1(new_n784), .A2(new_n791), .A3(new_n796), .A4(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G58), .A2(new_n787), .B1(new_n793), .B2(G77), .ZN(new_n803));
  INV_X1    g0603(.A(new_n800), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n201), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT96), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n783), .A2(G87), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n293), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G107), .B2(new_n790), .ZN(new_n809));
  INV_X1    g0609(.A(new_n777), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n810), .A2(G97), .B1(G68), .B2(new_n798), .ZN(new_n811));
  INV_X1    g0611(.A(G159), .ZN(new_n812));
  OAI21_X1  g0612(.A(KEYINPUT32), .B1(new_n794), .B2(new_n812), .ZN(new_n813));
  OR3_X1    g0613(.A1(new_n794), .A2(KEYINPUT32), .A3(new_n812), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n809), .A2(new_n811), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n802), .B1(new_n806), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n775), .B1(new_n816), .B2(new_n766), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n759), .B1(new_n764), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n706), .B1(G330), .B2(new_n703), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n759), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT97), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  INV_X1    g0622(.A(new_n759), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n382), .A2(new_n717), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(new_n667), .B2(new_n672), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n700), .B1(new_n667), .B2(new_n672), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n381), .A2(new_n700), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n369), .A2(new_n700), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n378), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n830), .B2(new_n381), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n826), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n752), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n823), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  INV_X1    g0635(.A(new_n766), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n761), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n823), .B1(G77), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT98), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n790), .A2(G87), .ZN(new_n840));
  INV_X1    g0640(.A(G294), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(new_n786), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n772), .B1(new_n777), .B2(new_n205), .C1(new_n206), .C2(new_n782), .ZN(new_n843));
  INV_X1    g0643(.A(new_n798), .ZN(new_n844));
  INV_X1    g0644(.A(G283), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n844), .A2(new_n845), .B1(new_n804), .B2(new_n471), .ZN(new_n846));
  INV_X1    g0646(.A(G311), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n792), .A2(new_n449), .B1(new_n794), .B2(new_n847), .ZN(new_n848));
  NOR4_X1   g0648(.A1(new_n842), .A2(new_n843), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT99), .B(G143), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n787), .A2(new_n850), .B1(new_n793), .B2(G159), .ZN(new_n851));
  INV_X1    g0651(.A(G137), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n851), .B1(new_n804), .B2(new_n852), .C1(new_n252), .C2(new_n844), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT34), .ZN(new_n854));
  INV_X1    g0654(.A(G132), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n293), .B1(new_n794), .B2(new_n855), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n782), .A2(new_n201), .B1(new_n789), .B2(new_n326), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n856), .B(new_n857), .C1(G58), .C2(new_n810), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n849), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n839), .B1(new_n836), .B2(new_n859), .C1(new_n831), .C2(new_n761), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n835), .A2(new_n860), .ZN(G384));
  NAND2_X1  g0661(.A1(new_n220), .A2(G116), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n526), .A2(new_n528), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n862), .B1(new_n863), .B2(KEYINPUT35), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(KEYINPUT35), .B2(new_n863), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT36), .ZN(new_n866));
  OAI21_X1  g0666(.A(G77), .B1(new_n202), .B2(new_n326), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n867), .A2(new_n221), .B1(G50), .B2(new_n326), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(G1), .A3(new_n260), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT100), .Z(new_n871));
  NAND2_X1  g0671(.A1(new_n684), .A2(new_n682), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n357), .A3(new_n700), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n360), .B1(new_n337), .B2(new_n717), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n828), .B(KEYINPUT101), .Z(new_n876));
  OAI21_X1  g0676(.A(new_n875), .B1(new_n825), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT102), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n427), .A2(new_n259), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n398), .A2(KEYINPUT16), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n429), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n698), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n679), .A2(new_n680), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n442), .B1(new_n886), .B2(KEYINPUT17), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n885), .B1(new_n887), .B2(new_n441), .ZN(new_n888));
  INV_X1    g0688(.A(new_n886), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n698), .B(KEYINPUT103), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n409), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n409), .A2(new_n437), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT37), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n883), .B1(new_n438), .B2(new_n884), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n679), .A3(new_n680), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n889), .A2(new_n894), .B1(new_n896), .B2(KEYINPUT37), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n880), .B1(new_n888), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n885), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n444), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n889), .A2(new_n894), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n900), .A2(new_n903), .A3(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n875), .B(KEYINPUT102), .C1(new_n825), .C2(new_n876), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n879), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n686), .A2(new_n891), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(KEYINPUT104), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT105), .B1(new_n681), .B2(new_n442), .ZN(new_n911));
  INV_X1    g0711(.A(new_n439), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n893), .A2(new_n432), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n912), .A2(new_n913), .A3(new_n892), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT105), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n431), .A2(new_n916), .A3(new_n443), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n911), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n677), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n919), .A2(new_n893), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n920), .A2(new_n892), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n910), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n901), .A2(new_n880), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n904), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n684), .A2(new_n700), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n898), .A2(new_n904), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT39), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n909), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT104), .B1(new_n907), .B2(new_n908), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n932), .A2(KEYINPUT106), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT106), .ZN(new_n935));
  INV_X1    g0735(.A(new_n924), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n914), .B1(new_n887), .B2(new_n916), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n921), .B1(new_n937), .B2(new_n911), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n936), .B1(new_n938), .B2(new_n910), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT39), .B1(new_n939), .B2(new_n904), .ZN(new_n940));
  INV_X1    g0740(.A(new_n928), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n905), .A2(new_n926), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n929), .B1(new_n877), .B2(new_n878), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n944), .A2(new_n906), .B1(new_n686), .B2(new_n891), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n943), .B1(new_n945), .B2(KEYINPUT104), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n907), .A2(new_n908), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT104), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n935), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n934), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n645), .B1(new_n734), .B2(new_n726), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n688), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n737), .A2(new_n751), .ZN(new_n955));
  INV_X1    g0755(.A(new_n831), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(new_n873), .B2(new_n874), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT40), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n958), .A2(new_n959), .A3(new_n905), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n955), .A2(new_n957), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n939), .B2(new_n904), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n960), .B1(new_n962), .B2(new_n959), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n955), .A2(new_n645), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n964), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(G330), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n954), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n264), .B2(new_n757), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n954), .A2(new_n967), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n871), .B1(new_n969), .B2(new_n970), .ZN(G367));
  NAND2_X1  g0771(.A1(new_n647), .A2(new_n700), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n541), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n662), .A2(new_n700), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n713), .A2(new_n715), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n652), .B1(new_n973), .B2(new_n630), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n976), .A2(KEYINPUT42), .B1(new_n717), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(KEYINPUT42), .B2(new_n976), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n559), .A2(new_n717), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n657), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n656), .B2(new_n980), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT107), .Z(new_n985));
  INV_X1    g0785(.A(new_n714), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n975), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n985), .B(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n720), .B(KEYINPUT41), .Z(new_n991));
  NAND2_X1  g0791(.A1(new_n716), .A2(new_n718), .ZN(new_n992));
  INV_X1    g0792(.A(new_n975), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT44), .Z(new_n995));
  NOR2_X1   g0795(.A1(new_n992), .A2(new_n993), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n986), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n713), .B(new_n715), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(new_n706), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n754), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n995), .A2(new_n714), .A3(new_n997), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n999), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n991), .B1(new_n1006), .B2(new_n754), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT108), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n758), .B(KEYINPUT109), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n990), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n982), .A2(new_n763), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n769), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(new_n241), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n767), .B1(new_n213), .B2(new_n366), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n293), .B1(new_n794), .B2(new_n852), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G159), .B2(new_n798), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n789), .A2(new_n226), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G50), .B2(new_n793), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G150), .A2(new_n787), .B1(new_n783), .B2(G58), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n810), .A2(G68), .B1(new_n800), .B2(new_n850), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n783), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1025), .B1(new_n206), .B2(new_n777), .C1(new_n844), .C2(new_n778), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT111), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n293), .B1(new_n795), .B2(G317), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n446), .B2(new_n789), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1026), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT46), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n782), .B2(new_n449), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT110), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT110), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n800), .A2(G311), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G303), .A2(new_n787), .B1(new_n793), .B2(G283), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1024), .B1(new_n1031), .B2(new_n1038), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT47), .Z(new_n1040));
  OAI221_X1 g0840(.A(new_n823), .B1(new_n1016), .B2(new_n1017), .C1(new_n1040), .C2(new_n836), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1014), .B1(new_n1041), .B2(KEYINPUT112), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(KEYINPUT112), .B2(new_n1041), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1013), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT113), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(G387));
  INV_X1    g0846(.A(new_n754), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n1001), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n1003), .A3(new_n720), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n710), .A2(new_n712), .A3(new_n765), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n773), .A2(new_n722), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(G107), .B2(new_n213), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n238), .A2(new_n276), .ZN(new_n1053));
  AOI211_X1 g0853(.A(G45), .B(new_n722), .C1(G68), .C2(G77), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n255), .A2(G50), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1015), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1052), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n823), .B1(new_n1058), .B2(new_n768), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n800), .A2(G159), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT114), .Z(new_n1061));
  OAI22_X1  g0861(.A1(new_n201), .A2(new_n786), .B1(new_n782), .B2(new_n226), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n789), .A2(new_n205), .B1(new_n794), .B2(new_n252), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n777), .A2(new_n366), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n293), .B1(new_n792), .B2(new_n326), .C1(new_n844), .C2(new_n255), .ZN(new_n1066));
  OR4_X1    g0866(.A1(new_n1061), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G317), .A2(new_n787), .B1(new_n793), .B2(G303), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n800), .A2(G322), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(new_n847), .C2(new_n844), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n782), .A2(new_n778), .B1(new_n777), .B2(new_n845), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n293), .B1(new_n795), .B2(G326), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n449), .C2(new_n789), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1067), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1059), .B1(new_n1080), .B2(new_n766), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1002), .A2(new_n1010), .B1(new_n1050), .B2(new_n1081), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1049), .A2(KEYINPUT116), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT116), .B1(new_n1049), .B2(new_n1082), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G393));
  NOR2_X1   g0886(.A1(new_n1015), .A2(new_n248), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n767), .B1(new_n213), .B2(new_n446), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n787), .A2(G311), .B1(G317), .B2(new_n800), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G283), .A2(new_n783), .B1(new_n795), .B2(G322), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1091), .A2(KEYINPUT117), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(KEYINPUT117), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n772), .B1(new_n789), .B2(new_n206), .ZN(new_n1094));
  NOR4_X1   g0894(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n792), .A2(new_n841), .B1(new_n777), .B2(new_n449), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G303), .B2(new_n798), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT118), .Z(new_n1098));
  OAI22_X1  g0898(.A1(new_n804), .A2(new_n252), .B1(new_n786), .B2(new_n812), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT51), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n782), .A2(new_n326), .B1(new_n792), .B2(new_n255), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n810), .A2(G77), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n798), .A2(G50), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n840), .A2(new_n1102), .A3(new_n293), .A4(new_n1103), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1101), .B(new_n1104), .C1(new_n795), .C2(new_n850), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1095), .A2(new_n1098), .B1(new_n1100), .B2(new_n1105), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n823), .B1(new_n1087), .B2(new_n1088), .C1(new_n1106), .C2(new_n836), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n993), .B2(new_n765), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n999), .A2(new_n1005), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n1010), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1004), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1006), .A2(new_n720), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(G390));
  NAND2_X1  g0913(.A1(new_n927), .A2(new_n930), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n877), .A2(new_n941), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n731), .A2(new_n700), .A3(new_n956), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT119), .B1(new_n1116), .B2(new_n876), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n661), .A2(new_n730), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n717), .B(new_n831), .C1(new_n1118), .C2(new_n729), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n876), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1117), .A2(new_n875), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n928), .B1(new_n939), .B2(new_n904), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1114), .A2(new_n1115), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n505), .A2(new_n643), .A3(new_n700), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n747), .A2(new_n700), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT31), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n748), .ZN(new_n1130));
  OAI211_X1 g0930(.A(G330), .B(new_n831), .C1(new_n1126), .C2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n875), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OR2_X1    g0934(.A1(new_n1125), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1115), .B1(new_n940), .B2(new_n942), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT120), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n752), .A2(KEYINPUT120), .A3(new_n831), .A4(new_n875), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1136), .A2(new_n1137), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n826), .A2(new_n1121), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n875), .B1(new_n752), .B2(new_n831), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1144), .B1(new_n1145), .B2(new_n1133), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1116), .A2(KEYINPUT119), .A3(new_n876), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1120), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1146), .B1(new_n1150), .B2(new_n1141), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n645), .B(G330), .C1(new_n1126), .C2(new_n1130), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(KEYINPUT121), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT121), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n752), .A2(new_n1154), .A3(new_n645), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1156), .A2(new_n688), .A3(new_n952), .ZN(new_n1157));
  AND3_X1   g0957(.A1(new_n1151), .A2(new_n1157), .A3(KEYINPUT122), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT122), .B1(new_n1151), .B2(new_n1157), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1135), .B(new_n1143), .C1(new_n1158), .C2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT122), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1143), .B1(new_n1125), .B2(new_n1134), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1151), .A2(new_n1157), .A3(KEYINPUT122), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1160), .A2(new_n720), .A3(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1164), .A2(new_n1011), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1114), .A2(new_n760), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n255), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n823), .B1(new_n1170), .B2(new_n837), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n782), .A2(new_n252), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1172), .B(KEYINPUT53), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G132), .A2(new_n787), .B1(new_n795), .B2(G125), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT54), .B(G143), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1173), .B(new_n1174), .C1(new_n792), .C2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n772), .B1(new_n790), .B2(G50), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n810), .A2(G159), .B1(G137), .B2(new_n798), .ZN(new_n1178));
  INV_X1    g0978(.A(G128), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1177), .B(new_n1178), .C1(new_n1179), .C2(new_n804), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G68), .A2(new_n790), .B1(new_n795), .B2(G294), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n449), .B2(new_n786), .C1(new_n446), .C2(new_n792), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G107), .A2(new_n798), .B1(new_n800), .B2(G283), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n807), .A2(new_n1183), .A3(new_n1102), .A4(new_n772), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1176), .A2(new_n1180), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1171), .B1(new_n1185), .B2(new_n766), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1168), .B1(new_n1169), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1167), .A2(new_n1187), .ZN(G378));
  NAND2_X1  g0988(.A1(new_n314), .A2(new_n363), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n304), .A2(new_n884), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1189), .B(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1191), .B(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n959), .B1(new_n958), .B2(new_n925), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n929), .A2(new_n961), .A3(KEYINPUT40), .ZN(new_n1195));
  OAI211_X1 g0995(.A(G330), .B(new_n1193), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1193), .B1(new_n963), .B2(G330), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n934), .B2(new_n950), .ZN(new_n1200));
  OAI21_X1  g1000(.A(KEYINPUT106), .B1(new_n932), .B2(new_n933), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n946), .A2(new_n935), .A3(new_n949), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1200), .A2(new_n1010), .A3(new_n1204), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1193), .A2(new_n761), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n823), .B1(G50), .B2(new_n837), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n772), .A2(new_n275), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G77), .B2(new_n783), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n202), .B2(new_n789), .C1(new_n845), .C2(new_n794), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT123), .Z(new_n1211));
  OAI22_X1  g1011(.A1(new_n786), .A2(new_n206), .B1(new_n792), .B2(new_n366), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G68), .B2(new_n810), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G97), .A2(new_n798), .B1(new_n800), .B2(G116), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1211), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n782), .A2(new_n1175), .B1(new_n792), .B2(new_n852), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G125), .A2(new_n800), .B1(new_n798), .B2(G132), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n252), .B2(new_n777), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(G128), .C2(new_n787), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1221), .B(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(G33), .B(G41), .C1(new_n795), .C2(G124), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n812), .C2(new_n789), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1208), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1217), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1207), .B1(new_n1228), .B2(new_n766), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1206), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1205), .A2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1203), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT57), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n1160), .B2(new_n1157), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n756), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1200), .A2(new_n1204), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1164), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1157), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1235), .B1(new_n1238), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1231), .B1(new_n1237), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(G375));
  OAI21_X1  g1044(.A(new_n293), .B1(new_n789), .B2(new_n202), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n855), .A2(new_n804), .B1(new_n844), .B2(new_n1175), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(G50), .C2(new_n810), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n852), .A2(new_n786), .B1(new_n782), .B2(new_n812), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n792), .A2(new_n252), .B1(new_n794), .B2(new_n1179), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n205), .A2(new_n782), .B1(new_n786), .B2(new_n845), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n792), .A2(new_n206), .B1(new_n794), .B2(new_n471), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n844), .A2(new_n449), .B1(new_n804), .B2(new_n841), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(new_n1254), .A2(new_n293), .A3(new_n1020), .A4(new_n1065), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1247), .A2(new_n1250), .B1(new_n1253), .B2(new_n1255), .ZN(new_n1256));
  OAI221_X1 g1056(.A(new_n823), .B1(G68), .B2(new_n837), .C1(new_n1256), .C2(new_n836), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1132), .B2(new_n760), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1151), .B2(new_n1010), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1151), .A2(new_n1157), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n991), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1259), .B1(new_n1260), .B2(new_n1263), .ZN(G381));
  INV_X1    g1064(.A(G378), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1085), .A2(new_n821), .ZN(new_n1266));
  NOR4_X1   g1066(.A1(G390), .A2(new_n1266), .A3(G384), .A4(G381), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1045), .A2(new_n1265), .A3(new_n1243), .A4(new_n1267), .ZN(G407));
  NAND2_X1  g1068(.A1(new_n699), .A2(G213), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1243), .A2(new_n1265), .A3(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G407), .A2(G213), .A3(new_n1271), .ZN(G409));
  NAND2_X1  g1072(.A1(G393), .A2(G396), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1273), .A2(new_n1266), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(G390), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT113), .B1(new_n1273), .B2(new_n1266), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1275), .B1(G390), .B2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(new_n1013), .A3(new_n1043), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1044), .B(new_n1275), .C1(G390), .C2(new_n1276), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(KEYINPUT61), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1230), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1282), .B1(new_n1234), .B2(new_n1010), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1160), .A2(new_n1157), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1234), .A2(new_n1262), .A3(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G378), .B1(new_n1283), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT57), .B1(new_n1234), .B2(new_n1284), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT57), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n720), .B1(new_n1238), .B2(new_n1289), .ZN(new_n1290));
  OAI211_X1 g1090(.A(G378), .B(new_n1283), .C1(new_n1288), .C2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT125), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT125), .B1(new_n1243), .B2(G378), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1287), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1295), .A2(new_n1296), .A3(new_n1269), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1237), .A2(new_n1242), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1299), .A2(KEYINPUT125), .A3(G378), .A4(new_n1283), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1286), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(KEYINPUT126), .B1(new_n1301), .B2(new_n1270), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT60), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1261), .B1(new_n1260), .B2(new_n1303), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1304), .B(new_n720), .C1(new_n1303), .C2(new_n1261), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1259), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1306), .B(G384), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1297), .A2(new_n1302), .A3(KEYINPUT63), .A4(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1295), .A2(new_n1269), .A3(new_n1307), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT63), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1270), .A2(G2897), .ZN(new_n1312));
  XOR2_X1   g1112(.A(new_n1307), .B(new_n1312), .Z(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n1270), .B2(new_n1301), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1281), .A2(new_n1308), .A3(new_n1311), .A4(new_n1314), .ZN(new_n1315));
  AND2_X1   g1115(.A1(new_n1307), .A2(KEYINPUT62), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1297), .A2(new_n1302), .A3(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1309), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT61), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1296), .B1(new_n1295), .B2(new_n1269), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1301), .A2(KEYINPUT126), .A3(new_n1270), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1313), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1320), .A2(KEYINPUT127), .A3(new_n1321), .A4(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(new_n1280), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1297), .A2(new_n1302), .ZN(new_n1327));
  AOI21_X1  g1127(.A(KEYINPUT61), .B1(new_n1327), .B2(new_n1313), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT127), .B1(new_n1328), .B2(new_n1320), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1315), .B1(new_n1326), .B2(new_n1329), .ZN(G405));
  OAI22_X1  g1130(.A1(new_n1293), .A2(new_n1294), .B1(G378), .B2(new_n1243), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(new_n1331), .B(new_n1307), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1280), .B(new_n1332), .ZN(G402));
endmodule


