//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:52 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n559, new_n560,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n604,
    new_n606, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1161;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT64), .B(G108), .Z(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G137), .ZN(new_n461));
  NAND2_X1  g036(.A1(G101), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT65), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n460), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n463), .B1(new_n473), .B2(G2105), .ZN(G160));
  NAND2_X1  g049(.A1(new_n465), .A2(new_n467), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n475), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT66), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(new_n476), .B2(G114), .ZN(new_n486));
  NOR2_X1   g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n489), .A2(new_n491), .A3(KEYINPUT67), .A4(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(KEYINPUT68), .B(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n460), .A2(new_n494), .A3(G138), .A4(new_n476), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n476), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n460), .A2(G126), .A3(G2105), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n493), .A2(new_n495), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT69), .A3(G651), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(new_n507), .B1(KEYINPUT6), .B2(new_n504), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(G50), .A3(G543), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n509), .B(KEYINPUT70), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(KEYINPUT71), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT5), .A3(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n517), .A2(new_n504), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n505), .A2(new_n507), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n513), .A2(new_n515), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n510), .A2(new_n518), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n521), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(new_n516), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n521), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n508), .A2(KEYINPUT72), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n534), .A2(G543), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(G51), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n530), .B(new_n532), .C1(new_n536), .C2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  INV_X1    g114(.A(new_n536), .ZN(new_n540));
  XOR2_X1   g115(.A(KEYINPUT73), .B(G52), .Z(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n504), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(G90), .B2(new_n523), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n536), .A2(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n508), .A2(new_n516), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n550), .A2(new_n551), .B1(new_n552), .B2(new_n504), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G188));
  NAND4_X1  g136(.A1(new_n534), .A2(G53), .A3(G543), .A4(new_n535), .ZN(new_n562));
  NAND2_X1  g137(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n563));
  OR2_X1    g138(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n522), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(G91), .A2(new_n523), .B1(new_n569), .B2(G651), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n570), .B1(new_n562), .B2(new_n563), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G299));
  NAND4_X1  g148(.A1(new_n534), .A2(G49), .A3(G543), .A4(new_n535), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n523), .A2(G87), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  AOI22_X1  g152(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(new_n504), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n516), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n521), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(G305));
  NAND2_X1  g157(.A1(new_n540), .A2(G47), .ZN(new_n583));
  NAND2_X1  g158(.A1(G72), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G60), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n522), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(G85), .A2(new_n523), .B1(new_n586), .B2(G651), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n508), .A2(G92), .A3(new_n516), .ZN(new_n590));
  XOR2_X1   g165(.A(new_n590), .B(KEYINPUT10), .Z(new_n591));
  NAND2_X1  g166(.A1(new_n540), .A2(G54), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n504), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n589), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n589), .B1(new_n596), .B2(G868), .ZN(G321));
  NAND2_X1  g173(.A1(G286), .A2(G868), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n572), .B(KEYINPUT76), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(G297));
  OAI21_X1  g176(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(G280));
  INV_X1    g177(.A(G860), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n595), .B1(G559), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT77), .ZN(G148));
  OR2_X1    g180(.A1(new_n595), .A2(G559), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g184(.A(new_n479), .ZN(new_n610));
  INV_X1    g185(.A(G135), .ZN(new_n611));
  OR3_X1    g186(.A1(new_n610), .A2(KEYINPUT79), .A3(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(KEYINPUT79), .B1(new_n610), .B2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n477), .A2(G123), .ZN(new_n614));
  OR2_X1    g189(.A1(G99), .A2(G2105), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n615), .B(G2104), .C1(G111), .C2(new_n476), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n612), .A2(new_n613), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(G2096), .Z(new_n618));
  NOR2_X1   g193(.A1(new_n464), .A2(G2105), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n460), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT78), .B(KEYINPUT13), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n618), .A2(new_n624), .ZN(G156));
  XOR2_X1   g200(.A(G2443), .B(G2446), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT81), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2451), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2435), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2438), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n629), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G14), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  NOR2_X1   g220(.A1(G2072), .A2(G2078), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n443), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT82), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT18), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n647), .A2(KEYINPUT83), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(KEYINPUT83), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(new_n645), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n647), .B(KEYINPUT84), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT17), .Z(new_n655));
  OAI211_X1 g230(.A(new_n653), .B(new_n644), .C1(new_n655), .C2(new_n645), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(new_n645), .A3(new_n643), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n650), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT85), .Z(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n663), .A2(new_n664), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n666), .A2(new_n668), .A3(new_n670), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n673), .B(new_n674), .C1(new_n672), .C2(new_n671), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1991), .B(G1996), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT22), .B(G1981), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(G229));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(KEYINPUT93), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(KEYINPUT93), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(G16), .A2(G22), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(G303), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(KEYINPUT91), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT91), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n692), .B(new_n688), .C1(G303), .C2(new_n689), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(G1971), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n691), .A2(G1971), .A3(new_n693), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AND3_X1   g273(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(KEYINPUT90), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT90), .ZN(new_n701));
  NAND2_X1  g276(.A1(G288), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G16), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT33), .B(G1976), .Z(new_n705));
  OAI211_X1 g280(.A(new_n704), .B(new_n705), .C1(G16), .C2(G23), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n704), .B1(G16), .B2(G23), .ZN(new_n707));
  INV_X1    g282(.A(new_n705), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n689), .A2(G6), .ZN(new_n710));
  INV_X1    g285(.A(G305), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n689), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT32), .B(G1981), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n698), .A2(new_n706), .A3(new_n709), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT89), .B(KEYINPUT34), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n477), .A2(G119), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT86), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n479), .A2(G131), .ZN(new_n724));
  NOR2_X1   g299(.A1(G95), .A2(G2105), .ZN(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(new_n476), .B2(G107), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OR3_X1    g302(.A1(new_n723), .A2(KEYINPUT87), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(KEYINPUT87), .B1(new_n723), .B2(new_n727), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n720), .B1(new_n731), .B2(new_n719), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT35), .B(G1991), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT88), .Z(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n732), .B(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT92), .ZN(new_n737));
  AND3_X1   g312(.A1(new_n715), .A2(new_n737), .A3(new_n716), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n715), .B2(new_n716), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n718), .B(new_n736), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G290), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G16), .B2(G24), .ZN(new_n743));
  INV_X1    g318(.A(G1986), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n685), .B(new_n687), .C1(new_n740), .C2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n739), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n715), .A2(new_n737), .A3(new_n716), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n717), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n745), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n749), .A2(new_n750), .A3(new_n736), .A4(new_n686), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n617), .A2(new_n719), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT101), .Z(new_n753));
  NOR2_X1   g328(.A1(G16), .A2(G21), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G168), .B2(G16), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT100), .B(G1966), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G35), .ZN(new_n758));
  OAI21_X1  g333(.A(KEYINPUT103), .B1(new_n758), .B2(G29), .ZN(new_n759));
  OR3_X1    g334(.A1(new_n758), .A2(KEYINPUT103), .A3(G29), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n759), .B(new_n760), .C1(G162), .C2(new_n719), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT29), .ZN(new_n762));
  OR3_X1    g337(.A1(new_n762), .A2(KEYINPUT104), .A3(G2090), .ZN(new_n763));
  NAND2_X1  g338(.A1(G164), .A2(G29), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G27), .B2(G29), .ZN(new_n765));
  INV_X1    g340(.A(G2078), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n479), .A2(G141), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT95), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n477), .A2(G129), .B1(G105), .B2(new_n619), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT96), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT26), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n769), .A2(new_n770), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n774), .A2(new_n719), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(KEYINPUT97), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G29), .B2(G32), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n776), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT27), .B(G1996), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT98), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  AND4_X1   g357(.A1(new_n757), .A2(new_n763), .A3(new_n767), .A4(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n689), .A2(KEYINPUT23), .A3(G20), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT23), .ZN(new_n785));
  INV_X1    g360(.A(G20), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(G16), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n787), .C1(new_n572), .C2(new_n689), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1956), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n762), .A2(G2090), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(KEYINPUT104), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n765), .A2(new_n766), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n762), .A2(G2090), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n783), .A2(new_n791), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n689), .A2(G5), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G171), .B2(new_n689), .ZN(new_n796));
  INV_X1    g371(.A(G1961), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G34), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n799), .A2(KEYINPUT24), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(KEYINPUT24), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n719), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G160), .B2(new_n719), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(G2084), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT102), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n798), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n719), .A2(G26), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n477), .A2(G128), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n479), .A2(G140), .ZN(new_n809));
  OR2_X1    g384(.A1(G104), .A2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n810), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n807), .B1(new_n813), .B2(new_n719), .ZN(new_n814));
  MUX2_X1   g389(.A(new_n807), .B(new_n814), .S(KEYINPUT28), .Z(new_n815));
  INV_X1    g390(.A(G2067), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT30), .B(G28), .Z(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(G29), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(KEYINPUT99), .B1(new_n779), .B2(new_n781), .ZN(new_n820));
  OR3_X1    g395(.A1(new_n779), .A2(KEYINPUT99), .A3(new_n781), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(KEYINPUT31), .B(G11), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n619), .A2(G103), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT25), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n479), .A2(G139), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n825), .B(new_n826), .C1(new_n476), .C2(new_n827), .ZN(new_n828));
  MUX2_X1   g403(.A(G33), .B(new_n828), .S(G29), .Z(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(G2072), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n803), .A2(G2084), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n822), .A2(new_n823), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n794), .A2(new_n806), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n746), .A2(new_n751), .A3(new_n753), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n554), .A2(new_n689), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n689), .B2(G19), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT94), .B(G1341), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n689), .A2(G4), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n596), .B2(new_n689), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(G1348), .Z(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n834), .A2(new_n838), .A3(new_n842), .ZN(G311));
  AND3_X1   g418(.A1(new_n746), .A2(new_n751), .A3(new_n833), .ZN(new_n844));
  INV_X1    g419(.A(new_n838), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n844), .A2(new_n845), .A3(new_n841), .A4(new_n753), .ZN(G150));
  NAND2_X1  g421(.A1(G80), .A2(G543), .ZN(new_n847));
  INV_X1    g422(.A(G67), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n522), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G651), .ZN(new_n850));
  INV_X1    g425(.A(G93), .ZN(new_n851));
  INV_X1    g426(.A(G55), .ZN(new_n852));
  OAI221_X1 g427(.A(new_n850), .B1(new_n851), .B2(new_n551), .C1(new_n536), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT37), .Z(new_n855));
  AOI22_X1  g430(.A1(G93), .A2(new_n523), .B1(new_n849), .B2(G651), .ZN(new_n856));
  OAI221_X1 g431(.A(new_n856), .B1(new_n852), .B2(new_n536), .C1(new_n549), .C2(new_n553), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n554), .A2(new_n853), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n596), .A2(G559), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT105), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n603), .B1(new_n862), .B2(KEYINPUT39), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n855), .B1(new_n864), .B2(new_n865), .ZN(G145));
  XNOR2_X1  g441(.A(G160), .B(KEYINPUT106), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(G162), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n617), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n476), .A2(G118), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT107), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n872));
  AOI22_X1  g447(.A1(G130), .A2(new_n477), .B1(new_n479), .B2(G142), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n869), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n730), .B(new_n774), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n828), .B(new_n813), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n621), .B(new_n501), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n876), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n875), .B(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g459(.A(KEYINPUT111), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT110), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n887));
  XNOR2_X1  g462(.A(G290), .B(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n700), .A2(G305), .A3(new_n702), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(G305), .B1(new_n700), .B2(new_n702), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G290), .B(KEYINPUT109), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n703), .A2(new_n711), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n889), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n895), .A3(G166), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(G166), .B1(new_n892), .B2(new_n895), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n892), .A2(new_n895), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(G303), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT42), .B1(new_n902), .B2(new_n896), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n886), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n899), .B1(new_n897), .B2(new_n898), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(KEYINPUT42), .A3(new_n896), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT110), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n606), .B(new_n859), .ZN(new_n908));
  NAND2_X1  g483(.A1(G299), .A2(new_n595), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n596), .A2(new_n572), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(KEYINPUT41), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n909), .A2(new_n915), .A3(new_n910), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(KEYINPUT108), .A3(new_n916), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n916), .A2(KEYINPUT108), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n908), .A3(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n904), .A2(new_n907), .A3(new_n913), .A4(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n900), .A2(new_n903), .ZN(new_n921));
  INV_X1    g496(.A(new_n919), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n921), .B(KEYINPUT110), .C1(new_n912), .C2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(G868), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n853), .A2(G868), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n885), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(G868), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(new_n920), .B2(new_n923), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n930), .A2(KEYINPUT111), .A3(new_n926), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n928), .A2(new_n931), .ZN(G295));
  NOR2_X1   g507(.A1(new_n930), .A2(new_n926), .ZN(G331));
  AOI21_X1  g508(.A(G286), .B1(new_n857), .B2(new_n858), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n857), .A2(new_n858), .A3(G286), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(G171), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n936), .ZN(new_n938));
  OAI21_X1  g513(.A(G301), .B1(new_n938), .B2(new_n934), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n917), .A2(new_n940), .A3(new_n918), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n902), .A2(new_n896), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n937), .A2(new_n939), .A3(new_n909), .A4(new_n910), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n882), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT43), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n942), .B1(new_n941), .B2(new_n943), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n942), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n914), .A2(new_n916), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n940), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n943), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n949), .A2(new_n952), .A3(KEYINPUT112), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT112), .B1(new_n949), .B2(new_n952), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n882), .B(new_n944), .C1(new_n954), .C2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n948), .B1(new_n956), .B2(new_n946), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n946), .B1(new_n945), .B2(new_n947), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(new_n956), .B2(new_n946), .ZN(new_n959));
  MUX2_X1   g534(.A(new_n957), .B(new_n959), .S(KEYINPUT44), .Z(G397));
  NAND2_X1  g535(.A1(new_n473), .A2(G2105), .ZN(new_n961));
  INV_X1    g536(.A(new_n463), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(G40), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n501), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT50), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n501), .A2(KEYINPUT50), .A3(new_n964), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G2090), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT115), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT114), .B(G1971), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n974), .A2(G40), .A3(G160), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT45), .B1(new_n501), .B2(new_n964), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n969), .A2(new_n978), .A3(new_n970), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n972), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT116), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n972), .A2(new_n982), .A3(new_n977), .A4(new_n979), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n981), .A2(G8), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G8), .ZN(new_n985));
  NOR2_X1   g560(.A1(G166), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(KEYINPUT117), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n989), .B1(new_n986), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n984), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1981), .ZN(new_n995));
  XNOR2_X1  g570(.A(G305), .B(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT49), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n963), .A2(new_n965), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(new_n985), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n703), .A2(G1976), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1002), .A2(KEYINPUT118), .A3(new_n999), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n699), .A2(G1976), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT52), .B1(new_n999), .B2(new_n1004), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1001), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n981), .A2(G8), .A3(new_n992), .A4(new_n983), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n756), .B1(new_n975), .B2(new_n976), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n961), .A2(G40), .A3(new_n962), .ZN(new_n1011));
  INV_X1    g586(.A(G2084), .ZN(new_n1012));
  INV_X1    g587(.A(new_n968), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT50), .B1(new_n501), .B2(new_n964), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n1011), .B(new_n1012), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1010), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G8), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G286), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n994), .A2(new_n1008), .A3(new_n1009), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT63), .ZN(new_n1020));
  INV_X1    g595(.A(G1976), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1021), .B(new_n699), .C1(new_n997), .C2(new_n1000), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n711), .A2(new_n995), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1000), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1009), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1024), .B1(new_n1025), .B2(new_n1008), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1020), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n975), .A2(new_n976), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n766), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1011), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1029), .A2(new_n1030), .B1(new_n797), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n965), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1033), .A2(KEYINPUT113), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(KEYINPUT113), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n975), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(KEYINPUT53), .A3(new_n766), .A4(new_n1038), .ZN(new_n1039));
  XOR2_X1   g614(.A(G301), .B(KEYINPUT54), .Z(new_n1040));
  AND3_X1   g615(.A1(new_n1032), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n998), .A2(new_n816), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n969), .B2(G1348), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1043), .A2(KEYINPUT60), .A3(new_n595), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n596), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1042), .B(new_n595), .C1(new_n969), .C2(G1348), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1044), .B1(new_n1047), .B2(KEYINPUT60), .ZN(new_n1048));
  XOR2_X1   g623(.A(KEYINPUT58), .B(G1341), .Z(new_n1049));
  OAI21_X1  g624(.A(new_n1049), .B1(new_n963), .B2(new_n965), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n976), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT121), .B(G1996), .Z(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1011), .A3(new_n974), .A4(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT122), .B(new_n1049), .C1(new_n963), .C2(new_n965), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1052), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1057), .A2(KEYINPUT59), .A3(new_n554), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT59), .B1(new_n1057), .B2(new_n554), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT61), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT56), .B(G2072), .ZN(new_n1062));
  INV_X1    g637(.A(G1956), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1028), .A2(new_n1062), .B1(new_n1031), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n571), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n569), .A2(G651), .ZN(new_n1067));
  INV_X1    g642(.A(G91), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1067), .B1(new_n551), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1066), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1065), .A2(new_n565), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n570), .B2(KEYINPUT119), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n566), .B2(new_n571), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1061), .B1(new_n1064), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1064), .A2(new_n1075), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1064), .A2(new_n1075), .A3(new_n1061), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1048), .A2(new_n1060), .A3(new_n1078), .A4(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1045), .B1(new_n1075), .B2(new_n1064), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1064), .B(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1075), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1041), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1032), .B1(new_n1030), .B2(new_n1029), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1040), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1016), .B2(G8), .ZN(new_n1092));
  AOI211_X1 g667(.A(KEYINPUT124), .B(new_n985), .C1(new_n1010), .C2(new_n1015), .ZN(new_n1093));
  NAND2_X1  g668(.A1(G286), .A2(G8), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT123), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n1094), .B(new_n1095), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1092), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1090), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1017), .A2(KEYINPUT124), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1096), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1016), .A2(new_n1091), .A3(G8), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(KEYINPUT125), .A3(KEYINPUT51), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1096), .A2(new_n1016), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1099), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1101), .A2(new_n1098), .A3(new_n1017), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1086), .A2(new_n1089), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  OR3_X1    g683(.A1(new_n1017), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n971), .A2(new_n977), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n993), .B1(new_n985), .B2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1008), .A2(new_n1009), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1027), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1106), .A2(KEYINPUT62), .A3(new_n1107), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n1117));
  AOI21_X1  g692(.A(G301), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1113), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1106), .A2(KEYINPUT126), .A3(KEYINPUT62), .A4(new_n1107), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1118), .A2(new_n1121), .A3(new_n1087), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1115), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1037), .A2(new_n963), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n731), .A2(new_n735), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n774), .A2(G1996), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n812), .B(new_n816), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n774), .A2(G1996), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1131), .B1(new_n734), .B2(new_n730), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1132), .B1(new_n744), .B2(new_n741), .ZN(new_n1133));
  NOR2_X1   g708(.A1(G290), .A2(G1986), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1125), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1124), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1125), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT46), .ZN(new_n1138));
  OR3_X1    g713(.A1(new_n1137), .A2(new_n1138), .A3(G1996), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1128), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1125), .B1(new_n774), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1138), .B1(new_n1137), .B2(G1996), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT47), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1130), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1145), .A2(new_n1126), .B1(G2067), .B2(new_n812), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1125), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1125), .A2(new_n1134), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT48), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1137), .B2(new_n1132), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1144), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT127), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1136), .A2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g728(.A1(new_n956), .A2(new_n946), .ZN(new_n1155));
  INV_X1    g729(.A(new_n948), .ZN(new_n1156));
  NAND3_X1  g730(.A1(new_n1155), .A2(G319), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g731(.A(new_n883), .ZN(new_n1158));
  NAND4_X1  g732(.A1(new_n641), .A2(new_n661), .A3(new_n682), .A4(new_n681), .ZN(new_n1159));
  NOR3_X1   g733(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(G308));
  INV_X1    g734(.A(new_n1159), .ZN(new_n1161));
  NAND4_X1  g735(.A1(new_n1161), .A2(new_n957), .A3(G319), .A4(new_n883), .ZN(G225));
endmodule


