//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1033, new_n1034;
  INV_X1    g000(.A(KEYINPUT4), .ZN(new_n202));
  AND2_X1   g001(.A1(G113gat), .A2(G120gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G113gat), .A2(G120gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT68), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G113gat), .ZN(new_n206));
  INV_X1    g005(.A(G120gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n209));
  NAND2_X1  g008(.A1(G113gat), .A2(G120gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n205), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G127gat), .A2(G134gat), .ZN(new_n214));
  INV_X1    g013(.A(G134gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT67), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G134gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n214), .B1(new_n219), .B2(G127gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n213), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(G127gat), .A2(G134gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n212), .B1(new_n222), .B2(new_n214), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n210), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT69), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n208), .A2(KEYINPUT69), .A3(new_n210), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G155gat), .B(G162gat), .ZN(new_n231));
  AND2_X1   g030(.A1(G141gat), .A2(G148gat), .ZN(new_n232));
  NOR2_X1   g031(.A1(G141gat), .A2(G148gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n235), .A2(KEYINPUT75), .A3(KEYINPUT2), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT75), .B1(new_n235), .B2(KEYINPUT2), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n231), .B(new_n234), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G141gat), .ZN(new_n239));
  INV_X1    g038(.A(G148gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT2), .ZN(new_n242));
  NAND2_X1  g041(.A1(G141gat), .A2(G148gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(G155gat), .A2(G162gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(G155gat), .A2(G162gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n244), .A2(KEYINPUT74), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT74), .B1(new_n244), .B2(new_n247), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n238), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n202), .B1(new_n230), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT74), .ZN(new_n252));
  NOR3_X1   g051(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT2), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(new_n231), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n244), .A2(KEYINPUT74), .A3(new_n247), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n236), .A2(new_n237), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n234), .A2(new_n231), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n254), .A2(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n223), .B1(new_n226), .B2(new_n225), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n259), .A2(new_n228), .B1(new_n213), .B2(new_n220), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT4), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n251), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT5), .ZN(new_n263));
  NAND2_X1  g062(.A1(G225gat), .A2(G233gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n266), .B(new_n238), .C1(new_n248), .C2(new_n249), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n230), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n262), .A2(new_n263), .A3(new_n264), .A4(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n268), .A2(new_n264), .A3(new_n251), .A4(new_n261), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n230), .A2(new_n250), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n255), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n272), .A2(new_n238), .A3(new_n221), .A4(new_n229), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n264), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n263), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n269), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G1gat), .B(G29gat), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n279), .B(KEYINPUT0), .ZN(new_n280));
  XNOR2_X1  g079(.A(G57gat), .B(G85gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n278), .A2(KEYINPUT6), .A3(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n277), .A3(new_n282), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(KEYINPUT76), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n282), .B1(new_n269), .B2(new_n277), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT76), .B1(new_n285), .B2(new_n286), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n284), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n293), .A2(G190gat), .ZN(new_n294));
  INV_X1    g093(.A(G190gat), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n295), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n294), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G169gat), .ZN(new_n300));
  INV_X1    g099(.A(G176gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT23), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n303), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n299), .B(new_n306), .C1(KEYINPUT64), .C2(KEYINPUT25), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT25), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n302), .A2(new_n304), .A3(KEYINPUT64), .A4(new_n305), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n295), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n293), .A2(G190gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n310), .B1(new_n311), .B2(new_n297), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n302), .A2(new_n304), .A3(new_n305), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n308), .B(new_n309), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT65), .ZN(new_n316));
  INV_X1    g115(.A(G183gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT27), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT27), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G183gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT66), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n316), .A2(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n317), .A2(KEYINPUT65), .A3(KEYINPUT27), .ZN(new_n323));
  NOR2_X1   g122(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n319), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  OR3_X1    g125(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n305), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n318), .A2(new_n320), .A3(new_n295), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n330), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n326), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G226gat), .ZN(new_n333));
  INV_X1    g132(.A(G233gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n315), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G197gat), .A2(G204gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(G197gat), .A2(G204gat), .ZN(new_n340));
  AND2_X1   g139(.A1(G211gat), .A2(G218gat), .ZN(new_n341));
  OAI22_X1  g140(.A1(new_n339), .A2(new_n340), .B1(new_n341), .B2(KEYINPUT22), .ZN(new_n342));
  NOR2_X1   g141(.A1(G211gat), .A2(G218gat), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT72), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  OR2_X1    g144(.A1(G197gat), .A2(G204gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT22), .ZN(new_n347));
  NAND2_X1  g146(.A1(G211gat), .A2(G218gat), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n346), .A2(new_n338), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OR2_X1    g148(.A1(G211gat), .A2(G218gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n351), .A3(new_n348), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n345), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n315), .A2(new_n332), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n335), .A2(KEYINPUT29), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n337), .B(new_n354), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n345), .A2(new_n353), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n315), .A2(new_n332), .A3(new_n336), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n356), .B1(new_n315), .B2(new_n332), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  NAND3_X1  g163(.A1(new_n357), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT73), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n366), .A2(KEYINPUT30), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n357), .A2(new_n361), .ZN(new_n368));
  INV_X1    g167(.A(new_n364), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(KEYINPUT30), .ZN(new_n371));
  AND3_X1   g170(.A1(new_n367), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n292), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT77), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n292), .A2(new_n375), .A3(new_n372), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT31), .B(G50gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G228gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(new_n334), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n341), .A2(new_n343), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n349), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n349), .B2(new_n385), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n266), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n389), .A2(new_n250), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n354), .B1(new_n267), .B2(new_n387), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n384), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n266), .B1(new_n358), .B2(KEYINPUT29), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n384), .B1(new_n394), .B2(new_n250), .ZN(new_n395));
  INV_X1    g194(.A(new_n391), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n393), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT3), .B1(new_n354), .B2(new_n387), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n383), .B1(new_n398), .B2(new_n258), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n399), .A2(new_n391), .A3(KEYINPUT79), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n392), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(G22gat), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n395), .A2(new_n393), .A3(new_n396), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT79), .B1(new_n399), .B2(new_n391), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G22gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(new_n392), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n381), .B1(new_n408), .B2(KEYINPUT78), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT78), .ZN(new_n410));
  AOI211_X1 g209(.A(new_n410), .B(new_n380), .C1(new_n402), .C2(new_n407), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n379), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n355), .A2(KEYINPUT70), .A3(new_n230), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n315), .A2(new_n332), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT70), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n260), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n230), .A2(KEYINPUT70), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n414), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n413), .A2(G227gat), .A3(G233gat), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT32), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  XOR2_X1   g221(.A(G15gat), .B(G43gat), .Z(new_n423));
  XNOR2_X1  g222(.A(G71gat), .B(G99gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n420), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n425), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n419), .B(KEYINPUT32), .C1(new_n421), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n413), .A2(new_n418), .B1(G227gat), .B2(G233gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT34), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT71), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n430), .B(KEYINPUT34), .Z(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(new_n426), .A3(new_n428), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n435), .B2(new_n432), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n401), .A2(G22gat), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n406), .B1(new_n405), .B2(new_n392), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT78), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n380), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n408), .A2(KEYINPUT78), .A3(new_n381), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n378), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n412), .A2(new_n436), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT35), .B1(new_n377), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n285), .A2(new_n286), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT80), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n278), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n269), .A2(new_n277), .A3(KEYINPUT80), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n445), .B1(new_n449), .B2(new_n283), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT82), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n284), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n288), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n372), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT83), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n372), .B(new_n457), .C1(new_n450), .C2(new_n454), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n429), .A2(new_n431), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n435), .A2(new_n460), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n412), .A2(new_n442), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AND3_X1   g263(.A1(new_n288), .A2(KEYINPUT82), .A3(KEYINPUT6), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT82), .B1(new_n288), .B2(KEYINPUT6), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(KEYINPUT37), .B1(new_n368), .B2(KEYINPUT81), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT38), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT81), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n357), .A2(new_n361), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n468), .A2(new_n469), .A3(new_n369), .A4(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n473), .A2(new_n365), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n269), .A2(new_n277), .A3(KEYINPUT80), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT80), .B1(new_n269), .B2(new_n277), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n283), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n445), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n468), .A2(new_n369), .A3(new_n472), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT38), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n467), .A2(new_n474), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n367), .A2(new_n370), .A3(new_n371), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n262), .A2(new_n268), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT39), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n275), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n282), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT40), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT39), .B1(new_n274), .B2(new_n275), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n489), .B1(new_n484), .B2(new_n275), .ZN(new_n490));
  OR3_X1    g289(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n488), .B1(new_n487), .B2(new_n490), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n483), .A2(new_n491), .A3(new_n477), .A4(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n482), .A2(new_n412), .A3(new_n442), .A4(new_n493), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n429), .A2(new_n432), .A3(new_n431), .ZN(new_n495));
  AOI22_X1  g294(.A1(new_n434), .A2(KEYINPUT71), .B1(new_n426), .B2(new_n428), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT36), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n435), .A2(new_n460), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n494), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n412), .A2(new_n442), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n377), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n444), .A2(new_n464), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G229gat), .A2(G233gat), .ZN(new_n506));
  AND2_X1   g305(.A1(G43gat), .A2(G50gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(G43gat), .A2(G50gat), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT15), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G29gat), .ZN(new_n511));
  INV_X1    g310(.A(G36gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT14), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT14), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(G29gat), .B2(G36gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT84), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT84), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n513), .A2(new_n515), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(G29gat), .A2(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AND4_X1   g320(.A1(new_n509), .A2(new_n515), .A3(new_n513), .A4(new_n520), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT15), .ZN(new_n523));
  OR2_X1    g322(.A1(KEYINPUT85), .A2(G43gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(KEYINPUT85), .A2(G43gat), .ZN(new_n525));
  AOI21_X1  g324(.A(G50gat), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g325(.A1(KEYINPUT86), .A2(G50gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(KEYINPUT86), .A2(G50gat), .ZN(new_n528));
  AOI21_X1  g327(.A(G43gat), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n523), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n510), .A2(new_n521), .B1(new_n522), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n531), .A2(KEYINPUT17), .ZN(new_n532));
  INV_X1    g331(.A(G1gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT16), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n406), .A2(G15gat), .ZN(new_n535));
  INV_X1    g334(.A(G15gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(G22gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT87), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n538), .B1(new_n535), .B2(new_n537), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n534), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G8gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n536), .A2(G22gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n406), .A2(G15gat), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT87), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n535), .A2(new_n537), .A3(new_n538), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n545), .A2(new_n533), .A3(new_n546), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n541), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n542), .B1(new_n541), .B2(new_n547), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n531), .A2(KEYINPUT17), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n532), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT88), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(new_n548), .B2(new_n549), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n539), .A2(new_n540), .A3(G1gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n534), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n556), .B1(new_n545), .B2(new_n546), .ZN(new_n557));
  OAI21_X1  g356(.A(G8gat), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n547), .A3(new_n542), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(KEYINPUT88), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n531), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT89), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT89), .ZN(new_n564));
  AOI211_X1 g363(.A(new_n564), .B(new_n531), .C1(new_n554), .C2(new_n560), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n506), .B(new_n552), .C1(new_n563), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT90), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT18), .ZN(new_n568));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G197gat), .ZN(new_n570));
  XOR2_X1   g369(.A(KEYINPUT11), .B(G169gat), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT12), .Z(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT18), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n566), .A2(KEYINPUT90), .A3(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(new_n506), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR3_X1   g378(.A1(new_n548), .A2(new_n549), .A3(new_n553), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT88), .B1(new_n558), .B2(new_n559), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n562), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n564), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n561), .A2(KEYINPUT89), .A3(new_n562), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n561), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n531), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n579), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n568), .A2(new_n574), .A3(new_n576), .A4(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n588), .B1(new_n567), .B2(KEYINPUT18), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n574), .B1(new_n592), .B2(new_n576), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT7), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(KEYINPUT96), .A2(KEYINPUT7), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n600), .A2(G85gat), .A3(G92gat), .A4(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G85gat), .ZN(new_n603));
  INV_X1    g402(.A(G92gat), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n598), .B(new_n599), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n606), .B1(new_n603), .B2(new_n604), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n608), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n606), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n602), .A2(new_n611), .A3(new_n605), .A4(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g412(.A(G57gat), .B(G64gat), .Z(new_n614));
  INV_X1    g413(.A(KEYINPUT9), .ZN(new_n615));
  INV_X1    g414(.A(G71gat), .ZN(new_n616));
  INV_X1    g415(.A(G78gat), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(KEYINPUT92), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G71gat), .B(G78gat), .Z(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n623));
  INV_X1    g422(.A(G64gat), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n624), .A2(G57gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(G57gat), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(new_n627), .A3(new_n618), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n621), .A2(new_n628), .A3(KEYINPUT93), .ZN(new_n629));
  AOI21_X1  g428(.A(KEYINPUT93), .B1(new_n621), .B2(new_n628), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n613), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n610), .A2(new_n612), .ZN(new_n632));
  INV_X1    g431(.A(new_n628), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n622), .B1(new_n627), .B2(new_n618), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n597), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n632), .B(KEYINPUT10), .C1(new_n629), .C2(new_n630), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n596), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n596), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n631), .A2(new_n635), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G176gat), .B(G204gat), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n642), .B(new_n643), .Z(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT102), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n639), .A2(new_n647), .A3(new_n641), .A4(new_n644), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n639), .A2(new_n641), .ZN(new_n650));
  INV_X1    g449(.A(new_n644), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G232gat), .A2(G233gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT95), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(KEYINPUT41), .ZN(new_n657));
  XNOR2_X1  g456(.A(G134gat), .B(G162gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  AND2_X1   g458(.A1(new_n659), .A2(KEYINPUT100), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(KEYINPUT100), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n613), .B(KEYINPUT97), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n663), .A2(new_n532), .A3(new_n551), .ZN(new_n664));
  AOI22_X1  g463(.A1(new_n562), .A2(new_n632), .B1(KEYINPUT41), .B2(new_n656), .ZN(new_n665));
  XNOR2_X1  g464(.A(G190gat), .B(G218gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n664), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n669), .B1(new_n664), .B2(new_n665), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n662), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n672), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n660), .A3(new_n670), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(G155gat), .Z(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT21), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n629), .A2(new_n630), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n586), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n683), .A2(KEYINPUT94), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(KEYINPUT94), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n680), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(G183gat), .B(G211gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n682), .A2(new_n681), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(G231gat), .A3(G233gat), .ZN(new_n690));
  INV_X1    g489(.A(G127gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(G231gat), .A2(G233gat), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n682), .A2(new_n681), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n690), .A2(new_n691), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n691), .B1(new_n690), .B2(new_n693), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n688), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n696), .ZN(new_n698));
  INV_X1    g497(.A(new_n688), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n699), .A3(new_n694), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n680), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n687), .A2(new_n697), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n697), .A2(new_n700), .ZN(new_n703));
  INV_X1    g502(.A(new_n701), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(new_n686), .ZN(new_n705));
  AOI211_X1 g504(.A(new_n653), .B(new_n677), .C1(new_n702), .C2(new_n705), .ZN(new_n706));
  AND3_X1   g505(.A1(new_n505), .A2(new_n595), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n292), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g509(.A(KEYINPUT16), .B(G8gat), .Z(new_n711));
  AND3_X1   g510(.A1(new_n707), .A2(new_n483), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n542), .B1(new_n707), .B2(new_n483), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT42), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(KEYINPUT42), .B2(new_n712), .ZN(G1325gat));
  INV_X1    g514(.A(new_n500), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n536), .B1(new_n707), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n461), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(G15gat), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n717), .B1(new_n707), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT103), .ZN(G1326gat));
  NAND2_X1  g520(.A1(new_n707), .A2(new_n502), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT43), .B(G22gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1327gat));
  NAND2_X1  g523(.A1(new_n702), .A2(new_n705), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n594), .A2(new_n725), .A3(new_n653), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n504), .A2(new_n676), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n708), .A2(new_n511), .ZN(new_n730));
  OR3_X1    g529(.A1(new_n729), .A2(KEYINPUT104), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT104), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n412), .A2(new_n442), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n736), .A2(new_n374), .A3(new_n376), .A4(new_n436), .ZN(new_n737));
  AOI21_X1  g536(.A(KEYINPUT35), .B1(new_n456), .B2(new_n458), .ZN(new_n738));
  AOI22_X1  g537(.A1(new_n737), .A2(KEYINPUT35), .B1(new_n738), .B2(new_n462), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n494), .A2(new_n500), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n377), .B2(new_n502), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT105), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n444), .A2(new_n464), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n501), .A2(new_n503), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n676), .A2(KEYINPUT44), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n742), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT44), .B1(new_n504), .B2(new_n676), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n727), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(G29gat), .B1(new_n751), .B2(new_n292), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n731), .A2(KEYINPUT45), .A3(new_n732), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n735), .A2(new_n752), .A3(new_n753), .ZN(G1328gat));
  OAI21_X1  g553(.A(G36gat), .B1(new_n751), .B2(new_n372), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n483), .A2(new_n512), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT46), .B1(new_n729), .B2(new_n756), .ZN(new_n757));
  OR3_X1    g556(.A1(new_n729), .A2(KEYINPUT46), .A3(new_n756), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(G1329gat));
  AOI22_X1  g558(.A1(new_n750), .A2(new_n716), .B1(new_n524), .B2(new_n525), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n461), .A2(new_n524), .A3(new_n525), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n505), .A2(new_n677), .A3(new_n726), .A4(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT47), .B1(new_n762), .B2(KEYINPUT106), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI211_X1 g566(.A(KEYINPUT107), .B(KEYINPUT47), .C1(new_n762), .C2(KEYINPUT106), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n760), .A2(new_n763), .B1(new_n767), .B2(new_n768), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(G1330gat));
  NAND2_X1  g571(.A1(new_n527), .A2(new_n528), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n729), .A2(new_n736), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI211_X1 g575(.A(new_n736), .B(new_n727), .C1(new_n748), .C2(new_n749), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n773), .B1(new_n777), .B2(KEYINPUT108), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n750), .A2(KEYINPUT108), .A3(new_n502), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n750), .A2(new_n502), .B1(new_n527), .B2(new_n528), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n775), .B1(new_n781), .B2(new_n774), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1331gat));
  AND2_X1   g582(.A1(new_n742), .A2(new_n746), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n292), .B(KEYINPUT109), .ZN(new_n785));
  INV_X1    g584(.A(new_n725), .ZN(new_n786));
  INV_X1    g585(.A(new_n653), .ZN(new_n787));
  NOR4_X1   g586(.A1(new_n595), .A2(new_n786), .A3(new_n677), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n784), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g589(.A(new_n372), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n784), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT110), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n784), .A2(new_n794), .A3(new_n788), .A4(new_n791), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(G1333gat));
  NAND2_X1  g597(.A1(new_n784), .A2(new_n788), .ZN(new_n799));
  OAI21_X1  g598(.A(G71gat), .B1(new_n799), .B2(new_n500), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n461), .A2(new_n616), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n800), .B(KEYINPUT50), .C1(new_n799), .C2(new_n801), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1334gat));
  NOR2_X1   g605(.A1(new_n799), .A2(new_n736), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(new_n617), .ZN(G1335gat));
  NOR2_X1   g607(.A1(new_n595), .A2(new_n787), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n786), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n748), .B2(new_n749), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G85gat), .B1(new_n812), .B2(new_n292), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n504), .B2(new_n676), .ZN(new_n815));
  OAI211_X1 g614(.A(KEYINPUT111), .B(new_n677), .C1(new_n739), .C2(new_n741), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n595), .A2(new_n725), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n815), .A2(KEYINPUT51), .A3(new_n816), .A4(new_n817), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n653), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n708), .A2(new_n603), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n813), .B1(new_n823), .B2(new_n824), .ZN(G1336gat));
  NOR2_X1   g624(.A1(new_n372), .A2(G92gat), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n818), .A2(new_n819), .ZN(new_n828));
  AOI211_X1 g627(.A(new_n787), .B(new_n827), .C1(new_n828), .C2(new_n821), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n604), .B1(new_n811), .B2(new_n483), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT52), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n653), .B(new_n826), .C1(new_n820), .C2(new_n822), .ZN(new_n832));
  INV_X1    g631(.A(new_n830), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n831), .A2(new_n835), .ZN(G1337gat));
  OAI21_X1  g635(.A(G99gat), .B1(new_n812), .B2(new_n500), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n718), .A2(G99gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n823), .B2(new_n838), .ZN(G1338gat));
  INV_X1    g638(.A(G106gat), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n502), .A2(new_n840), .A3(new_n653), .ZN(new_n841));
  XOR2_X1   g640(.A(new_n841), .B(KEYINPUT112), .Z(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n843), .B1(new_n828), .B2(new_n821), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n840), .B1(new_n811), .B2(new_n502), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT53), .B1(new_n844), .B2(new_n845), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1339gat));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n706), .A2(new_n594), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  INV_X1    g652(.A(new_n597), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT93), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n633), .B2(new_n634), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n621), .A2(new_n628), .A3(KEYINPUT93), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n632), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n613), .B1(new_n628), .B2(new_n621), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n640), .A3(new_n637), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n861), .A2(new_n639), .A3(KEYINPUT54), .ZN(new_n862));
  XOR2_X1   g661(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n651), .B1(new_n639), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n853), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n640), .B1(new_n860), .B2(new_n637), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n644), .B1(new_n867), .B2(new_n863), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n861), .A2(new_n639), .A3(KEYINPUT54), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n869), .A3(KEYINPUT55), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n866), .A2(new_n649), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n585), .A2(new_n587), .A3(new_n579), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n532), .A2(new_n551), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n583), .A2(new_n584), .B1(new_n873), .B2(new_n550), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n872), .B1(new_n874), .B2(new_n506), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n572), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n871), .A2(new_n590), .A3(new_n677), .A4(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n871), .B1(new_n591), .B2(new_n593), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n590), .A2(new_n653), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT114), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT114), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n590), .A2(new_n653), .A3(new_n882), .A4(new_n876), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n879), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n878), .B1(new_n884), .B2(new_n676), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n852), .B1(new_n885), .B2(new_n725), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(new_n462), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n708), .A2(new_n372), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n595), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n851), .B1(new_n892), .B2(G113gat), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT115), .B(new_n206), .C1(new_n891), .C2(new_n595), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n886), .A2(new_n785), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n443), .A2(new_n483), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT116), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n595), .A2(new_n206), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n893), .A2(new_n894), .B1(new_n898), .B2(new_n899), .ZN(G1340gat));
  OAI21_X1  g699(.A(G120gat), .B1(new_n890), .B2(new_n787), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n653), .A2(new_n207), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n898), .B2(new_n902), .ZN(G1341gat));
  OAI21_X1  g702(.A(new_n691), .B1(new_n897), .B2(new_n786), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n786), .A2(new_n691), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT117), .B1(new_n890), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n890), .A2(KEYINPUT117), .A3(new_n906), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(G1342gat));
  NOR2_X1   g709(.A1(new_n676), .A2(new_n219), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n896), .A3(new_n911), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(KEYINPUT118), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(KEYINPUT118), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT56), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G134gat), .B1(new_n890), .B2(new_n676), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n913), .A2(KEYINPUT56), .A3(new_n914), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(G1343gat));
  NOR3_X1   g719(.A1(new_n716), .A2(new_n483), .A3(new_n736), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n895), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n239), .A3(new_n595), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n716), .A2(new_n888), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT57), .B1(new_n886), .B2(new_n502), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n502), .A2(KEYINPUT57), .ZN(new_n926));
  XOR2_X1   g725(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n927));
  OAI21_X1  g726(.A(new_n927), .B1(new_n862), .B2(new_n865), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(new_n649), .A3(new_n870), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n929), .B1(new_n591), .B2(new_n593), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n677), .B1(new_n930), .B2(new_n880), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n786), .B1(new_n931), .B2(new_n878), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n926), .B1(new_n932), .B2(new_n852), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n595), .B(new_n924), .C1(new_n925), .C2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n923), .B1(new_n239), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT58), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(KEYINPUT120), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n239), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT58), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n923), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n937), .B1(new_n941), .B2(new_n943), .ZN(G1344gat));
  INV_X1    g743(.A(KEYINPUT59), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n924), .B1(new_n925), .B2(new_n933), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n945), .B(G148gat), .C1(new_n946), .C2(new_n787), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n928), .A2(new_n649), .A3(new_n870), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n568), .A2(new_n576), .A3(new_n589), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n573), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n948), .B1(new_n950), .B2(new_n590), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n590), .A2(new_n653), .A3(new_n876), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n676), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n725), .B1(new_n953), .B2(new_n877), .ZN(new_n954));
  INV_X1    g753(.A(new_n852), .ZN(new_n955));
  OAI21_X1  g754(.A(KEYINPUT122), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n932), .A2(new_n957), .A3(new_n852), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n956), .A2(new_n958), .A3(new_n502), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT57), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT121), .ZN(new_n962));
  INV_X1    g761(.A(new_n926), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n886), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n886), .A2(new_n963), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT121), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n961), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n716), .A2(new_n787), .A3(new_n888), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n240), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n947), .B1(new_n969), .B2(new_n945), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n922), .A2(new_n240), .A3(new_n653), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(G1345gat));
  OAI21_X1  g771(.A(G155gat), .B1(new_n946), .B2(new_n786), .ZN(new_n973));
  INV_X1    g772(.A(new_n922), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n786), .A2(G155gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n973), .B1(new_n974), .B2(new_n975), .ZN(G1346gat));
  INV_X1    g775(.A(G162gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n977), .B1(new_n974), .B2(new_n676), .ZN(new_n978));
  OR3_X1    g777(.A1(new_n946), .A2(new_n977), .A3(new_n676), .ZN(new_n979));
  AND2_X1   g778(.A1(new_n978), .A2(new_n979), .ZN(G1347gat));
  NOR2_X1   g779(.A1(new_n785), .A2(new_n372), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n887), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n982), .A2(new_n300), .A3(new_n594), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n886), .A2(new_n292), .A3(new_n483), .ZN(new_n984));
  INV_X1    g783(.A(new_n443), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(new_n595), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n983), .B1(new_n988), .B2(new_n300), .ZN(G1348gat));
  OAI21_X1  g788(.A(new_n301), .B1(new_n986), .B2(new_n787), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n653), .A2(G176gat), .ZN(new_n991));
  OAI21_X1  g790(.A(KEYINPUT123), .B1(new_n982), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  NOR3_X1   g792(.A1(new_n982), .A2(KEYINPUT123), .A3(new_n991), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n993), .A2(new_n994), .ZN(G1349gat));
  OAI21_X1  g794(.A(G183gat), .B1(new_n982), .B2(new_n786), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n725), .A2(new_n318), .A3(new_n320), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n996), .B1(new_n986), .B2(new_n997), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n998), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g798(.A1(new_n886), .A2(new_n462), .A3(new_n677), .A4(new_n981), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(G190gat), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n1002));
  OR3_X1    g801(.A1(new_n1001), .A2(new_n1002), .A3(KEYINPUT61), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1001), .A2(KEYINPUT61), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT124), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1001), .A2(KEYINPUT124), .A3(KEYINPUT61), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1002), .B1(new_n1001), .B2(KEYINPUT61), .ZN(new_n1008));
  NAND4_X1  g807(.A1(new_n1003), .A2(new_n1006), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n987), .A2(new_n295), .A3(new_n677), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(G1351gat));
  NOR3_X1   g810(.A1(new_n716), .A2(new_n785), .A3(new_n372), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n967), .A2(new_n595), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1013), .A2(KEYINPUT126), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1015));
  NAND4_X1  g814(.A1(new_n967), .A2(new_n1015), .A3(new_n595), .A4(new_n1012), .ZN(new_n1016));
  NAND3_X1  g815(.A1(new_n1014), .A2(G197gat), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g816(.A1(new_n716), .A2(new_n736), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n984), .A2(new_n1018), .ZN(new_n1019));
  OR3_X1    g818(.A1(new_n1019), .A2(G197gat), .A3(new_n594), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1017), .A2(new_n1020), .ZN(G1352gat));
  XOR2_X1   g820(.A(KEYINPUT127), .B(G204gat), .Z(new_n1022));
  NOR3_X1   g821(.A1(new_n1019), .A2(new_n787), .A3(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g822(.A(new_n1023), .B(KEYINPUT62), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n967), .A2(new_n1012), .ZN(new_n1025));
  OAI21_X1  g824(.A(new_n1022), .B1(new_n1025), .B2(new_n787), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1024), .A2(new_n1026), .ZN(G1353gat));
  OR3_X1    g826(.A1(new_n1019), .A2(G211gat), .A3(new_n786), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n967), .A2(new_n725), .A3(new_n1012), .ZN(new_n1029));
  AND3_X1   g828(.A1(new_n1029), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1030));
  AOI21_X1  g829(.A(KEYINPUT63), .B1(new_n1029), .B2(G211gat), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n1028), .B1(new_n1030), .B2(new_n1031), .ZN(G1354gat));
  OAI21_X1  g831(.A(G218gat), .B1(new_n1025), .B2(new_n676), .ZN(new_n1033));
  OR2_X1    g832(.A1(new_n676), .A2(G218gat), .ZN(new_n1034));
  OAI21_X1  g833(.A(new_n1033), .B1(new_n1019), .B2(new_n1034), .ZN(G1355gat));
endmodule


