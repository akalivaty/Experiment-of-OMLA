//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203));
  INV_X1    g002(.A(G71gat), .ZN(new_n204));
  INV_X1    g003(.A(G78gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(G71gat), .B(G78gat), .Z(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G231gat), .A2(G233gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(G127gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT93), .ZN(new_n216));
  INV_X1    g015(.A(G1gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(KEYINPUT93), .A3(G1gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n218), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(G8gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(new_n210), .B2(new_n209), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT95), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n214), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(G155gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(G183gat), .B(G211gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n227), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G190gat), .B(G218gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G85gat), .A2(G92gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT7), .ZN(new_n236));
  XNOR2_X1  g035(.A(G99gat), .B(G106gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(G99gat), .A2(G106gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n238), .B1(KEYINPUT8), .B2(new_n239), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n236), .A2(new_n237), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n237), .B1(new_n236), .B2(new_n240), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XOR2_X1   g042(.A(G43gat), .B(G50gat), .Z(new_n244));
  INV_X1    g043(.A(KEYINPUT15), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G29gat), .ZN(new_n247));
  INV_X1    g046(.A(G36gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  OR3_X1    g049(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n244), .A2(KEYINPUT92), .A3(new_n245), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT92), .B1(new_n244), .B2(new_n245), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n250), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n251), .A2(KEYINPUT91), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n252), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n251), .A2(KEYINPUT91), .ZN(new_n259));
  OAI22_X1  g058(.A1(new_n258), .A2(new_n259), .B1(new_n247), .B2(new_n248), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n246), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT17), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT17), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n256), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n243), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(G232gat), .A2(G233gat), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n262), .A2(new_n243), .B1(KEYINPUT41), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n234), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(new_n241), .A2(new_n242), .ZN(new_n271));
  INV_X1    g070(.A(new_n265), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n264), .B1(new_n256), .B2(new_n261), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n274), .A2(new_n268), .A3(new_n233), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n267), .A2(KEYINPUT41), .ZN(new_n276));
  XNOR2_X1  g075(.A(G134gat), .B(G162gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n276), .B(new_n277), .Z(new_n278));
  XOR2_X1   g077(.A(new_n278), .B(KEYINPUT96), .Z(new_n279));
  NAND3_X1  g078(.A1(new_n270), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT97), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n270), .A2(new_n275), .ZN(new_n282));
  INV_X1    g081(.A(new_n278), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT97), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n270), .A2(new_n285), .A3(new_n275), .A4(new_n279), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n281), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G230gat), .A2(G233gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n209), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT10), .ZN(new_n292));
  INV_X1    g091(.A(new_n208), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n207), .B(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n243), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n291), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n243), .A3(KEYINPUT10), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n290), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n291), .A2(new_n295), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n298), .B1(new_n299), .B2(new_n290), .ZN(new_n300));
  XNOR2_X1  g099(.A(G120gat), .B(G148gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(G176gat), .B(G204gat), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n301), .B(new_n302), .Z(new_n303));
  OR2_X1    g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n296), .A2(new_n297), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(new_n289), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n299), .A2(new_n290), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n307), .A3(new_n303), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n232), .A2(new_n288), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT98), .ZN(new_n313));
  INV_X1    g112(.A(new_n262), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(new_n224), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n222), .B(G8gat), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n316), .B1(new_n263), .B2(new_n265), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT94), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n315), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G229gat), .A2(G233gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n224), .B1(new_n272), .B2(new_n273), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT94), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT18), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n319), .A2(new_n322), .A3(KEYINPUT18), .A4(new_n320), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n316), .B(new_n262), .ZN(new_n327));
  XOR2_X1   g126(.A(new_n320), .B(KEYINPUT13), .Z(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G113gat), .B(G141gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(G197gat), .ZN(new_n332));
  XOR2_X1   g131(.A(KEYINPUT11), .B(G169gat), .Z(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n334), .B(KEYINPUT12), .Z(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  AOI22_X1  g135(.A1(new_n323), .A2(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n337));
  INV_X1    g136(.A(new_n335), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n326), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT98), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n311), .A2(new_n341), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n313), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G127gat), .B(G134gat), .Z(new_n344));
  XNOR2_X1  g143(.A(G113gat), .B(G120gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(KEYINPUT1), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G113gat), .B(G120gat), .Z(new_n347));
  INV_X1    g146(.A(KEYINPUT1), .ZN(new_n348));
  XNOR2_X1  g147(.A(G127gat), .B(G134gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G141gat), .B(G148gat), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n353));
  NAND2_X1  g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n353), .B1(new_n354), .B2(KEYINPUT2), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  OR2_X1    g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(new_n354), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n354), .A2(new_n353), .A3(KEYINPUT2), .ZN(new_n360));
  AND2_X1   g159(.A1(G155gat), .A2(G162gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT79), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n356), .A2(new_n359), .A3(new_n360), .A4(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT2), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT78), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n354), .A2(new_n367), .A3(KEYINPUT2), .ZN(new_n368));
  AND2_X1   g167(.A1(G141gat), .A2(G148gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n361), .A2(new_n362), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n364), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n351), .B1(new_n375), .B2(KEYINPUT3), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n359), .A2(new_n363), .A3(new_n360), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n378), .A2(new_n356), .B1(new_n373), .B2(new_n372), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n377), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AND4_X1   g180(.A1(new_n377), .A2(new_n364), .A3(new_n374), .A4(new_n380), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n376), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT5), .ZN(new_n384));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n351), .A2(new_n374), .A3(new_n364), .ZN(new_n387));
  OR3_X1    g186(.A1(new_n387), .A2(KEYINPUT86), .A3(KEYINPUT4), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n346), .A2(new_n350), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT4), .B1(new_n375), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n379), .A2(new_n391), .A3(new_n351), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n390), .A2(new_n392), .A3(KEYINPUT86), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n386), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n390), .A2(new_n392), .A3(KEYINPUT82), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT82), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n387), .A2(new_n397), .A3(KEYINPUT4), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n383), .A2(new_n385), .A3(new_n396), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n375), .A2(new_n389), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n387), .ZN(new_n401));
  INV_X1    g200(.A(new_n385), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n384), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(KEYINPUT83), .A3(new_n403), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n395), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  XOR2_X1   g207(.A(G1gat), .B(G29gat), .Z(new_n409));
  XNOR2_X1  g208(.A(new_n409), .B(KEYINPUT85), .ZN(new_n410));
  XOR2_X1   g209(.A(G57gat), .B(G85gat), .Z(new_n411));
  XNOR2_X1  g210(.A(new_n410), .B(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT87), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT6), .B1(new_n408), .B2(new_n414), .ZN(new_n416));
  INV_X1    g215(.A(new_n395), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n399), .A2(KEYINPUT83), .A3(new_n403), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT83), .B1(new_n399), .B2(new_n403), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n421));
  INV_X1    g220(.A(new_n414), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n415), .A2(new_n416), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n420), .A2(KEYINPUT6), .A3(new_n422), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  XOR2_X1   g228(.A(new_n429), .B(KEYINPUT76), .Z(new_n430));
  INV_X1    g229(.A(KEYINPUT72), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT22), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n431), .A2(new_n432), .B1(G211gat), .B2(G218gat), .ZN(new_n433));
  NAND2_X1  g232(.A1(KEYINPUT72), .A2(KEYINPUT22), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT73), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(G211gat), .B(G218gat), .Z(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n431), .A2(new_n432), .ZN(new_n440));
  NAND2_X1  g239(.A1(G211gat), .A2(G218gat), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n440), .A2(KEYINPUT73), .A3(new_n441), .A4(new_n434), .ZN(new_n442));
  XNOR2_X1  g241(.A(G197gat), .B(G204gat), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n437), .A2(new_n439), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n443), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT73), .B1(new_n433), .B2(new_n434), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n438), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(G226gat), .ZN(new_n449));
  INV_X1    g248(.A(G233gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(G169gat), .ZN(new_n452));
  INV_X1    g251(.A(G176gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT26), .ZN(new_n455));
  NAND2_X1  g254(.A1(G169gat), .A2(G176gat), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(G169gat), .A2(G176gat), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n458), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n457), .A2(new_n459), .A3(KEYINPUT68), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT27), .B(G183gat), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT28), .ZN(new_n465));
  INV_X1    g264(.A(G190gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n466), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT28), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n462), .A2(new_n463), .A3(new_n467), .A4(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(G183gat), .A2(G190gat), .ZN(new_n471));
  AND2_X1   g270(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n471), .B1(new_n472), .B2(G190gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(G183gat), .A2(G190gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT24), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT66), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n473), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n452), .A2(new_n453), .A3(KEYINPUT23), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT23), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(G169gat), .B2(G176gat), .ZN(new_n484));
  AND4_X1   g283(.A1(KEYINPUT25), .A2(new_n482), .A3(new_n484), .A4(new_n456), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT67), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n481), .A2(new_n485), .A3(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(G183gat), .B2(G190gat), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT64), .B1(new_n474), .B2(new_n475), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT64), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n482), .A2(new_n484), .A3(new_n456), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n494), .A2(new_n495), .B1(new_n496), .B2(KEYINPUT65), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n482), .A2(new_n484), .A3(new_n498), .A4(new_n456), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT25), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n470), .B1(new_n490), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT29), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n451), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND4_X1   g302(.A1(new_n462), .A2(new_n463), .A3(new_n467), .A4(new_n469), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n481), .A2(new_n485), .A3(KEYINPUT67), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT67), .B1(new_n481), .B2(new_n485), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT64), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n476), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n473), .A2(new_n509), .A3(new_n495), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n456), .B1(new_n458), .B2(KEYINPUT23), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n483), .A2(G169gat), .A3(G176gat), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT65), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n513), .A3(new_n499), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT25), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n504), .B1(new_n507), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n451), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT74), .B1(new_n503), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT74), .B1(new_n501), .B2(new_n451), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n448), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT75), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(new_n488), .A3(new_n489), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT29), .B1(new_n525), .B2(new_n470), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n524), .B1(new_n526), .B2(new_n451), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n501), .A2(new_n451), .ZN(new_n528));
  OAI211_X1 g327(.A(KEYINPUT75), .B(new_n518), .C1(new_n517), .C2(KEYINPUT29), .ZN(new_n529));
  AND4_X1   g328(.A1(new_n448), .A2(new_n527), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n430), .B1(new_n523), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT77), .ZN(new_n532));
  INV_X1    g331(.A(new_n448), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT74), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n518), .B1(new_n517), .B2(KEYINPUT29), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(new_n528), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n533), .B1(new_n536), .B2(new_n521), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n527), .A2(new_n529), .A3(new_n448), .A4(new_n528), .ZN(new_n538));
  INV_X1    g337(.A(new_n429), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n531), .A2(new_n532), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n538), .A3(new_n429), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n540), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n532), .B1(new_n531), .B2(new_n542), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n525), .A2(new_n351), .A3(new_n470), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT69), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G227gat), .A2(G233gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n501), .A2(new_n389), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n525), .A2(KEYINPUT69), .A3(new_n351), .A4(new_n470), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT70), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n557), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(KEYINPUT70), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT32), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n551), .A2(new_n554), .A3(new_n553), .ZN(new_n563));
  INV_X1    g362(.A(new_n552), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT33), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  XOR2_X1   g365(.A(G15gat), .B(G43gat), .Z(new_n567));
  XNOR2_X1  g366(.A(G71gat), .B(G99gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n565), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  AOI221_X4 g370(.A(new_n562), .B1(KEYINPUT33), .B2(new_n569), .C1(new_n563), .C2(new_n564), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n561), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n563), .A2(new_n564), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT33), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n570), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n565), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n572), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n555), .A2(KEYINPUT70), .A3(new_n559), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n559), .B1(new_n555), .B2(KEYINPUT70), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT29), .B1(new_n444), .B2(new_n447), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n375), .ZN(new_n585));
  NAND2_X1  g384(.A1(G228gat), .A2(G233gat), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(new_n375), .B2(KEYINPUT3), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n502), .B1(new_n381), .B2(new_n382), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n589), .B2(new_n533), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n448), .A2(new_n502), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT88), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n584), .A2(KEYINPUT88), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n594), .A2(new_n380), .A3(new_n595), .ZN(new_n596));
  AOI22_X1  g395(.A1(new_n596), .A2(new_n375), .B1(new_n589), .B2(new_n533), .ZN(new_n597));
  INV_X1    g396(.A(new_n586), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n591), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G78gat), .B(G106gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT31), .B(G50gat), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n600), .B(new_n601), .Z(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT89), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(G22gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n595), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n380), .B1(new_n584), .B2(KEYINPUT88), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n375), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n533), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n590), .B1(new_n610), .B2(new_n586), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n605), .B1(new_n611), .B2(new_n602), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n598), .B1(new_n608), .B2(new_n609), .ZN(new_n613));
  NOR4_X1   g412(.A1(new_n613), .A2(G22gat), .A3(new_n603), .A4(new_n590), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n604), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT89), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(new_n611), .B2(new_n602), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n591), .B(new_n602), .C1(new_n597), .C2(new_n598), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(G22gat), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n611), .A2(new_n605), .A3(new_n602), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n573), .A2(new_n583), .B1(new_n615), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n426), .A2(new_n548), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT35), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n545), .A2(new_n531), .A3(new_n542), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(KEYINPUT35), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n420), .A2(new_n422), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n416), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n425), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n622), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n621), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n425), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT6), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n420), .B2(new_n422), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n421), .B1(new_n420), .B2(new_n422), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n634), .B1(new_n638), .B2(new_n423), .ZN(new_n639));
  INV_X1    g438(.A(new_n547), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n640), .A2(new_n545), .A3(new_n543), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n633), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n383), .A2(new_n388), .A3(new_n393), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n402), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n400), .A2(new_n387), .A3(new_n385), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT39), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT90), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n646), .A2(KEYINPUT90), .A3(KEYINPUT39), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n645), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n644), .A2(new_n652), .A3(new_n402), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n414), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n643), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n645), .A2(new_n649), .A3(new_n650), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n656), .A2(KEYINPUT40), .A3(new_n414), .A4(new_n653), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n627), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n659), .A2(new_n625), .B1(new_n615), .B2(new_n621), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT37), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n537), .A2(new_n661), .A3(new_n538), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n527), .A2(new_n529), .A3(new_n533), .A4(new_n528), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n528), .B1(new_n451), .B2(new_n526), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n521), .B1(new_n664), .B2(KEYINPUT74), .ZN(new_n665));
  OAI211_X1 g464(.A(KEYINPUT37), .B(new_n663), .C1(new_n665), .C2(new_n533), .ZN(new_n666));
  INV_X1    g465(.A(new_n430), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(KEYINPUT38), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n662), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n669), .A2(new_n544), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n662), .A2(new_n539), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n661), .B1(new_n537), .B2(new_n538), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT38), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n670), .A2(new_n425), .A3(new_n673), .A4(new_n628), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n660), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT36), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n571), .A2(new_n561), .A3(new_n572), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n582), .B1(new_n578), .B2(new_n579), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n573), .A2(KEYINPUT36), .A3(new_n583), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n642), .A2(new_n675), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n631), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n343), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n426), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(new_n217), .ZN(G1324gat));
  INV_X1    g486(.A(KEYINPUT42), .ZN(new_n688));
  INV_X1    g487(.A(new_n625), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT16), .B(G8gat), .Z(new_n691));
  AOI21_X1  g490(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G8gat), .B1(new_n685), .B2(new_n689), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT99), .A2(KEYINPUT42), .ZN(new_n694));
  MUX2_X1   g493(.A(KEYINPUT99), .B(new_n694), .S(new_n691), .Z(new_n695));
  AOI22_X1  g494(.A1(new_n692), .A2(new_n693), .B1(new_n690), .B2(new_n695), .ZN(G1325gat));
  OAI21_X1  g495(.A(G15gat), .B1(new_n685), .B2(new_n682), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n573), .A2(new_n583), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n699), .A2(G15gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n697), .B1(new_n685), .B2(new_n700), .ZN(G1326gat));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n632), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT43), .B(G22gat), .Z(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n426), .A2(new_n548), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n681), .B1(new_n706), .B2(new_n633), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n675), .A2(new_n707), .B1(new_n624), .B2(new_n630), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n705), .B1(new_n708), .B2(new_n288), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n642), .A2(new_n675), .A3(new_n682), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n626), .A2(new_n629), .ZN(new_n711));
  AOI22_X1  g510(.A1(KEYINPUT35), .A2(new_n623), .B1(new_n711), .B2(new_n622), .ZN(new_n712));
  OAI211_X1 g511(.A(KEYINPUT44), .B(new_n287), .C1(new_n710), .C2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n330), .A2(new_n335), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n338), .B1(new_n337), .B2(new_n326), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(new_n232), .A3(new_n309), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n709), .A2(new_n639), .A3(new_n713), .A4(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n247), .B1(new_n718), .B2(KEYINPUT100), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT44), .B1(new_n684), .B2(new_n287), .ZN(new_n720));
  AOI211_X1 g519(.A(new_n705), .B(new_n288), .C1(new_n631), .C2(new_n683), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT100), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n722), .A2(new_n723), .A3(new_n639), .A4(new_n717), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n684), .A2(new_n287), .A3(new_n717), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n426), .A2(G29gat), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n725), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT101), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT101), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n725), .A2(new_n734), .A3(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1328gat));
  NOR3_X1   g535(.A1(new_n726), .A2(G36gat), .A3(new_n689), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT46), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n722), .A2(new_n625), .A3(new_n717), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n248), .B2(new_n739), .ZN(G1329gat));
  INV_X1    g539(.A(G43gat), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n709), .A2(new_n681), .A3(new_n713), .A4(new_n717), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT103), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n743), .B2(new_n742), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n708), .A2(new_n288), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n746), .A2(new_n741), .A3(new_n698), .A4(new_n717), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(KEYINPUT47), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n742), .A2(G43gat), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n749), .A2(new_n747), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT102), .B(KEYINPUT47), .Z(new_n751));
  OAI21_X1  g550(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(G1330gat));
  NAND3_X1  g551(.A1(new_n722), .A2(new_n633), .A3(new_n717), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G50gat), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT104), .ZN(new_n755));
  OR3_X1    g554(.A1(new_n726), .A2(G50gat), .A3(new_n632), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n754), .B(new_n756), .C1(KEYINPUT104), .C2(KEYINPUT48), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1331gat));
  NAND3_X1  g560(.A1(new_n232), .A2(new_n288), .A3(new_n309), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n708), .A2(new_n340), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n639), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n625), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT49), .B(G64gat), .Z(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n766), .B2(new_n768), .ZN(G1333gat));
  XNOR2_X1  g568(.A(new_n698), .B(KEYINPUT105), .ZN(new_n770));
  AOI21_X1  g569(.A(G71gat), .B1(new_n763), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n682), .A2(new_n204), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n771), .B1(new_n763), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n773), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g573(.A1(new_n763), .A2(new_n633), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g575(.A1(new_n232), .A2(new_n340), .A3(new_n310), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n722), .A2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778), .B2(new_n426), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n232), .A2(new_n340), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n684), .A2(new_n287), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT106), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT106), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n746), .A2(new_n784), .A3(KEYINPUT51), .A4(new_n780), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(new_n782), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n426), .A2(G85gat), .A3(new_n310), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT107), .Z(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n779), .A2(new_n790), .ZN(G1336gat));
  NOR3_X1   g590(.A1(new_n689), .A2(G92gat), .A3(new_n310), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(KEYINPUT109), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT109), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n787), .A2(new_n795), .A3(new_n792), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n722), .A2(new_n625), .A3(new_n777), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT52), .B1(new_n797), .B2(G92gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n794), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n797), .A2(G92gat), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n781), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT51), .B1(new_n781), .B2(KEYINPUT108), .ZN(new_n802));
  INV_X1    g601(.A(new_n792), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n799), .A2(new_n805), .ZN(G1337gat));
  XNOR2_X1  g605(.A(KEYINPUT110), .B(G99gat), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n787), .A2(new_n698), .A3(new_n309), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n778), .A2(new_n682), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n808), .B1(new_n809), .B2(new_n807), .ZN(G1338gat));
  INV_X1    g609(.A(G106gat), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n709), .A2(new_n633), .A3(new_n713), .A4(new_n777), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(KEYINPUT111), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(KEYINPUT111), .B2(new_n812), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n632), .A2(G106gat), .A3(new_n310), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT53), .B1(new_n787), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n815), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n801), .A2(new_n802), .A3(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n812), .A2(G106gat), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT53), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n821), .ZN(G1339gat));
  OR2_X1    g621(.A1(new_n327), .A2(new_n328), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n320), .B1(new_n319), .B2(new_n322), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(KEYINPUT112), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n826));
  AOI211_X1 g625(.A(new_n826), .B(new_n320), .C1(new_n319), .C2(new_n322), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n334), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n296), .A2(new_n297), .A3(new_n290), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n306), .A2(KEYINPUT54), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n303), .B1(new_n298), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n832), .ZN(new_n836));
  AND3_X1   g635(.A1(new_n835), .A2(new_n308), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n828), .A2(new_n339), .A3(new_n837), .A4(new_n287), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT113), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(new_n308), .A3(new_n836), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n284), .A2(new_n286), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n840), .B1(new_n841), .B2(new_n281), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n842), .A2(new_n843), .A3(new_n339), .A4(new_n828), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n837), .B1(new_n714), .B2(new_n715), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n828), .A2(new_n339), .A3(new_n309), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n287), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT114), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n828), .A2(new_n339), .A3(new_n309), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n840), .B1(new_n336), .B2(new_n339), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n288), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n852), .A2(new_n853), .A3(new_n839), .A4(new_n844), .ZN(new_n854));
  INV_X1    g653(.A(new_n232), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n849), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n311), .A2(new_n340), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n426), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n859), .A2(new_n689), .A3(new_n622), .ZN(new_n860));
  INV_X1    g659(.A(G113gat), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n340), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT116), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n633), .B1(new_n856), .B2(new_n858), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n426), .A2(new_n699), .A3(new_n625), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n865), .A2(KEYINPUT115), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT115), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n867), .A2(new_n868), .A3(new_n716), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n864), .B1(new_n869), .B2(new_n861), .ZN(G1340gat));
  AOI21_X1  g669(.A(G120gat), .B1(new_n860), .B2(new_n309), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n867), .A2(new_n868), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n309), .A2(G120gat), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(G1341gat));
  INV_X1    g673(.A(G127gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n875), .A3(new_n232), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n867), .A2(new_n868), .A3(new_n855), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n875), .ZN(G1342gat));
  NAND2_X1  g677(.A1(new_n689), .A2(new_n287), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(G134gat), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n859), .A2(new_n622), .A3(new_n880), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT56), .Z(new_n882));
  NOR3_X1   g681(.A1(new_n867), .A2(new_n868), .A3(new_n288), .ZN(new_n883));
  INV_X1    g682(.A(G134gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(G1343gat));
  NOR3_X1   g684(.A1(new_n681), .A2(new_n426), .A3(new_n625), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n839), .A2(new_n844), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n840), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n835), .A2(KEYINPUT117), .A3(new_n308), .A4(new_n836), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n847), .B1(new_n716), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n288), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n857), .B1(new_n894), .B2(new_n855), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n632), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT118), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT118), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n232), .B1(new_n887), .B2(new_n893), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n900), .B(new_n897), .C1(new_n901), .C2(new_n857), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n856), .A2(new_n858), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n904), .B2(new_n633), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n340), .B(new_n886), .C1(new_n903), .C2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G141gat), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n682), .A2(new_n633), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n716), .A2(G141gat), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n859), .A2(new_n689), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n912), .A2(KEYINPUT120), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT58), .B1(new_n912), .B2(KEYINPUT120), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n907), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(KEYINPUT119), .ZN(new_n916));
  AOI211_X1 g715(.A(new_n426), .B(new_n908), .C1(new_n856), .C2(new_n858), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n917), .A2(new_n918), .A3(new_n689), .A4(new_n910), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(G141gat), .B2(new_n906), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT58), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n915), .B1(new_n921), .B2(new_n922), .ZN(G1344gat));
  INV_X1    g722(.A(new_n917), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n625), .ZN(new_n925));
  INV_X1    g724(.A(G148gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n925), .A2(new_n926), .A3(new_n309), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT59), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G148gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n886), .B1(new_n903), .B2(new_n905), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n929), .B1(new_n931), .B2(new_n309), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n313), .A2(new_n716), .A3(new_n342), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n232), .B1(new_n893), .B2(new_n838), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n896), .B(new_n633), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n886), .A2(KEYINPUT121), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n886), .A2(KEYINPUT121), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n936), .A2(new_n937), .A3(new_n310), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n632), .B1(new_n856), .B2(new_n858), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n935), .B(new_n938), .C1(new_n939), .C2(new_n896), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n928), .B1(new_n940), .B2(G148gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n927), .B1(new_n932), .B2(new_n941), .ZN(G1345gat));
  OAI21_X1  g741(.A(G155gat), .B1(new_n930), .B2(new_n855), .ZN(new_n943));
  INV_X1    g742(.A(G155gat), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n925), .A2(new_n944), .A3(new_n232), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1346gat));
  OAI21_X1  g745(.A(G162gat), .B1(new_n930), .B2(new_n288), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n879), .A2(G162gat), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n924), .B2(new_n948), .ZN(G1347gat));
  NOR2_X1   g748(.A1(new_n639), .A2(new_n689), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n770), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n865), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(G169gat), .B1(new_n952), .B2(new_n716), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n950), .A2(new_n622), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n954), .B1(new_n856), .B2(new_n858), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n955), .A2(new_n452), .A3(new_n340), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT122), .Z(G1348gat));
  OAI21_X1  g757(.A(G176gat), .B1(new_n952), .B2(new_n310), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n453), .A3(new_n309), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1349gat));
  OAI21_X1  g760(.A(G183gat), .B1(new_n952), .B2(new_n855), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n955), .A2(new_n464), .A3(new_n232), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g764(.A1(new_n865), .A2(new_n287), .A3(new_n951), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT123), .B1(new_n966), .B2(G190gat), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n967), .A2(new_n968), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n466), .A3(new_n287), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(G1351gat));
  NAND2_X1  g773(.A1(new_n950), .A2(new_n682), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n939), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n977), .A2(new_n340), .ZN(new_n978));
  OAI211_X1 g777(.A(new_n935), .B(new_n976), .C1(new_n939), .C2(new_n896), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n340), .A2(G197gat), .ZN(new_n980));
  OAI22_X1  g779(.A1(new_n978), .A2(G197gat), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(new_n981), .ZN(G1352gat));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n310), .A2(G204gat), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n977), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n983), .B1(new_n985), .B2(KEYINPUT62), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n977), .A2(KEYINPUT125), .A3(new_n987), .A4(new_n984), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g788(.A(G204gat), .B1(new_n979), .B2(new_n310), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT124), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n991), .B1(new_n985), .B2(KEYINPUT62), .ZN(new_n992));
  AOI211_X1 g791(.A(KEYINPUT124), .B(new_n987), .C1(new_n977), .C2(new_n984), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n989), .B(new_n990), .C1(new_n992), .C2(new_n993), .ZN(G1353gat));
  INV_X1    g793(.A(G211gat), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n977), .A2(new_n995), .A3(new_n232), .ZN(new_n996));
  INV_X1    g795(.A(new_n979), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n997), .A2(new_n232), .ZN(new_n998));
  AOI21_X1  g797(.A(KEYINPUT63), .B1(new_n998), .B2(G211gat), .ZN(new_n999));
  OAI211_X1 g798(.A(KEYINPUT63), .B(G211gat), .C1(new_n979), .C2(new_n855), .ZN(new_n1000));
  INV_X1    g799(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n996), .B1(new_n999), .B2(new_n1001), .ZN(G1354gat));
  NAND2_X1  g801(.A1(new_n977), .A2(new_n287), .ZN(new_n1003));
  INV_X1    g802(.A(G218gat), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1005), .A2(KEYINPUT126), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT126), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1003), .A2(new_n1007), .A3(new_n1004), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n287), .A2(G218gat), .ZN(new_n1009));
  XOR2_X1   g808(.A(new_n1009), .B(KEYINPUT127), .Z(new_n1010));
  AOI22_X1  g809(.A1(new_n1006), .A2(new_n1008), .B1(new_n997), .B2(new_n1010), .ZN(G1355gat));
endmodule


