

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590;

  INV_X1 U322 ( .A(G78GAT), .ZN(n377) );
  XNOR2_X1 U323 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U324 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U325 ( .A(KEYINPUT119), .B(KEYINPUT55), .ZN(n290) );
  XNOR2_X1 U326 ( .A(n446), .B(n372), .ZN(n374) );
  XNOR2_X1 U327 ( .A(KEYINPUT54), .B(KEYINPUT118), .ZN(n417) );
  XNOR2_X1 U328 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U329 ( .A(n380), .B(n379), .ZN(n382) );
  XNOR2_X1 U330 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n415) );
  XNOR2_X1 U331 ( .A(n416), .B(n415), .ZN(n548) );
  XOR2_X1 U332 ( .A(n450), .B(KEYINPUT120), .Z(n566) );
  XOR2_X1 U333 ( .A(n403), .B(n402), .Z(n575) );
  XNOR2_X1 U334 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U335 ( .A(n454), .B(n453), .ZN(G1349GAT) );
  XOR2_X1 U336 ( .A(G78GAT), .B(G148GAT), .Z(n292) );
  XNOR2_X1 U337 ( .A(G106GAT), .B(G204GAT), .ZN(n291) );
  XNOR2_X1 U338 ( .A(n292), .B(n291), .ZN(n422) );
  XNOR2_X1 U339 ( .A(G176GAT), .B(G92GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n293), .B(G64GAT), .ZN(n342) );
  XNOR2_X1 U341 ( .A(n422), .B(n342), .ZN(n312) );
  INV_X1 U342 ( .A(KEYINPUT13), .ZN(n294) );
  NAND2_X1 U343 ( .A1(KEYINPUT73), .A2(n294), .ZN(n297) );
  INV_X1 U344 ( .A(KEYINPUT73), .ZN(n295) );
  NAND2_X1 U345 ( .A1(n295), .A2(KEYINPUT13), .ZN(n296) );
  NAND2_X1 U346 ( .A1(n297), .A2(n296), .ZN(n299) );
  XNOR2_X1 U347 ( .A(G71GAT), .B(G57GAT), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n373) );
  XOR2_X1 U349 ( .A(n373), .B(KEYINPUT78), .Z(n301) );
  XOR2_X1 U350 ( .A(G99GAT), .B(G85GAT), .Z(n354) );
  XNOR2_X1 U351 ( .A(G120GAT), .B(n354), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U353 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n303) );
  NAND2_X1 U354 ( .A1(G230GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U355 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U356 ( .A(n305), .B(n304), .Z(n310) );
  XOR2_X1 U357 ( .A(KEYINPUT32), .B(KEYINPUT74), .Z(n307) );
  XNOR2_X1 U358 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n308), .B(KEYINPUT31), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U362 ( .A(n312), .B(n311), .ZN(n578) );
  XNOR2_X1 U363 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n313) );
  XNOR2_X1 U364 ( .A(n578), .B(n313), .ZN(n552) );
  XOR2_X1 U365 ( .A(n552), .B(KEYINPUT104), .Z(n538) );
  XOR2_X1 U366 ( .A(G85GAT), .B(G162GAT), .Z(n315) );
  XNOR2_X1 U367 ( .A(G29GAT), .B(G127GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U369 ( .A(KEYINPUT88), .B(G148GAT), .Z(n317) );
  XNOR2_X1 U370 ( .A(G1GAT), .B(G155GAT), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U372 ( .A(n319), .B(n318), .Z(n324) );
  XOR2_X1 U373 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n321) );
  NAND2_X1 U374 ( .A1(G225GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U376 ( .A(KEYINPUT6), .B(n322), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U378 ( .A(KEYINPUT87), .B(KEYINPUT89), .Z(n326) );
  XNOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U381 ( .A(n328), .B(n327), .Z(n334) );
  XOR2_X1 U382 ( .A(G120GAT), .B(KEYINPUT0), .Z(n330) );
  XNOR2_X1 U383 ( .A(G113GAT), .B(G134GAT), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n442) );
  XOR2_X1 U385 ( .A(KEYINPUT3), .B(KEYINPUT86), .Z(n332) );
  XNOR2_X1 U386 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n331) );
  XNOR2_X1 U387 ( .A(n332), .B(n331), .ZN(n420) );
  XNOR2_X1 U388 ( .A(n442), .B(n420), .ZN(n333) );
  XOR2_X1 U389 ( .A(n334), .B(n333), .Z(n505) );
  INV_X1 U390 ( .A(n505), .ZN(n521) );
  XNOR2_X1 U391 ( .A(G8GAT), .B(G183GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n335), .B(G211GAT), .ZN(n376) );
  INV_X1 U393 ( .A(G190GAT), .ZN(n336) );
  NAND2_X1 U394 ( .A1(G36GAT), .A2(n336), .ZN(n339) );
  INV_X1 U395 ( .A(G36GAT), .ZN(n337) );
  NAND2_X1 U396 ( .A1(n337), .A2(G190GAT), .ZN(n338) );
  NAND2_X1 U397 ( .A1(n339), .A2(n338), .ZN(n353) );
  XOR2_X1 U398 ( .A(n353), .B(G204GAT), .Z(n341) );
  NAND2_X1 U399 ( .A1(G226GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U400 ( .A(n341), .B(n340), .ZN(n343) );
  XOR2_X1 U401 ( .A(n343), .B(n342), .Z(n349) );
  XOR2_X1 U402 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n345) );
  XNOR2_X1 U403 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n441) );
  XOR2_X1 U405 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n347) );
  XNOR2_X1 U406 ( .A(G197GAT), .B(G218GAT), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n421) );
  XNOR2_X1 U408 ( .A(n441), .B(n421), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U410 ( .A(n376), .B(n350), .Z(n509) );
  INV_X1 U411 ( .A(n509), .ZN(n525) );
  XOR2_X1 U412 ( .A(KEYINPUT80), .B(KEYINPUT10), .Z(n352) );
  XNOR2_X1 U413 ( .A(G106GAT), .B(G92GAT), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n356) );
  XOR2_X1 U416 ( .A(G134GAT), .B(G218GAT), .Z(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U418 ( .A(n358), .B(n357), .Z(n360) );
  NAND2_X1 U419 ( .A1(G232GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U421 ( .A(n361), .B(KEYINPUT11), .Z(n364) );
  XNOR2_X1 U422 ( .A(G50GAT), .B(KEYINPUT79), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n362), .B(G162GAT), .ZN(n423) );
  XNOR2_X1 U424 ( .A(n423), .B(KEYINPUT9), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n369) );
  XOR2_X1 U426 ( .A(KEYINPUT71), .B(KEYINPUT8), .Z(n366) );
  XNOR2_X1 U427 ( .A(G43GAT), .B(G29GAT), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U429 ( .A(KEYINPUT7), .B(n367), .ZN(n403) );
  INV_X1 U430 ( .A(n403), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n369), .B(n368), .ZN(n408) );
  INV_X1 U432 ( .A(n408), .ZN(n470) );
  XOR2_X1 U433 ( .A(KEYINPUT15), .B(KEYINPUT82), .Z(n371) );
  XNOR2_X1 U434 ( .A(G64GAT), .B(KEYINPUT81), .ZN(n370) );
  XOR2_X1 U435 ( .A(n371), .B(n370), .Z(n384) );
  XOR2_X1 U436 ( .A(G15GAT), .B(G127GAT), .Z(n446) );
  AND2_X1 U437 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U438 ( .A(n375), .B(KEYINPUT12), .ZN(n380) );
  XOR2_X1 U439 ( .A(n376), .B(KEYINPUT14), .Z(n378) );
  XOR2_X1 U440 ( .A(G22GAT), .B(G155GAT), .Z(n429) );
  XNOR2_X1 U441 ( .A(G1GAT), .B(n429), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n556) );
  XOR2_X1 U444 ( .A(KEYINPUT112), .B(n556), .Z(n564) );
  XOR2_X1 U445 ( .A(G197GAT), .B(G141GAT), .Z(n386) );
  XNOR2_X1 U446 ( .A(G15GAT), .B(G22GAT), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U448 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n388) );
  XNOR2_X1 U449 ( .A(G1GAT), .B(G8GAT), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U451 ( .A(n390), .B(n389), .Z(n401) );
  XOR2_X1 U452 ( .A(KEYINPUT29), .B(KEYINPUT72), .Z(n392) );
  XNOR2_X1 U453 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n399) );
  XOR2_X1 U455 ( .A(G113GAT), .B(G36GAT), .Z(n394) );
  XNOR2_X1 U456 ( .A(G169GAT), .B(G50GAT), .ZN(n393) );
  XNOR2_X1 U457 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U458 ( .A(KEYINPUT68), .B(n395), .Z(n397) );
  NAND2_X1 U459 ( .A1(G229GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U460 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U461 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n402) );
  INV_X1 U463 ( .A(n575), .ZN(n503) );
  NOR2_X1 U464 ( .A1(n503), .A2(n552), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n404), .B(KEYINPUT46), .ZN(n405) );
  NOR2_X1 U466 ( .A1(n564), .A2(n405), .ZN(n406) );
  NAND2_X1 U467 ( .A1(n470), .A2(n406), .ZN(n407) );
  XNOR2_X1 U468 ( .A(n407), .B(KEYINPUT47), .ZN(n414) );
  XNOR2_X1 U469 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n410) );
  XOR2_X1 U470 ( .A(n408), .B(KEYINPUT36), .Z(n587) );
  NOR2_X1 U471 ( .A1(n587), .A2(n556), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n412) );
  OR2_X1 U473 ( .A1(n575), .A2(n578), .ZN(n411) );
  NOR2_X1 U474 ( .A1(n412), .A2(n411), .ZN(n413) );
  NOR2_X1 U475 ( .A1(n414), .A2(n413), .ZN(n416) );
  NAND2_X1 U476 ( .A1(n525), .A2(n548), .ZN(n418) );
  NOR2_X1 U477 ( .A1(n521), .A2(n419), .ZN(n573) );
  XOR2_X1 U478 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n433) );
  XOR2_X1 U481 ( .A(G211GAT), .B(KEYINPUT23), .Z(n427) );
  XNOR2_X1 U482 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U484 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n462) );
  AND2_X1 U488 ( .A1(n573), .A2(n462), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n434), .B(n290), .ZN(n449) );
  XOR2_X1 U490 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n436) );
  XNOR2_X1 U491 ( .A(G176GAT), .B(G71GAT), .ZN(n435) );
  XNOR2_X1 U492 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U493 ( .A(G183GAT), .B(G99GAT), .Z(n438) );
  XNOR2_X1 U494 ( .A(G43GAT), .B(G190GAT), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U496 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U499 ( .A(n446), .B(n445), .Z(n448) );
  NAND2_X1 U500 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XOR2_X1 U501 ( .A(n448), .B(n447), .Z(n511) );
  INV_X1 U502 ( .A(n511), .ZN(n534) );
  NAND2_X1 U503 ( .A1(n449), .A2(n534), .ZN(n450) );
  NAND2_X1 U504 ( .A1(n538), .A2(n566), .ZN(n454) );
  XOR2_X1 U505 ( .A(G176GAT), .B(KEYINPUT121), .Z(n452) );
  XOR2_X1 U506 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n451) );
  XOR2_X1 U507 ( .A(KEYINPUT34), .B(KEYINPUT94), .Z(n456) );
  XNOR2_X1 U508 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n475) );
  NOR2_X1 U510 ( .A1(n503), .A2(n578), .ZN(n489) );
  XOR2_X1 U511 ( .A(KEYINPUT27), .B(n509), .Z(n464) );
  AND2_X1 U512 ( .A1(n521), .A2(n464), .ZN(n546) );
  XNOR2_X1 U513 ( .A(KEYINPUT28), .B(KEYINPUT66), .ZN(n457) );
  XOR2_X1 U514 ( .A(n457), .B(n462), .Z(n529) );
  INV_X1 U515 ( .A(n529), .ZN(n515) );
  NAND2_X1 U516 ( .A1(n546), .A2(n515), .ZN(n536) );
  NOR2_X1 U517 ( .A1(n534), .A2(n536), .ZN(n458) );
  XOR2_X1 U518 ( .A(KEYINPUT90), .B(n458), .Z(n469) );
  NAND2_X1 U519 ( .A1(n525), .A2(n534), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n459), .A2(n462), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT25), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n461), .B(KEYINPUT91), .ZN(n466) );
  NOR2_X1 U523 ( .A1(n462), .A2(n534), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT26), .ZN(n572) );
  NAND2_X1 U525 ( .A1(n464), .A2(n572), .ZN(n465) );
  NAND2_X1 U526 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n505), .A2(n467), .ZN(n468) );
  NAND2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n484) );
  NOR2_X1 U529 ( .A1(n408), .A2(n556), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT83), .ZN(n472) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(n472), .Z(n473) );
  AND2_X1 U532 ( .A1(n484), .A2(n473), .ZN(n504) );
  NAND2_X1 U533 ( .A1(n489), .A2(n504), .ZN(n482) );
  NOR2_X1 U534 ( .A1(n505), .A2(n482), .ZN(n474) );
  XOR2_X1 U535 ( .A(n475), .B(n474), .Z(n476) );
  XNOR2_X1 U536 ( .A(KEYINPUT92), .B(n476), .ZN(G1324GAT) );
  NOR2_X1 U537 ( .A1(n509), .A2(n482), .ZN(n477) );
  XOR2_X1 U538 ( .A(G8GAT), .B(n477), .Z(G1325GAT) );
  NOR2_X1 U539 ( .A1(n482), .A2(n511), .ZN(n481) );
  XOR2_X1 U540 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n479) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n478) );
  XNOR2_X1 U542 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NOR2_X1 U544 ( .A1(n515), .A2(n482), .ZN(n483) );
  XOR2_X1 U545 ( .A(G22GAT), .B(n483), .Z(G1327GAT) );
  NAND2_X1 U546 ( .A1(n556), .A2(n484), .ZN(n485) );
  XNOR2_X1 U547 ( .A(KEYINPUT98), .B(n485), .ZN(n486) );
  NOR2_X1 U548 ( .A1(n587), .A2(n486), .ZN(n488) );
  XNOR2_X1 U549 ( .A(KEYINPUT99), .B(KEYINPUT37), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(n518) );
  NAND2_X1 U551 ( .A1(n518), .A2(n489), .ZN(n491) );
  XOR2_X1 U552 ( .A(KEYINPUT100), .B(KEYINPUT38), .Z(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(n501) );
  NAND2_X1 U554 ( .A1(n501), .A2(n521), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT97), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n492), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  XOR2_X1 U558 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n496) );
  NAND2_X1 U559 ( .A1(n501), .A2(n525), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n499) );
  NAND2_X1 U563 ( .A1(n501), .A2(n534), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n500), .ZN(G1330GAT) );
  NAND2_X1 U566 ( .A1(n501), .A2(n529), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n502), .B(G50GAT), .ZN(G1331GAT) );
  AND2_X1 U568 ( .A1(n503), .A2(n538), .ZN(n519) );
  NAND2_X1 U569 ( .A1(n519), .A2(n504), .ZN(n514) );
  NOR2_X1 U570 ( .A1(n505), .A2(n514), .ZN(n507) );
  XNOR2_X1 U571 ( .A(KEYINPUT42), .B(KEYINPUT105), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n508), .ZN(G1332GAT) );
  NOR2_X1 U574 ( .A1(n509), .A2(n514), .ZN(n510) );
  XOR2_X1 U575 ( .A(G64GAT), .B(n510), .Z(G1333GAT) );
  NOR2_X1 U576 ( .A1(n511), .A2(n514), .ZN(n512) );
  XOR2_X1 U577 ( .A(KEYINPUT106), .B(n512), .Z(n513) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(n513), .ZN(G1334GAT) );
  NOR2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n523) );
  NAND2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(KEYINPUT107), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n530), .A2(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n530), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n526), .B(KEYINPUT110), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(n527), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n530), .A2(n534), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n532) );
  NAND2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NAND2_X1 U597 ( .A1(n534), .A2(n548), .ZN(n535) );
  NOR2_X1 U598 ( .A1(n536), .A2(n535), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n575), .A2(n543), .ZN(n537) );
  XNOR2_X1 U600 ( .A(n537), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U602 ( .A1(n543), .A2(n538), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NAND2_X1 U604 ( .A1(n543), .A2(n564), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n541), .B(KEYINPUT50), .ZN(n542) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n542), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U608 ( .A1(n543), .A2(n408), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT114), .ZN(n550) );
  AND2_X1 U611 ( .A1(n546), .A2(n572), .ZN(n547) );
  NAND2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n551) );
  INV_X1 U613 ( .A(n551), .ZN(n560) );
  NAND2_X1 U614 ( .A1(n560), .A2(n575), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1344GAT) );
  NOR2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n554) );
  XNOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n558) );
  INV_X1 U621 ( .A(n556), .ZN(n583) );
  NAND2_X1 U622 ( .A1(n560), .A2(n583), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(n559), .ZN(G1346GAT) );
  XOR2_X1 U625 ( .A(G162GAT), .B(KEYINPUT117), .Z(n562) );
  NAND2_X1 U626 ( .A1(n560), .A2(n408), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n575), .A2(n566), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n566), .A2(n564), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n566), .A2(n408), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n570) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U638 ( .A(KEYINPUT123), .B(n571), .Z(n577) );
  NAND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U640 ( .A(KEYINPUT122), .B(n574), .ZN(n588) );
  INV_X1 U641 ( .A(n588), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n584), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U645 ( .A1(n578), .A2(n584), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n582) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT125), .Z(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  XOR2_X1 U649 ( .A(G211GAT), .B(KEYINPUT127), .Z(n586) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

