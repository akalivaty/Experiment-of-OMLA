//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G107), .ZN(new_n199));
  INV_X1    g013(.A(G107), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G104), .ZN(new_n201));
  OAI21_X1  g015(.A(G101), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT72), .A2(G101), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n198), .A2(G107), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT72), .A2(G101), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT3), .B1(new_n198), .B2(G107), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n200), .A3(G104), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n202), .B1(new_n207), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT1), .B1(new_n213), .B2(G146), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G143), .ZN(new_n217));
  OAI211_X1 g031(.A(G128), .B(new_n214), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(G143), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(G146), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n219), .B(new_n220), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n212), .A2(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT72), .A2(G101), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(new_n203), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n226), .A2(new_n208), .A3(new_n210), .A4(new_n205), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n227), .A2(new_n202), .B1(new_n218), .B2(new_n222), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n197), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT12), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n212), .A2(new_n223), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n227), .A2(new_n222), .A3(new_n218), .A4(new_n202), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n234), .A2(KEYINPUT74), .A3(KEYINPUT12), .A4(new_n197), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n194), .A2(new_n196), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(new_n233), .B2(new_n232), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT74), .B1(new_n238), .B2(KEYINPUT12), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT75), .B1(new_n236), .B2(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(KEYINPUT12), .B(new_n197), .C1(new_n224), .C2(new_n228), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT74), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n243), .A2(new_n231), .A3(new_n244), .A4(new_n235), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n197), .A2(KEYINPUT73), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT73), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n194), .A2(new_n247), .A3(new_n196), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  XNOR2_X1  g064(.A(G143), .B(G146), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n250), .B1(new_n251), .B2(KEYINPUT64), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n219), .A2(new_n220), .ZN(new_n253));
  NOR2_X1   g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT64), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n208), .A2(new_n210), .A3(new_n205), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n227), .A2(KEYINPUT4), .B1(G101), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(KEYINPUT4), .A3(G101), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n258), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT10), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n233), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n223), .ZN(new_n266));
  INV_X1    g080(.A(new_n211), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n201), .A2(new_n225), .A3(new_n203), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n200), .A2(G104), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n205), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n267), .A2(new_n268), .B1(G101), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n266), .A2(new_n271), .A3(KEYINPUT10), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n249), .A2(new_n263), .A3(new_n265), .A4(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G953), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G227), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT71), .ZN(new_n276));
  XNOR2_X1  g090(.A(G110), .B(G140), .ZN(new_n277));
  XOR2_X1   g091(.A(new_n276), .B(new_n277), .Z(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n240), .A2(new_n245), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n272), .A2(new_n265), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n252), .A2(new_n257), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n227), .A2(KEYINPUT4), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n259), .A2(G101), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(new_n286), .B2(new_n261), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n197), .B1(new_n282), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n278), .B1(new_n288), .B2(new_n273), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n281), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n292), .A2(new_n293), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n243), .A2(new_n231), .A3(new_n235), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n278), .B1(new_n297), .B2(new_n273), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n288), .A2(new_n273), .A3(new_n278), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n298), .A2(new_n292), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n294), .A2(new_n296), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT9), .B(G234), .ZN(new_n303));
  OAI21_X1  g117(.A(G221), .B1(new_n303), .B2(G902), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n304), .B(KEYINPUT70), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G214), .B1(G237), .B2(G902), .ZN(new_n308));
  INV_X1    g122(.A(G125), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n252), .B2(new_n257), .ZN(new_n310));
  OR2_X1    g124(.A1(new_n310), .A2(KEYINPUT78), .ZN(new_n311));
  AOI21_X1  g125(.A(G125), .B1(new_n218), .B2(new_n222), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT78), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G224), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G953), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT79), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n311), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n316), .B1(new_n311), .B2(new_n313), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G116), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(G119), .ZN(new_n321));
  AND2_X1   g135(.A1(KEYINPUT65), .A2(G116), .ZN(new_n322));
  NOR2_X1   g136(.A1(KEYINPUT65), .A2(G116), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n321), .B1(new_n324), .B2(G119), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT2), .B(G113), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G119), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n322), .A2(new_n323), .A3(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n326), .B1(new_n330), .B2(new_n321), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n260), .B2(new_n262), .ZN(new_n333));
  OR2_X1    g147(.A1(KEYINPUT65), .A2(G116), .ZN(new_n334));
  NAND2_X1  g148(.A1(KEYINPUT65), .A2(G116), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(G119), .A3(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n336), .B(KEYINPUT5), .C1(new_n320), .C2(G119), .ZN(new_n337));
  INV_X1    g151(.A(G113), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT5), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n329), .A3(G116), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT76), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT76), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n342), .A2(new_n339), .A3(new_n329), .A4(G116), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n338), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n337), .A2(new_n344), .B1(new_n325), .B2(new_n327), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n271), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n333), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G110), .B(G122), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n333), .A2(new_n346), .A3(new_n348), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n350), .A2(KEYINPUT6), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n348), .B1(new_n333), .B2(new_n346), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT6), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n353), .A2(KEYINPUT77), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT77), .B1(new_n353), .B2(new_n354), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n319), .B(new_n352), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(G210), .B1(G237), .B2(G902), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n348), .B(KEYINPUT8), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n345), .A2(new_n271), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n337), .A2(new_n344), .ZN(new_n361));
  AND3_X1   g175(.A1(new_n361), .A2(new_n271), .A3(new_n328), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT7), .B1(new_n314), .B2(G953), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n311), .A2(new_n313), .A3(new_n365), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n364), .B1(new_n310), .B2(new_n312), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n351), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(G902), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n357), .A2(new_n358), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n358), .B1(new_n357), .B2(new_n370), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n308), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n307), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n324), .A2(G122), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n320), .A2(G122), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n200), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n200), .B1(new_n375), .B2(new_n376), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n380));
  OAI22_X1  g194(.A1(new_n380), .A2(KEYINPUT13), .B1(new_n213), .B2(G128), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT13), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(KEYINPUT84), .ZN(new_n383));
  OAI21_X1  g197(.A(G134), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(G128), .B(G143), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g201(.A1(KEYINPUT84), .A2(new_n382), .B1(new_n221), .B2(G143), .ZN(new_n388));
  INV_X1    g202(.A(new_n383), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n385), .B1(new_n390), .B2(G134), .ZN(new_n391));
  OAI22_X1  g205(.A1(new_n378), .A2(new_n379), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n385), .B(new_n188), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n375), .A2(new_n394), .A3(new_n376), .ZN(new_n395));
  OAI21_X1  g209(.A(G107), .B1(new_n375), .B2(new_n394), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n377), .B(new_n393), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G217), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n303), .A2(new_n399), .A3(G953), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n392), .A2(new_n397), .A3(new_n400), .ZN(new_n403));
  AOI21_X1  g217(.A(G902), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G478), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(KEYINPUT15), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G952), .ZN(new_n407));
  AOI211_X1 g221(.A(G953), .B(new_n407), .C1(G234), .C2(G237), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI211_X1 g223(.A(new_n293), .B(new_n274), .C1(G234), .C2(G237), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  XOR2_X1   g225(.A(KEYINPUT21), .B(G898), .Z(new_n412));
  OAI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n403), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n400), .B1(new_n392), .B2(new_n397), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n293), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n405), .A2(KEYINPUT15), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n406), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G113), .B(G122), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(new_n198), .ZN(new_n421));
  INV_X1    g235(.A(G237), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(new_n274), .A3(G214), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n213), .ZN(new_n424));
  NOR2_X1   g238(.A1(G237), .A2(G953), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n425), .A2(G143), .A3(G214), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(KEYINPUT18), .A2(G131), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G140), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G125), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n309), .A2(G140), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n216), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT69), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n431), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n430), .A2(KEYINPUT69), .A3(G125), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n434), .B1(new_n438), .B2(new_n216), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n429), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n436), .A2(KEYINPUT16), .A3(new_n437), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT16), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n431), .A2(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n441), .A2(new_n216), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n216), .B1(new_n441), .B2(new_n443), .ZN(new_n445));
  OAI21_X1  g259(.A(KEYINPUT80), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n441), .A2(new_n443), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G146), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n441), .A2(new_n216), .A3(new_n443), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT80), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n426), .ZN(new_n453));
  AOI21_X1  g267(.A(G143), .B1(new_n425), .B2(G214), .ZN(new_n454));
  OAI21_X1  g268(.A(G131), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n424), .A2(new_n195), .A3(new_n426), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT81), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n427), .A2(KEYINPUT17), .A3(G131), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n455), .A2(KEYINPUT81), .A3(new_n456), .A4(new_n457), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n421), .B(new_n440), .C1(new_n452), .C2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n462), .A2(new_n461), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n466), .A2(new_n446), .A3(new_n451), .A4(new_n460), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n421), .B1(new_n467), .B2(new_n440), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n293), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G475), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n455), .A2(new_n457), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n433), .A2(KEYINPUT19), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n438), .B2(KEYINPUT19), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n448), .B(new_n471), .C1(new_n473), .C2(G146), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n440), .ZN(new_n475));
  INV_X1    g289(.A(new_n421), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n464), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(G475), .A2(G902), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n480), .A2(KEYINPUT82), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT20), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(KEYINPUT82), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n478), .A2(KEYINPUT83), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n480), .B1(new_n464), .B2(new_n477), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n486), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT83), .B1(new_n478), .B2(new_n485), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n419), .B(new_n470), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT85), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n478), .A2(new_n485), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT83), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n478), .A2(new_n479), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT20), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n496), .A3(new_n486), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT85), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n497), .A2(new_n498), .A3(new_n470), .A4(new_n419), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n374), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT32), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n328), .A2(new_n331), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n188), .A2(G137), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n190), .A2(G134), .ZN(new_n505));
  OAI21_X1  g319(.A(G131), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n218), .A2(new_n196), .A3(new_n506), .A4(new_n222), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n237), .B2(new_n283), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT30), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n258), .A2(new_n197), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n507), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n503), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n508), .A2(new_n332), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n425), .A2(G210), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT27), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT26), .B(G101), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NOR4_X1   g333(.A1(new_n513), .A2(KEYINPUT31), .A3(new_n514), .A4(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT28), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n508), .A2(new_n332), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n503), .A2(new_n510), .A3(new_n507), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n196), .A2(new_n506), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n258), .A2(new_n197), .B1(new_n266), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT28), .B1(new_n526), .B2(new_n503), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n519), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT31), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n513), .A2(new_n514), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n518), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n520), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(G472), .A2(G902), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n502), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n503), .B1(new_n510), .B2(new_n507), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT28), .B1(new_n514), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n527), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n518), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n519), .B1(new_n513), .B2(new_n514), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT29), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n293), .B1(new_n540), .B2(new_n542), .ZN(new_n544));
  OAI21_X1  g358(.A(G472), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n513), .A2(new_n514), .A3(new_n519), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n529), .B2(new_n528), .ZN(new_n547));
  OAI211_X1 g361(.A(KEYINPUT32), .B(new_n534), .C1(new_n547), .C2(new_n520), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n536), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT66), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT66), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n536), .A2(new_n545), .A3(new_n548), .A4(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(G234), .ZN(new_n553));
  OAI21_X1  g367(.A(G217), .B1(new_n553), .B2(G902), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT67), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT22), .B(G137), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n274), .A2(G221), .A3(G234), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT24), .B(G110), .Z(new_n561));
  INV_X1    g375(.A(KEYINPUT68), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n221), .A2(G119), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n329), .A2(G128), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n329), .A2(G128), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n221), .A2(G119), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(KEYINPUT68), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n561), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n221), .A2(KEYINPUT23), .A3(G119), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n566), .B(new_n570), .C1(new_n564), .C2(KEYINPUT23), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(G110), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n434), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(new_n445), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n565), .A2(new_n568), .A3(new_n561), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n571), .A2(G110), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n577), .B1(new_n448), .B2(new_n449), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n560), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n448), .B(new_n434), .C1(new_n572), .C2(new_n569), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n575), .B(new_n576), .C1(new_n444), .C2(new_n445), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n559), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n579), .A2(new_n582), .A3(new_n293), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT25), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n579), .A2(new_n582), .A3(KEYINPUT25), .A4(new_n293), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n556), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n579), .A2(new_n582), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n588), .A2(G902), .A3(new_n555), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n550), .A2(new_n552), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n501), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(new_n226), .ZN(G3));
  INV_X1    g407(.A(KEYINPUT88), .ZN(new_n594));
  INV_X1    g408(.A(new_n308), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n357), .A2(new_n370), .ZN(new_n596));
  INV_X1    g410(.A(new_n358), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n357), .A2(new_n358), .A3(new_n370), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n413), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n497), .A2(new_n470), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n293), .A2(G478), .ZN(new_n603));
  OAI21_X1  g417(.A(KEYINPUT33), .B1(new_n414), .B2(new_n415), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n402), .A2(new_n605), .A3(new_n403), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n603), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT87), .B1(new_n404), .B2(G478), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI211_X1 g423(.A(KEYINPUT87), .B(new_n603), .C1(new_n604), .C2(new_n606), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n602), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n594), .B1(new_n601), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT87), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n607), .B2(new_n608), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n497), .B2(new_n470), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n617), .A2(KEYINPUT88), .A3(new_n413), .A4(new_n600), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT86), .ZN(new_n620));
  INV_X1    g434(.A(G472), .ZN(new_n621));
  OAI221_X1 g435(.A(new_n293), .B1(new_n620), .B2(new_n621), .C1(new_n547), .C2(new_n520), .ZN(new_n622));
  OAI211_X1 g436(.A(KEYINPUT86), .B(G472), .C1(new_n533), .C2(G902), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n590), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n307), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(new_n198), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT89), .B(KEYINPUT34), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  INV_X1    g444(.A(new_n601), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n487), .A2(new_n482), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n496), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n470), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n406), .A2(new_n418), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n626), .A2(new_n631), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G107), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT90), .B(KEYINPUT35), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G9));
  NOR2_X1   g455(.A1(new_n555), .A2(G902), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT91), .B1(new_n574), .B2(new_n578), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT91), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n580), .A2(new_n581), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n560), .A2(KEYINPUT36), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n646), .B1(new_n643), .B2(new_n645), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n642), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(KEYINPUT92), .ZN(new_n651));
  INV_X1    g465(.A(new_n587), .ZN(new_n652));
  INV_X1    g466(.A(new_n649), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n647), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT92), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n655), .A3(new_n642), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n651), .A2(new_n652), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n624), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n374), .A2(new_n500), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT37), .B(G110), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT93), .B(KEYINPUT94), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  AOI21_X1  g478(.A(G902), .B1(new_n281), .B2(new_n290), .ZN(new_n665));
  AOI211_X1 g479(.A(new_n295), .B(new_n300), .C1(new_n665), .C2(new_n292), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT95), .B(G900), .Z(new_n667));
  AOI21_X1  g481(.A(new_n408), .B1(new_n410), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n633), .A2(new_n470), .A3(new_n635), .A4(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n666), .A2(new_n670), .A3(new_n305), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n658), .A2(new_n373), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n671), .A2(new_n550), .A3(new_n552), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  NOR2_X1   g488(.A1(new_n371), .A2(new_n372), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n602), .ZN(new_n678));
  NOR4_X1   g492(.A1(new_n677), .A2(new_n678), .A3(new_n636), .A4(new_n595), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n295), .B1(new_n665), .B2(new_n292), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n305), .B1(new_n680), .B2(new_n301), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT97), .B(KEYINPUT39), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n668), .B(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n531), .A2(new_n519), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n522), .A2(new_n523), .A3(new_n519), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n293), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n536), .A2(new_n548), .A3(new_n690), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n691), .A2(new_n658), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n679), .A2(new_n685), .A3(new_n686), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  AOI21_X1  g508(.A(new_n482), .B1(new_n478), .B2(new_n479), .ZN(new_n695));
  AOI211_X1 g509(.A(new_n493), .B(new_n484), .C1(new_n464), .C2(new_n477), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n489), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n470), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n611), .B(new_n669), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n307), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n550), .A3(new_n552), .A4(new_n672), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  AOI21_X1  g516(.A(new_n279), .B1(new_n297), .B2(KEYINPUT75), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n289), .B1(new_n703), .B2(new_n245), .ZN(new_n704));
  OAI21_X1  g518(.A(G469), .B1(new_n704), .B2(G902), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n294), .A2(new_n705), .A3(new_n306), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n550), .A2(new_n552), .A3(new_n590), .A4(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n619), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT41), .B(G113), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NOR3_X1   g526(.A1(new_n601), .A2(new_n636), .A3(new_n634), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  AND4_X1   g529(.A1(new_n550), .A2(new_n500), .A3(new_n552), .A4(new_n657), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n717));
  AOI211_X1 g531(.A(G469), .B(G902), .C1(new_n281), .C2(new_n290), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n600), .A3(KEYINPUT98), .A4(new_n306), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT98), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n294), .A2(new_n705), .A3(new_n306), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n721), .B1(new_n722), .B2(new_n373), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n716), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  NAND2_X1  g540(.A1(new_n706), .A2(new_n413), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT100), .ZN(new_n728));
  INV_X1    g542(.A(new_n589), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n652), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT100), .B1(new_n587), .B2(new_n589), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(G472), .B1(new_n533), .B2(G902), .ZN(new_n733));
  INV_X1    g547(.A(new_n520), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n538), .A2(new_n539), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT31), .B1(new_n735), .B2(new_n519), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n734), .B(KEYINPUT99), .C1(new_n736), .C2(new_n546), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT99), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n547), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n739), .A3(new_n534), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n732), .A2(new_n733), .A3(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n600), .A2(new_n602), .A3(new_n635), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n727), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  XOR2_X1   g557(.A(new_n743), .B(G122), .Z(G24));
  NAND3_X1  g558(.A1(new_n740), .A2(new_n657), .A3(new_n733), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n699), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT98), .B1(new_n706), .B2(new_n600), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n722), .A2(new_n373), .A3(new_n721), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n746), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT101), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n724), .A2(KEYINPUT101), .A3(new_n746), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G125), .ZN(G27));
  NAND4_X1  g568(.A1(new_n549), .A2(new_n617), .A3(new_n669), .A4(new_n732), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT102), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n298), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n299), .B1(new_n298), .B2(new_n756), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(G469), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n680), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n305), .A2(new_n595), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n675), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT42), .B1(new_n755), .B2(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n598), .A2(new_n599), .A3(new_n761), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n680), .B2(new_n759), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n550), .A2(new_n765), .A3(new_n552), .A4(new_n590), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n699), .A2(KEYINPUT42), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n763), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT103), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n763), .B(KEYINPUT103), .C1(new_n766), .C2(new_n767), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G131), .ZN(G33));
  NOR2_X1   g587(.A1(new_n766), .A2(new_n670), .ZN(new_n774));
  XOR2_X1   g588(.A(KEYINPUT104), .B(G134), .Z(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(G36));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n678), .A2(new_n611), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT43), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT105), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n678), .A2(KEYINPUT106), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT106), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n602), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n782), .A2(KEYINPUT43), .A3(new_n611), .A4(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT105), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n778), .A2(new_n786), .A3(new_n779), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n781), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT107), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n658), .B1(new_n622), .B2(new_n623), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n788), .B2(KEYINPUT107), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n777), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n788), .A2(KEYINPUT107), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(KEYINPUT44), .A3(new_n789), .A4(new_n791), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n371), .A2(new_n372), .A3(new_n595), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n298), .A2(new_n299), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT45), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n292), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n757), .A2(KEYINPUT45), .A3(new_n758), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n295), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(KEYINPUT46), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n294), .B1(new_n801), .B2(KEYINPUT46), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n306), .B(new_n683), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n793), .A2(new_n795), .A3(new_n796), .A4(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT108), .B(G137), .Z(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(G39));
  NAND2_X1  g622(.A1(new_n550), .A2(new_n552), .ZN(new_n809));
  INV_X1    g623(.A(new_n699), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n625), .A3(new_n810), .A4(new_n796), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n306), .B1(new_n802), .B2(new_n803), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT47), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(new_n813), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n811), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(new_n430), .ZN(G42));
  NAND2_X1  g631(.A1(new_n719), .A2(KEYINPUT109), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT109), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n717), .B2(new_n718), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  XOR2_X1   g635(.A(new_n821), .B(KEYINPUT49), .Z(new_n822));
  AND3_X1   g636(.A1(new_n782), .A2(new_n611), .A3(new_n784), .ZN(new_n823));
  INV_X1    g637(.A(new_n677), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n732), .A2(new_n761), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n824), .A2(new_n691), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n822), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT116), .B1(new_n788), .B2(new_n408), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n788), .A2(KEYINPUT116), .A3(new_n408), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n741), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n724), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n691), .A2(new_n625), .A3(new_n409), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n706), .A2(new_n796), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n407), .B(G953), .C1(new_n835), .C2(new_n617), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n549), .A2(new_n732), .ZN(new_n837));
  INV_X1    g651(.A(new_n830), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n837), .B(new_n834), .C1(new_n838), .C2(new_n828), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n839), .A2(KEYINPUT48), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(KEYINPUT48), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n832), .B(new_n836), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n824), .A2(new_n308), .A3(new_n722), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n831), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n831), .A2(KEYINPUT50), .A3(new_n843), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n741), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n838), .B2(new_n828), .ZN(new_n850));
  INV_X1    g664(.A(new_n821), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n851), .A2(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(KEYINPUT117), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n305), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n854), .A2(new_n815), .A3(new_n814), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n796), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT51), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n745), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n858), .B(new_n834), .C1(new_n838), .C2(new_n828), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n835), .A2(new_n678), .A3(new_n616), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT120), .Z(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n857), .A2(new_n862), .B1(KEYINPUT119), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n842), .B1(new_n848), .B2(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n846), .A2(KEYINPUT119), .A3(new_n847), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n850), .B2(new_n856), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n831), .A2(KEYINPUT118), .A3(new_n796), .A4(new_n855), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n859), .A4(new_n861), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n865), .B1(new_n871), .B2(new_n863), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n874));
  INV_X1    g688(.A(new_n742), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n305), .B(new_n668), .C1(new_n680), .C2(new_n759), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n692), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n701), .A2(new_n673), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n874), .B1(new_n753), .B2(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n724), .A2(KEYINPUT101), .A3(new_n746), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT101), .B1(new_n724), .B2(new_n746), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n701), .A2(new_n673), .A3(new_n877), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT112), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT112), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n753), .A2(new_n878), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n879), .B1(new_n887), .B2(new_n874), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n716), .A2(new_n724), .B1(new_n707), .B2(new_n713), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n743), .B1(new_n707), .B2(new_n619), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n770), .A2(new_n889), .A3(new_n771), .A4(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n746), .ZN(new_n892));
  OAI22_X1  g706(.A1(new_n766), .A2(new_n670), .B1(new_n892), .B2(new_n762), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n634), .A2(new_n668), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n587), .B1(KEYINPUT92), .B2(new_n650), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n635), .B1(new_n896), .B2(new_n656), .ZN(new_n897));
  AND4_X1   g711(.A1(new_n681), .A2(new_n895), .A3(new_n796), .A4(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(KEYINPUT111), .A3(new_n550), .A4(new_n552), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT111), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n681), .A2(new_n895), .A3(new_n897), .A4(new_n796), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n900), .B1(new_n809), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n591), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n500), .B(new_n374), .C1(new_n904), .C2(new_n659), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT110), .B1(new_n602), .B2(new_n636), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT110), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n497), .A2(new_n907), .A3(new_n470), .A4(new_n635), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n906), .A2(new_n612), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n626), .A2(new_n631), .A3(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n894), .A2(new_n903), .A3(new_n905), .A4(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n891), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT53), .B1(new_n888), .B2(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n753), .A2(new_n878), .A3(new_n885), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n885), .B1(new_n753), .B2(new_n878), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n874), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n884), .A2(KEYINPUT52), .A3(new_n886), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n912), .A3(KEYINPUT53), .A4(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT113), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n913), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n918), .A2(new_n919), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n873), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n916), .A2(new_n917), .A3(new_n912), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT53), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n660), .B1(new_n501), .B2(new_n591), .ZN(new_n926));
  INV_X1    g740(.A(new_n910), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n763), .B(KEYINPUT53), .C1(new_n766), .C2(new_n767), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n928), .A2(new_n930), .A3(new_n903), .A4(new_n894), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n889), .A2(new_n890), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT114), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n889), .A2(KEYINPUT114), .A3(new_n890), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n888), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n925), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(KEYINPUT54), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n872), .A2(new_n922), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(G952), .A2(G953), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n827), .B1(new_n940), .B2(new_n941), .ZN(G75));
  AOI22_X1  g756(.A1(new_n923), .A2(new_n924), .B1(new_n888), .B2(new_n936), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(new_n293), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(G210), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT56), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n352), .B1(new_n355), .B2(new_n356), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(new_n319), .Z(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT55), .Z(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n274), .A2(G952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n950), .B1(new_n945), .B2(new_n946), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(G51));
  XNOR2_X1  g769(.A(new_n943), .B(KEYINPUT54), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n295), .B(KEYINPUT57), .Z(new_n957));
  OAI21_X1  g771(.A(new_n291), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n799), .A2(new_n800), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT121), .Z(new_n960));
  NAND2_X1  g774(.A1(new_n944), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n953), .B1(new_n958), .B2(new_n961), .ZN(G54));
  AND2_X1   g776(.A1(KEYINPUT58), .A2(G475), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n944), .A2(new_n478), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n478), .B1(new_n944), .B2(new_n963), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(new_n953), .ZN(G60));
  INV_X1    g780(.A(new_n953), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n604), .A2(new_n606), .ZN(new_n968));
  NAND2_X1  g782(.A1(G478), .A2(G902), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT59), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n967), .B1(new_n956), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n968), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n970), .B1(new_n922), .B2(new_n939), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(G63));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT122), .ZN(new_n977));
  NAND2_X1  g791(.A1(G217), .A2(G902), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT60), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n938), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT122), .B1(new_n943), .B2(new_n979), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n981), .A2(new_n982), .A3(new_n588), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n967), .ZN(new_n984));
  AOI22_X1  g798(.A1(new_n981), .A2(new_n982), .B1(new_n647), .B2(new_n653), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n976), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n981), .A2(new_n982), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n654), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n988), .A2(KEYINPUT61), .A3(new_n967), .A4(new_n983), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n986), .A2(new_n989), .ZN(G66));
  AOI21_X1  g804(.A(new_n274), .B1(new_n412), .B2(G224), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n928), .A2(new_n890), .A3(new_n889), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n991), .B1(new_n992), .B2(new_n274), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n948), .B1(G898), .B2(new_n274), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n993), .B(new_n994), .Z(G69));
  NAND2_X1  g809(.A1(new_n509), .A2(new_n512), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT123), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(new_n473), .ZN(new_n998));
  INV_X1    g812(.A(new_n772), .ZN(new_n999));
  AND2_X1   g813(.A1(new_n701), .A2(new_n673), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n753), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n837), .A2(new_n875), .ZN(new_n1002));
  OAI22_X1  g816(.A1(new_n804), .A2(new_n1002), .B1(new_n670), .B2(new_n766), .ZN(new_n1003));
  NOR4_X1   g817(.A1(new_n816), .A2(new_n999), .A3(new_n1001), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(G953), .B1(new_n1004), .B2(new_n806), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n274), .A2(G900), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT126), .Z(new_n1007));
  OAI21_X1  g821(.A(new_n998), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1001), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n693), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(KEYINPUT62), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT62), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1009), .A2(new_n1012), .A3(new_n693), .ZN(new_n1013));
  INV_X1    g827(.A(new_n684), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n904), .A2(new_n1014), .A3(new_n796), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n816), .B1(new_n909), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n806), .A2(new_n1011), .A3(new_n1013), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n274), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n998), .B(KEYINPUT124), .ZN(new_n1019));
  AOI21_X1  g833(.A(KEYINPUT125), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT125), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1019), .ZN(new_n1022));
  AOI211_X1 g836(.A(new_n1021), .B(new_n1022), .C1(new_n1017), .C2(new_n274), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1008), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n274), .B1(G227), .B2(G900), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1024), .B(new_n1025), .ZN(G72));
  NAND2_X1  g840(.A1(G472), .A2(G902), .ZN(new_n1027));
  XOR2_X1   g841(.A(new_n1027), .B(KEYINPUT63), .Z(new_n1028));
  NAND2_X1  g842(.A1(new_n1004), .A2(new_n806), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1028), .B1(new_n1029), .B2(new_n992), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1030), .A2(new_n531), .A3(new_n519), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1028), .B1(new_n1017), .B2(new_n992), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(new_n687), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1031), .A2(new_n967), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n920), .A2(new_n921), .ZN(new_n1035));
  INV_X1    g849(.A(new_n687), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n531), .A2(new_n519), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1036), .A2(new_n1037), .A3(new_n1028), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(KEYINPUT127), .Z(new_n1039));
  AOI21_X1  g853(.A(new_n1034), .B1(new_n1035), .B2(new_n1039), .ZN(G57));
endmodule


