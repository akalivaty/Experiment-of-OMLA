//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G43gat), .ZN(new_n204));
  INV_X1    g003(.A(G43gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G50gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT15), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208));
  INV_X1    g007(.A(G29gat), .ZN(new_n209));
  INV_X1    g008(.A(G36gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT86), .ZN(new_n212));
  NOR3_X1   g011(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT86), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(KEYINPUT87), .A2(G29gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(KEYINPUT87), .A2(G29gat), .ZN(new_n219));
  OAI21_X1  g018(.A(G36gat), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n207), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT89), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT15), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n205), .A2(G50gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n203), .A2(G43gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(new_n207), .A3(new_n220), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n216), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT88), .B1(new_n230), .B2(new_n213), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT88), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n211), .A2(new_n232), .A3(new_n216), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n223), .B1(new_n229), .B2(new_n234), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n211), .A2(new_n232), .A3(new_n216), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n232), .B1(new_n211), .B2(new_n216), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NOR3_X1   g037(.A1(new_n238), .A2(new_n228), .A3(KEYINPUT89), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n222), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT90), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G15gat), .B(G22gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT91), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G8gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT16), .ZN(new_n248));
  AOI21_X1  g047(.A(G1gat), .B1(new_n243), .B2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n247), .B(new_n249), .Z(new_n250));
  OAI21_X1  g049(.A(KEYINPUT89), .B1(new_n238), .B2(new_n228), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n220), .A2(new_n207), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n234), .A2(new_n252), .A3(new_n223), .A4(new_n227), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n221), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT90), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n242), .A2(new_n250), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G229gat), .A2(G233gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(new_n253), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT90), .B1(new_n258), .B2(new_n222), .ZN(new_n259));
  AOI211_X1 g058(.A(new_n241), .B(new_n221), .C1(new_n251), .C2(new_n253), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n259), .A2(new_n260), .A3(KEYINPUT17), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(KEYINPUT17), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n247), .B(new_n249), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n256), .B(new_n257), .C1(new_n261), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT18), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT17), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n242), .A2(new_n267), .A3(new_n255), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n262), .A2(new_n263), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n259), .A2(new_n260), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n268), .A2(new_n269), .B1(new_n270), .B2(new_n250), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT18), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n257), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n257), .B(KEYINPUT13), .Z(new_n275));
  AOI21_X1  g074(.A(new_n250), .B1(new_n242), .B2(new_n255), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n259), .A2(new_n260), .A3(new_n263), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT92), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n263), .B1(new_n259), .B2(new_n260), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n256), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(KEYINPUT92), .A3(new_n275), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G113gat), .B(G141gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(G197gat), .ZN(new_n286));
  XOR2_X1   g085(.A(KEYINPUT11), .B(G169gat), .Z(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n288), .B(KEYINPUT12), .Z(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n274), .A2(new_n284), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n290), .B1(new_n274), .B2(new_n284), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n202), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n265), .A2(KEYINPUT18), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n272), .B1(new_n271), .B2(new_n257), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT92), .B1(new_n282), .B2(new_n275), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n282), .A2(KEYINPUT92), .A3(new_n275), .ZN(new_n297));
  OAI22_X1  g096(.A1(new_n294), .A2(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n289), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n274), .A2(new_n284), .A3(new_n290), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n299), .A2(KEYINPUT93), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n293), .A2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(KEYINPUT68), .B(KEYINPUT36), .Z(new_n303));
  OR2_X1    g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(KEYINPUT24), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(KEYINPUT24), .B2(new_n305), .ZN(new_n307));
  NOR2_X1   g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(G169gat), .B2(G176gat), .ZN(new_n311));
  INV_X1    g110(.A(G169gat), .ZN(new_n312));
  INV_X1    g111(.A(G176gat), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n309), .B(new_n311), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT25), .B1(new_n314), .B2(KEYINPUT64), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT27), .B(G183gat), .ZN(new_n318));
  INV_X1    g117(.A(G190gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(new_n320), .B(KEYINPUT28), .Z(new_n321));
  INV_X1    g120(.A(new_n305), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n312), .A2(new_n313), .ZN(new_n323));
  NOR3_X1   g122(.A1(new_n323), .A2(KEYINPUT26), .A3(new_n308), .ZN(new_n324));
  AOI211_X1 g123(.A(new_n322), .B(new_n324), .C1(KEYINPUT26), .C2(new_n308), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n317), .A2(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(KEYINPUT66), .B(G113gat), .Z(new_n328));
  INV_X1    g127(.A(G120gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(KEYINPUT65), .B(G120gat), .ZN(new_n330));
  INV_X1    g129(.A(G113gat), .ZN(new_n331));
  OAI22_X1  g130(.A1(new_n328), .A2(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT1), .ZN(new_n333));
  XNOR2_X1  g132(.A(G127gat), .B(G134gat), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G113gat), .A2(G120gat), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT1), .B1(new_n331), .B2(new_n329), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n327), .A2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n339), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n317), .A2(new_n341), .A3(new_n326), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT34), .ZN(new_n344));
  INV_X1    g143(.A(G227gat), .ZN(new_n345));
  INV_X1    g144(.A(G233gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n343), .A2(new_n344), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n342), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n341), .B1(new_n317), .B2(new_n326), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT34), .B1(new_n352), .B2(new_n347), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT33), .B1(new_n352), .B2(new_n347), .ZN(new_n354));
  XNOR2_X1  g153(.A(G15gat), .B(G43gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(G71gat), .B(G99gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n355), .B(new_n356), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n349), .B(new_n353), .C1(new_n354), .C2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n347), .A3(new_n342), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT32), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT33), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n357), .B1(new_n359), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n344), .B1(new_n343), .B2(new_n348), .ZN(new_n364));
  AOI211_X1 g163(.A(KEYINPUT34), .B(new_n347), .C1(new_n340), .C2(new_n342), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n358), .A2(new_n361), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n361), .B1(new_n358), .B2(new_n366), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n303), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT69), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT69), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n371), .B(new_n303), .C1(new_n367), .C2(new_n368), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n366), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n360), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n358), .A2(new_n361), .A3(new_n366), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(KEYINPUT36), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT67), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n376), .A2(KEYINPUT67), .A3(KEYINPUT36), .A4(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n373), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT5), .ZN(new_n384));
  INV_X1    g183(.A(G141gat), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT74), .B1(new_n385), .B2(G148gat), .ZN(new_n386));
  OR3_X1    g185(.A1(new_n385), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n387));
  XOR2_X1   g186(.A(KEYINPUT73), .B(G141gat), .Z(new_n388));
  INV_X1    g187(.A(G148gat), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT75), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(G155gat), .A2(G162gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n394), .A2(KEYINPUT2), .ZN(new_n395));
  INV_X1    g194(.A(G155gat), .ZN(new_n396));
  INV_X1    g195(.A(G162gat), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n392), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G141gat), .B(G148gat), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n399), .B(new_n394), .C1(new_n402), .C2(KEYINPUT2), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n341), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(new_n403), .A3(new_n339), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n384), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT4), .ZN(new_n411));
  OR2_X1    g210(.A1(new_n390), .A2(new_n391), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n391), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n412), .A2(new_n413), .B1(new_n399), .B2(new_n395), .ZN(new_n414));
  INV_X1    g213(.A(new_n403), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n411), .B1(new_n416), .B2(new_n339), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n406), .A2(KEYINPUT4), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n408), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT3), .B1(new_n414), .B2(new_n415), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n341), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT76), .B1(new_n404), .B2(KEYINPUT3), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT76), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT3), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n416), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n421), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n410), .B1(new_n419), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n423), .B1(new_n416), .B2(new_n424), .ZN(new_n428));
  NOR4_X1   g227(.A1(new_n414), .A2(KEYINPUT76), .A3(KEYINPUT3), .A4(new_n415), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n341), .B(new_n420), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT77), .B1(new_n406), .B2(KEYINPUT4), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n406), .A2(KEYINPUT4), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT77), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n416), .A2(new_n433), .A3(new_n411), .A4(new_n339), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n430), .A2(new_n435), .A3(new_n384), .A4(new_n408), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n427), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G1gat), .B(G29gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT0), .ZN(new_n439));
  XNOR2_X1  g238(.A(G57gat), .B(G85gat), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n439), .B(new_n440), .Z(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AND4_X1   g241(.A1(KEYINPUT84), .A2(new_n437), .A3(KEYINPUT6), .A4(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n441), .B1(new_n427), .B2(new_n436), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT84), .B1(new_n444), .B2(KEYINPUT6), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g245(.A(new_n441), .B(KEYINPUT80), .Z(new_n447));
  INV_X1    g246(.A(KEYINPUT82), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n427), .A2(new_n436), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n448), .B1(new_n427), .B2(new_n436), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n427), .A2(new_n436), .A3(new_n441), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g254(.A(KEYINPUT83), .B(KEYINPUT38), .ZN(new_n456));
  XNOR2_X1  g255(.A(G8gat), .B(G36gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(G64gat), .B(G92gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n457), .B(new_n458), .Z(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G197gat), .B(G204gat), .ZN(new_n461));
  INV_X1    g260(.A(G211gat), .ZN(new_n462));
  INV_X1    g261(.A(G218gat), .ZN(new_n463));
  OAI22_X1  g262(.A1(new_n462), .A2(new_n463), .B1(KEYINPUT70), .B2(KEYINPUT22), .ZN(new_n464));
  AND2_X1   g263(.A1(KEYINPUT70), .A2(KEYINPUT22), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(G211gat), .B(G218gat), .Z(new_n467));
  AND2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n466), .A2(new_n467), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G226gat), .A2(G233gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n471), .B(KEYINPUT71), .Z(new_n472));
  INV_X1    g271(.A(KEYINPUT29), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n472), .B1(new_n327), .B2(new_n473), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n315), .A2(new_n316), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n315), .A2(new_n316), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n475), .A2(new_n476), .B1(new_n321), .B2(new_n325), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n477), .A2(new_n471), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n470), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n471), .B1(new_n477), .B2(KEYINPUT29), .ZN(new_n480));
  INV_X1    g279(.A(new_n470), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n327), .A2(new_n472), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n460), .B1(new_n484), .B2(KEYINPUT37), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(KEYINPUT37), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n456), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n479), .A2(new_n483), .A3(new_n459), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n481), .B1(new_n474), .B2(new_n478), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n480), .A2(new_n470), .A3(new_n482), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(KEYINPUT37), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n456), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n489), .B1(new_n485), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n446), .A2(new_n455), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT3), .B1(new_n481), .B2(new_n473), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n416), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n473), .B1(new_n428), .B2(new_n429), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(new_n470), .ZN(new_n500));
  NAND2_X1  g299(.A1(G228gat), .A2(G233gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n422), .A2(new_n425), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n481), .B1(new_n502), .B2(new_n473), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n470), .A2(KEYINPUT78), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT78), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT29), .B1(new_n468), .B2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n504), .B(new_n506), .C1(new_n414), .C2(new_n415), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n507), .A2(KEYINPUT79), .A3(new_n420), .ZN(new_n508));
  AOI21_X1  g307(.A(KEYINPUT79), .B1(new_n507), .B2(new_n420), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n501), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  OAI22_X1  g309(.A1(new_n500), .A2(new_n501), .B1(new_n503), .B2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT31), .B(G50gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n512), .ZN(new_n514));
  OAI221_X1 g313(.A(new_n514), .B1(new_n503), .B2(new_n510), .C1(new_n500), .C2(new_n501), .ZN(new_n515));
  XNOR2_X1  g314(.A(G78gat), .B(G106gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(G22gat), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n513), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n513), .B2(new_n515), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n408), .B1(new_n430), .B2(new_n435), .ZN(new_n521));
  OAI211_X1 g320(.A(KEYINPUT81), .B(KEYINPUT39), .C1(new_n407), .C2(new_n409), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT39), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n447), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT81), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT40), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n523), .B(KEYINPUT40), .C1(new_n525), .C2(new_n526), .ZN(new_n530));
  INV_X1    g329(.A(new_n483), .ZN(new_n531));
  INV_X1    g330(.A(new_n472), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(new_n477), .B2(KEYINPUT29), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n327), .A2(G226gat), .A3(G233gat), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n481), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n460), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n479), .A2(KEYINPUT30), .A3(new_n483), .A4(new_n459), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n489), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n529), .A2(new_n530), .A3(new_n451), .A4(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n496), .A2(new_n520), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT72), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT72), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n547), .A3(new_n541), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n437), .A2(new_n442), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(new_n453), .A3(new_n452), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n444), .A2(KEYINPUT6), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n383), .B(new_n544), .C1(new_n520), .C2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n519), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n513), .A2(new_n515), .A3(new_n517), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n367), .A2(new_n368), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n550), .A2(new_n551), .ZN(new_n558));
  INV_X1    g357(.A(new_n548), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT35), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n446), .A2(new_n455), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT85), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n563), .B1(new_n367), .B2(new_n368), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n376), .A2(KEYINPUT85), .A3(new_n377), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n542), .A2(KEYINPUT35), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n562), .A2(new_n520), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n302), .B1(new_n553), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT100), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  OR2_X1    g371(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n573));
  INV_X1    g372(.A(G85gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(KEYINPUT98), .A2(G92gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT8), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(G92gat), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT7), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT7), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(G85gat), .A3(G92gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n572), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n584), .A2(new_n572), .A3(new_n576), .A4(new_n578), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n584), .A2(new_n576), .A3(new_n578), .ZN(new_n590));
  INV_X1    g389(.A(new_n572), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(KEYINPUT99), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n571), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(new_n591), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(new_n587), .A3(new_n586), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(KEYINPUT100), .A3(new_n592), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n268), .A2(new_n262), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI22_X1  g401(.A1(new_n270), .A2(new_n598), .B1(KEYINPUT41), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G190gat), .B(G218gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n600), .A2(new_n603), .A3(new_n605), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(KEYINPUT97), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT101), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n607), .A2(new_n611), .A3(new_n608), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n602), .A2(KEYINPUT41), .ZN(new_n613));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n609), .A2(KEYINPUT101), .A3(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  OR2_X1    g420(.A1(G71gat), .A2(G78gat), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT9), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(G57gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(G64gat), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(G64gat), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n627), .B2(KEYINPUT94), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT94), .ZN(new_n629));
  NOR3_X1   g428(.A1(new_n629), .A2(new_n625), .A3(G64gat), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n624), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(G64gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(G57gat), .ZN(new_n633));
  OAI21_X1  g432(.A(KEYINPUT9), .B1(new_n627), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n621), .A3(new_n622), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT21), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT95), .ZN(new_n639));
  XNOR2_X1  g438(.A(G127gat), .B(G155gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n640), .B(KEYINPUT96), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g441(.A(G183gat), .B(G211gat), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n263), .B1(new_n637), .B2(new_n636), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n646));
  NAND2_X1  g445(.A1(G231gat), .A2(G233gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n645), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n644), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n620), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n636), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(new_n594), .B2(new_n597), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n596), .A2(new_n636), .A3(new_n592), .ZN(new_n661));
  INV_X1    g460(.A(new_n636), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(new_n595), .A3(new_n586), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n661), .A2(new_n663), .A3(new_n657), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n656), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n656), .B1(new_n661), .B2(new_n663), .ZN(new_n667));
  XNOR2_X1  g466(.A(G120gat), .B(G148gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(G176gat), .B(G204gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  OR3_X1    g470(.A1(new_n666), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n666), .B2(new_n667), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n655), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n570), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n558), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g479(.A(new_n246), .B1(new_n677), .B2(new_n542), .ZN(new_n681));
  INV_X1    g480(.A(new_n542), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT16), .B(G8gat), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n676), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT42), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(KEYINPUT42), .B2(new_n684), .ZN(G1325gat));
  AOI21_X1  g485(.A(G15gat), .B1(new_n677), .B2(new_n566), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT102), .ZN(new_n688));
  INV_X1    g487(.A(new_n383), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n689), .A2(G15gat), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n688), .B1(new_n677), .B2(new_n690), .ZN(G1326gat));
  NAND2_X1  g490(.A1(new_n554), .A2(new_n555), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT103), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT43), .B(G22gat), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n694), .B(new_n696), .ZN(G1327gat));
  INV_X1    g496(.A(new_n674), .ZN(new_n698));
  AND4_X1   g497(.A1(new_n570), .A2(new_n653), .A3(new_n619), .A4(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n218), .A2(new_n219), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n699), .A2(new_n678), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT45), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n383), .A2(new_n544), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT105), .B1(new_n520), .B2(new_n552), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n692), .A2(new_n560), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n569), .B1(new_n703), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n619), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n553), .A2(new_n569), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(KEYINPUT44), .A3(new_n619), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n674), .B(KEYINPUT104), .Z(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n291), .A2(new_n292), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n715), .A2(new_n716), .A3(new_n654), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n711), .A2(new_n713), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT106), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n711), .A2(new_n720), .A3(new_n713), .A4(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n558), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n702), .B1(new_n723), .B2(new_n700), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n699), .A2(new_n210), .A3(new_n542), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT46), .Z(new_n726));
  OAI21_X1  g525(.A(G36gat), .B1(new_n722), .B2(new_n682), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(G1329gat));
  OAI21_X1  g527(.A(G43gat), .B1(new_n718), .B2(new_n383), .ZN(new_n729));
  INV_X1    g528(.A(new_n566), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(G43gat), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n699), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n729), .A2(KEYINPUT47), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n719), .A2(new_n689), .A3(new_n721), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n734), .A2(G43gat), .B1(new_n699), .B2(new_n731), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n735), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g535(.A(KEYINPUT48), .B(G50gat), .C1(new_n718), .C2(new_n520), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n699), .A2(new_n203), .A3(new_n692), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n737), .B(new_n738), .C1(KEYINPUT107), .C2(KEYINPUT48), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(KEYINPUT107), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n719), .A2(new_n692), .A3(new_n721), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n741), .B2(G50gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n742), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g542(.A(new_n716), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n655), .A2(new_n744), .A3(new_n714), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n708), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n678), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n542), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n752));
  XOR2_X1   g551(.A(KEYINPUT49), .B(G64gat), .Z(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n751), .B2(new_n753), .ZN(G1333gat));
  NAND2_X1  g553(.A1(new_n748), .A2(new_n689), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n730), .A2(G71gat), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n755), .A2(G71gat), .B1(new_n748), .B2(new_n756), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g557(.A1(new_n748), .A2(new_n692), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT109), .B(G78gat), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1335gat));
  NOR3_X1   g560(.A1(new_n744), .A2(new_n654), .A3(new_n698), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n711), .A2(new_n713), .A3(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(G85gat), .B1(new_n763), .B2(new_n558), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n744), .A2(new_n654), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n708), .A2(new_n619), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n708), .A2(KEYINPUT51), .A3(new_n619), .A4(new_n765), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n678), .A2(new_n574), .A3(new_n674), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n764), .B1(new_n770), .B2(new_n771), .ZN(G1336gat));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n768), .A2(new_n773), .A3(new_n769), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n766), .A2(KEYINPUT110), .A3(new_n767), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n714), .A2(new_n682), .A3(G92gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n774), .A2(KEYINPUT111), .A3(new_n775), .A4(new_n776), .ZN(new_n780));
  INV_X1    g579(.A(new_n573), .ZN(new_n781));
  INV_X1    g580(.A(new_n575), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n763), .A2(new_n682), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT52), .ZN(new_n785));
  INV_X1    g584(.A(new_n770), .ZN(new_n786));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(new_n786), .B2(new_n776), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n783), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(G1337gat));
  OAI21_X1  g588(.A(G99gat), .B1(new_n763), .B2(new_n383), .ZN(new_n790));
  OR3_X1    g589(.A1(new_n730), .A2(G99gat), .A3(new_n698), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n770), .B2(new_n791), .ZN(G1338gat));
  OAI21_X1  g591(.A(G106gat), .B1(new_n763), .B2(new_n520), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n520), .A2(G106gat), .A3(new_n714), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n774), .A2(new_n775), .A3(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(KEYINPUT112), .B(G106gat), .C1(new_n763), .C2(new_n520), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n795), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT53), .B1(new_n786), .B2(new_n796), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n793), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1339gat));
  OAI22_X1  g602(.A1(new_n271), .A2(new_n257), .B1(new_n282), .B2(new_n275), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n288), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n300), .A2(new_n674), .A3(new_n805), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n596), .A2(KEYINPUT100), .A3(new_n592), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT100), .B1(new_n596), .B2(new_n592), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n658), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n661), .A2(new_n663), .A3(new_n657), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n812), .A3(new_n656), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n813), .A2(KEYINPUT55), .A3(new_n671), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n811), .B2(new_n656), .ZN(new_n815));
  INV_X1    g614(.A(new_n656), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n809), .A2(new_n810), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT113), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  AND4_X1   g617(.A1(KEYINPUT113), .A2(new_n665), .A3(KEYINPUT54), .A4(new_n817), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n814), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n813), .A2(new_n671), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n665), .A2(KEYINPUT54), .A3(new_n817), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n815), .A2(KEYINPUT113), .A3(new_n817), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n820), .B(new_n672), .C1(new_n826), .C2(KEYINPUT55), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n806), .B1(new_n716), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n620), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n300), .A2(new_n805), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n617), .B2(new_n618), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n820), .A2(new_n672), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n824), .A2(new_n825), .ZN(new_n833));
  INV_X1    g632(.A(new_n821), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT55), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n654), .B1(new_n829), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n620), .A2(new_n716), .A3(new_n654), .A4(new_n698), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT114), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n828), .A2(new_n620), .B1(new_n831), .B2(new_n836), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n842), .B(new_n839), .C1(new_n843), .C2(new_n654), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n678), .A2(new_n682), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n730), .A2(new_n692), .ZN(new_n849));
  INV_X1    g648(.A(new_n302), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n848), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(KEYINPUT115), .A3(G113gat), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT115), .B1(new_n851), .B2(G113gat), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n848), .A2(new_n520), .A3(new_n556), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n716), .A2(new_n328), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT116), .ZN(new_n857));
  OAI22_X1  g656(.A1(new_n853), .A2(new_n854), .B1(new_n855), .B2(new_n857), .ZN(G1340gat));
  OR3_X1    g657(.A1(new_n855), .A2(new_n330), .A3(new_n698), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n848), .A2(new_n849), .A3(new_n715), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n861), .A3(G120gat), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n861), .B1(new_n860), .B2(G120gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(G1341gat));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n849), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n654), .A2(G127gat), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT118), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n855), .A2(new_n653), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n869), .B2(G127gat), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n866), .A2(KEYINPUT118), .A3(new_n867), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(G1342gat));
  AND2_X1   g671(.A1(new_n845), .A2(new_n678), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n620), .A2(new_n542), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n557), .A2(G134gat), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  XOR2_X1   g675(.A(new_n876), .B(KEYINPUT56), .Z(new_n877));
  OAI21_X1  g676(.A(G134gat), .B1(new_n866), .B2(new_n620), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1343gat));
  NAND3_X1  g678(.A1(new_n841), .A2(new_n692), .A3(new_n844), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT57), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n293), .A2(new_n301), .A3(new_n836), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n619), .B1(new_n883), .B2(new_n806), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n831), .A2(new_n836), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n653), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n839), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n520), .A2(new_n881), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT119), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n882), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n383), .A2(new_n847), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n388), .B1(new_n896), .B2(new_n302), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n689), .A2(new_n520), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n302), .A2(G141gat), .ZN(new_n900));
  AND4_X1   g699(.A1(new_n847), .A2(new_n845), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n897), .A2(new_n898), .A3(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n891), .B1(new_n887), .B2(new_n888), .ZN(new_n905));
  INV_X1    g704(.A(new_n888), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT119), .B(new_n906), .C1(new_n886), .C2(new_n839), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  AOI211_X1 g707(.A(new_n716), .B(new_n894), .C1(new_n908), .C2(new_n882), .ZN(new_n909));
  INV_X1    g708(.A(new_n388), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n902), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n904), .B1(new_n911), .B2(KEYINPUT58), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n893), .A2(new_n744), .A3(new_n895), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n901), .B1(new_n913), .B2(new_n388), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n914), .A2(KEYINPUT120), .A3(new_n898), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n903), .B1(new_n912), .B2(new_n915), .ZN(G1344gat));
  AND2_X1   g715(.A1(new_n848), .A2(new_n899), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n917), .A2(new_n389), .A3(new_n674), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n895), .A2(new_n674), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n675), .A2(new_n302), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n886), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT57), .B1(new_n922), .B2(new_n692), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n841), .A2(new_n844), .A3(new_n888), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n923), .B1(KEYINPUT122), .B2(new_n924), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(KEYINPUT122), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n927), .A2(KEYINPUT123), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n389), .B1(new_n927), .B2(KEYINPUT123), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n919), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n893), .A2(new_n674), .A3(new_n895), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n389), .A2(KEYINPUT59), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n931), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n918), .B1(new_n930), .B2(new_n936), .ZN(G1345gat));
  NAND3_X1  g736(.A1(new_n917), .A2(new_n396), .A3(new_n654), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n896), .A2(new_n653), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n396), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g741(.A(new_n938), .B(KEYINPUT124), .C1(new_n939), .C2(new_n396), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1346gat));
  OAI21_X1  g743(.A(G162gat), .B1(new_n896), .B2(new_n620), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n873), .A2(new_n397), .A3(new_n874), .A4(new_n899), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1347gat));
  NOR2_X1   g746(.A1(new_n678), .A2(new_n682), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n841), .A2(new_n844), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n849), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n950), .A2(new_n312), .A3(new_n302), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n949), .A2(new_n520), .A3(new_n556), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n744), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n953), .B2(new_n312), .ZN(G1348gat));
  NAND3_X1  g753(.A1(new_n952), .A2(new_n313), .A3(new_n674), .ZN(new_n955));
  OAI21_X1  g754(.A(G176gat), .B1(new_n950), .B2(new_n714), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1349gat));
  NAND3_X1  g756(.A1(new_n952), .A2(new_n318), .A3(new_n654), .ZN(new_n958));
  OAI21_X1  g757(.A(G183gat), .B1(new_n950), .B2(new_n653), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n961));
  XOR2_X1   g760(.A(new_n960), .B(new_n961), .Z(G1350gat));
  NAND3_X1  g761(.A1(new_n952), .A2(new_n319), .A3(new_n619), .ZN(new_n963));
  OAI21_X1  g762(.A(G190gat), .B1(new_n950), .B2(new_n620), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n964), .A2(KEYINPUT61), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n964), .A2(KEYINPUT61), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(G1351gat));
  INV_X1    g767(.A(G197gat), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n383), .A2(new_n948), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n970), .B1(new_n925), .B2(new_n926), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n971), .B2(new_n850), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT127), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n949), .A2(new_n899), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n744), .A2(new_n969), .ZN(new_n976));
  OR3_X1    g775(.A1(new_n975), .A2(KEYINPUT126), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(KEYINPUT126), .B1(new_n975), .B2(new_n976), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n973), .A2(new_n974), .A3(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n979), .ZN(new_n981));
  OAI21_X1  g780(.A(KEYINPUT127), .B1(new_n981), .B2(new_n972), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n982), .ZN(G1352gat));
  INV_X1    g782(.A(new_n971), .ZN(new_n984));
  OAI21_X1  g783(.A(G204gat), .B1(new_n984), .B2(new_n714), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n698), .A2(G204gat), .ZN(new_n986));
  OAI21_X1  g785(.A(KEYINPUT62), .B1(new_n975), .B2(new_n986), .ZN(new_n987));
  OR3_X1    g786(.A1(new_n975), .A2(KEYINPUT62), .A3(new_n986), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(G1353gat));
  INV_X1    g788(.A(new_n975), .ZN(new_n990));
  NAND3_X1  g789(.A1(new_n990), .A2(new_n462), .A3(new_n654), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n971), .A2(new_n654), .ZN(new_n992));
  AND3_X1   g791(.A1(new_n992), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n993));
  AOI21_X1  g792(.A(KEYINPUT63), .B1(new_n992), .B2(G211gat), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n991), .B1(new_n993), .B2(new_n994), .ZN(G1354gat));
  OAI21_X1  g794(.A(G218gat), .B1(new_n984), .B2(new_n620), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n990), .A2(new_n463), .A3(new_n619), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(G1355gat));
endmodule


