//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  INV_X1    g000(.A(G134), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G137), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT66), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n187), .A2(KEYINPUT66), .A3(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(KEYINPUT1), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(KEYINPUT1), .A3(G146), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n202), .B(new_n203), .C1(G128), .C2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT11), .B1(new_n187), .B2(G137), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT11), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(new_n191), .A3(G134), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(new_n188), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n195), .A2(new_n205), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n191), .A2(G134), .ZN(new_n215));
  AOI211_X1 g029(.A(G131), .B(new_n215), .C1(new_n206), .C2(new_n208), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n210), .B1(new_n209), .B2(new_n188), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n207), .B1(G134), .B2(new_n191), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n187), .A2(KEYINPUT11), .A3(G137), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n188), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G131), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(KEYINPUT68), .A3(new_n211), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(KEYINPUT0), .A2(G128), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n199), .A2(new_n201), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT0), .B(G128), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n226), .B(new_n227), .C1(new_n204), .C2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n199), .A2(new_n201), .ZN(new_n230));
  INV_X1    g044(.A(new_n225), .ZN(new_n231));
  OR2_X1    g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n230), .A2(KEYINPUT65), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n213), .B1(new_n224), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT67), .B(G119), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G116), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(G116), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n236), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n242), .B1(new_n246), .B2(new_n240), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n235), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G237), .A2(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G210), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(KEYINPUT27), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(G101), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  AND2_X1   g071(.A1(new_n229), .A2(new_n233), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n218), .B2(new_n223), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT30), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n259), .A2(new_n260), .A3(new_n213), .ZN(new_n261));
  XOR2_X1   g075(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n222), .A2(new_n211), .B1(new_n229), .B2(new_n233), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n263), .B1(new_n213), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n248), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n261), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n224), .A2(new_n234), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT30), .A3(new_n212), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n222), .A2(new_n211), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n234), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n212), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n249), .B1(new_n273), .B2(new_n263), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT69), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n257), .B1(new_n268), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n255), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n273), .A2(new_n248), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(new_n235), .B2(new_n249), .ZN(new_n280));
  NOR4_X1   g094(.A1(new_n259), .A2(KEYINPUT28), .A3(new_n213), .A4(new_n248), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n276), .A2(KEYINPUT31), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT31), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n257), .B(new_n284), .C1(new_n268), .C2(new_n275), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT70), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT70), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n267), .B1(new_n261), .B2(new_n266), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n270), .A2(new_n274), .A3(KEYINPUT69), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n256), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n287), .B1(new_n290), .B2(new_n284), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n283), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(G472), .A2(G902), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(KEYINPUT32), .A3(new_n293), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n250), .B(new_n277), .C1(new_n268), .C2(new_n275), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n282), .A2(new_n255), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT29), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n248), .B1(new_n259), .B2(new_n213), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n299), .B1(new_n280), .B2(new_n281), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n255), .A2(KEYINPUT29), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G472), .B1(new_n297), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT72), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(KEYINPUT72), .B(G472), .C1(new_n297), .C2(new_n302), .ZN(new_n306));
  AND3_X1   g120(.A1(new_n294), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n282), .A2(new_n277), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(new_n290), .B2(new_n284), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n290), .A2(new_n287), .A3(new_n284), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n285), .A2(KEYINPUT70), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n293), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n308), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n292), .A2(KEYINPUT71), .A3(new_n293), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT32), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n307), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  INV_X1    g134(.A(G953), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G214), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n200), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n251), .A2(G143), .A3(G214), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(KEYINPUT18), .A2(G131), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G125), .B(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n198), .ZN(new_n329));
  NOR2_X1   g143(.A1(G125), .A2(G140), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT75), .B(G125), .ZN(new_n332));
  INV_X1    g146(.A(G140), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n329), .B1(new_n334), .B2(new_n198), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n327), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G113), .B(G122), .ZN(new_n337));
  INV_X1    g151(.A(G104), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT88), .ZN(new_n340));
  INV_X1    g154(.A(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT75), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT75), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G125), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n333), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT16), .B1(new_n345), .B2(new_n330), .ZN(new_n346));
  OR2_X1    g160(.A1(KEYINPUT16), .A2(G140), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(new_n342), .B2(new_n344), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n198), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n346), .A2(G146), .A3(new_n349), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n325), .A2(KEYINPUT17), .A3(G131), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AND4_X1   g168(.A1(G143), .A2(new_n320), .A3(new_n321), .A4(G214), .ZN(new_n355));
  AOI21_X1  g169(.A(G143), .B1(new_n251), .B2(G214), .ZN(new_n356));
  OAI21_X1  g170(.A(G131), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT17), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n323), .A2(new_n210), .A3(new_n324), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT89), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n357), .A2(new_n359), .A3(KEYINPUT89), .A4(new_n358), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n336), .B(new_n340), .C1(new_n354), .C2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT90), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI211_X1 g181(.A(new_n198), .B(new_n348), .C1(new_n334), .C2(KEYINPUT16), .ZN(new_n368));
  AOI21_X1  g182(.A(G146), .B1(new_n346), .B2(new_n349), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n370), .A2(new_n353), .A3(new_n362), .A4(new_n363), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n371), .A2(KEYINPUT90), .A3(new_n336), .A4(new_n340), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT19), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n328), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n198), .B(new_n375), .C1(new_n334), .C2(new_n374), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n352), .A2(new_n376), .A3(KEYINPUT87), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n357), .A2(new_n359), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT87), .B1(new_n352), .B2(new_n376), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n336), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n339), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n373), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT20), .ZN(new_n385));
  NOR2_X1   g199(.A1(G475), .A2(G902), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT91), .ZN(new_n388));
  INV_X1    g202(.A(new_n386), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n373), .B2(new_n383), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT91), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(new_n385), .ZN(new_n392));
  AOI22_X1  g206(.A1(new_n367), .A2(new_n372), .B1(new_n382), .B2(new_n381), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT20), .B1(new_n393), .B2(new_n389), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n388), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT94), .ZN(new_n396));
  INV_X1    g210(.A(G475), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n336), .B1(new_n354), .B2(new_n364), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n339), .B1(new_n398), .B2(KEYINPUT92), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT92), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n371), .A2(new_n400), .A3(new_n336), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(G902), .B1(new_n402), .B2(new_n373), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n397), .B1(new_n403), .B2(KEYINPUT93), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT93), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n401), .A2(new_n399), .B1(new_n367), .B2(new_n372), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(G902), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n395), .A2(new_n396), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n396), .B1(new_n395), .B2(new_n408), .ZN(new_n410));
  INV_X1    g224(.A(G107), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n245), .A2(G122), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n411), .B1(new_n412), .B2(KEYINPUT14), .ZN(new_n413));
  XNOR2_X1  g227(.A(G116), .B(G122), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n413), .B(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(G128), .B(G143), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT96), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n417), .A2(new_n187), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n187), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n200), .A2(KEYINPUT13), .A3(G128), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n421), .B(KEYINPUT95), .C1(G128), .C2(new_n200), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT13), .B1(new_n200), .B2(G128), .ZN(new_n423));
  OAI221_X1 g237(.A(G134), .B1(KEYINPUT95), .B2(new_n421), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n414), .B(new_n411), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n420), .B1(new_n418), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT9), .B(G234), .ZN(new_n428));
  INV_X1    g242(.A(G217), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n428), .A2(new_n429), .A3(G953), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n427), .B(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G478), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(KEYINPUT15), .ZN(new_n433));
  OR3_X1    g247(.A1(new_n431), .A2(G902), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n431), .B2(G902), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(G234), .A2(G237), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(G952), .A3(new_n321), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT97), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n440), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n438), .A2(G902), .A3(G953), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(G898), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n437), .A2(new_n448), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n409), .A2(new_n410), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n239), .A2(G128), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n237), .B2(G128), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT24), .B(G110), .Z(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT73), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(KEYINPUT73), .A3(new_n453), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n370), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT23), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n237), .B2(G128), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n452), .B2(new_n459), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT74), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT74), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n460), .C1(new_n452), .C2(new_n459), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(G110), .A3(new_n464), .ZN(new_n465));
  OAI22_X1  g279(.A1(new_n461), .A2(G110), .B1(new_n452), .B2(new_n453), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n352), .A2(new_n329), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n458), .A2(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT22), .B(G137), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n321), .A2(G221), .A3(G234), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n470), .B(new_n471), .ZN(new_n472));
  XOR2_X1   g286(.A(new_n472), .B(KEYINPUT76), .Z(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n458), .A2(new_n465), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n466), .A2(new_n467), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n472), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n429), .B1(G234), .B2(new_n298), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(G902), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n478), .B(new_n298), .C1(new_n468), .C2(new_n473), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT25), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n475), .A2(KEYINPUT25), .A3(new_n298), .A4(new_n478), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n482), .B1(new_n487), .B2(new_n479), .ZN(new_n488));
  OAI21_X1  g302(.A(G214), .B1(G237), .B2(G902), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n238), .A2(KEYINPUT5), .A3(new_n241), .ZN(new_n490));
  INV_X1    g304(.A(G113), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT5), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n246), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT3), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n411), .A3(G104), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT79), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n495), .A2(new_n411), .A3(KEYINPUT79), .A4(G104), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G101), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT78), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n502), .B(KEYINPUT3), .C1(new_n338), .C2(G107), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n411), .A2(G104), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT3), .B1(new_n338), .B2(G107), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n504), .B1(new_n505), .B2(KEYINPUT78), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n500), .A2(new_n501), .A3(new_n503), .A4(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n338), .A2(G107), .ZN(new_n508));
  OAI21_X1  g322(.A(G101), .B1(new_n508), .B2(new_n504), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n494), .A2(new_n244), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(G110), .B(G122), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT80), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n498), .A2(new_n499), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n505), .A2(KEYINPUT78), .ZN(new_n514));
  INV_X1    g328(.A(new_n504), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n503), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n512), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT4), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n500), .A2(KEYINPUT80), .A3(new_n503), .A4(new_n506), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n517), .A2(new_n518), .A3(G101), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n248), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n500), .A2(new_n503), .A3(new_n506), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n501), .B1(new_n523), .B2(new_n512), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n522), .B1(new_n524), .B2(new_n519), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n510), .B(new_n511), .C1(new_n521), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT84), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n517), .A2(G101), .A3(new_n519), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n248), .A3(new_n520), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT84), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n510), .A4(new_n511), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT6), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n510), .B1(new_n521), .B2(new_n525), .ZN(new_n536));
  INV_X1    g350(.A(new_n511), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n534), .A2(new_n538), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n536), .A2(new_n535), .A3(new_n537), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n205), .A2(new_n332), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n332), .B1(new_n229), .B2(new_n233), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G224), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G953), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n544), .B(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n539), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT7), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT86), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(KEYINPUT86), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n544), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(KEYINPUT86), .B(new_n550), .C1(new_n542), .C2(new_n543), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT85), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n510), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n510), .A2(new_n556), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n494), .A2(new_n244), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n507), .A2(new_n509), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n557), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n511), .B(KEYINPUT8), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n555), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(G902), .B1(new_n564), .B2(new_n534), .ZN(new_n565));
  OAI21_X1  g379(.A(G210), .B1(G237), .B2(G902), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n548), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n566), .B1(new_n548), .B2(new_n565), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n489), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G469), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT82), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n205), .A2(KEYINPUT10), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n571), .B1(new_n560), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n205), .A2(KEYINPUT10), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n574), .A2(new_n507), .A3(KEYINPUT82), .A4(new_n509), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT10), .ZN(new_n576));
  AOI21_X1  g390(.A(G128), .B1(new_n199), .B2(new_n201), .ZN(new_n577));
  INV_X1    g391(.A(new_n203), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT81), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT81), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n580), .B(new_n203), .C1(new_n204), .C2(G128), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n202), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(new_n507), .A3(new_n509), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n573), .A2(new_n575), .B1(new_n576), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n530), .A2(new_n234), .A3(new_n520), .ZN(new_n585));
  INV_X1    g399(.A(new_n224), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(G110), .B(G140), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n321), .A2(G227), .ZN(new_n589));
  XOR2_X1   g403(.A(new_n588), .B(new_n589), .Z(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n205), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n560), .A2(new_n592), .ZN(new_n593));
  AOI22_X1  g407(.A1(new_n593), .A2(new_n583), .B1(new_n223), .B2(new_n218), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n271), .A2(KEYINPUT12), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n593), .B2(new_n583), .ZN(new_n596));
  OAI22_X1  g410(.A1(new_n594), .A2(KEYINPUT12), .B1(new_n596), .B2(KEYINPUT83), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n596), .A2(KEYINPUT83), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n587), .B(new_n591), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n573), .A2(new_n575), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n583), .A2(new_n576), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n520), .A2(new_n234), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(new_n525), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n224), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n591), .B1(new_n606), .B2(new_n587), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n570), .B(new_n298), .C1(new_n600), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(G469), .A2(G902), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n587), .B1(new_n597), .B2(new_n598), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n590), .B(KEYINPUT77), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n606), .A2(new_n587), .A3(new_n591), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(G469), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(G221), .B1(new_n428), .B2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n569), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n319), .A2(new_n450), .A3(new_n488), .A4(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT98), .B(G101), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G3));
  NOR2_X1   g435(.A1(new_n431), .A2(G902), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT99), .B(G478), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n431), .B(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n432), .A2(G902), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n391), .B1(new_n390), .B2(new_n385), .ZN(new_n629));
  NOR4_X1   g443(.A1(new_n393), .A2(KEYINPUT91), .A3(KEYINPUT20), .A4(new_n389), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n390), .A2(new_n385), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n403), .A2(KEYINPUT93), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n633), .A2(new_n407), .A3(G475), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT94), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n395), .A2(new_n396), .A3(new_n408), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n628), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n569), .B1(new_n444), .B2(new_n447), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(G472), .B1(new_n313), .B2(G902), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n315), .A2(new_n640), .A3(new_n316), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n488), .A2(new_n616), .A3(new_n615), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n639), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT34), .B(G104), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  XOR2_X1   g460(.A(new_n448), .B(KEYINPUT100), .Z(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n387), .A2(new_n394), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n408), .A2(new_n649), .A3(new_n436), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n569), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n643), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n651), .A2(new_n641), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NAND2_X1  g469(.A1(new_n487), .A2(new_n479), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n474), .A2(KEYINPUT36), .ZN(new_n657));
  XOR2_X1   g471(.A(new_n468), .B(new_n657), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n480), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n450), .A2(new_n618), .A3(new_n641), .A4(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  INV_X1    g477(.A(new_n660), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n307), .B2(new_n318), .ZN(new_n665));
  OR2_X1    g479(.A1(KEYINPUT101), .A2(G900), .ZN(new_n666));
  NAND2_X1  g480(.A1(KEYINPUT101), .A2(G900), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n445), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n444), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n387), .B2(new_n394), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n408), .A2(new_n436), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n665), .A2(new_n618), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  INV_X1    g488(.A(new_n617), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n669), .B(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT40), .Z(new_n679));
  AOI21_X1  g493(.A(new_n255), .B1(new_n250), .B2(new_n299), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n680), .A2(KEYINPUT103), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(KEYINPUT103), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n276), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(G902), .B1(new_n683), .B2(KEYINPUT104), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(KEYINPUT104), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n312), .A2(new_n311), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n314), .B1(new_n686), .B2(new_n283), .ZN(new_n687));
  AOI22_X1  g501(.A1(new_n685), .A2(G472), .B1(new_n687), .B2(KEYINPUT32), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n660), .B1(new_n688), .B2(new_n318), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n409), .A2(new_n410), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n436), .A2(new_n489), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n566), .ZN(new_n693));
  INV_X1    g507(.A(new_n547), .ZN(new_n694));
  AOI211_X1 g508(.A(new_n694), .B(new_n540), .C1(new_n534), .C2(new_n538), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n564), .A2(new_n534), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n298), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n693), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n548), .A2(new_n565), .A3(new_n566), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n679), .A2(new_n689), .A3(new_n692), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  AOI211_X1 g518(.A(new_n670), .B(new_n628), .C1(new_n635), .C2(new_n636), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n665), .A2(new_n705), .A3(new_n618), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G146), .ZN(G48));
  AND3_X1   g521(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n586), .B1(new_n584), .B2(new_n585), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n590), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n599), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n298), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G469), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n713), .A2(new_n616), .A3(new_n608), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n315), .A2(new_n317), .A3(new_n316), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n294), .A2(new_n305), .A3(new_n306), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n488), .B(new_n714), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n639), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT41), .B(G113), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  INV_X1    g534(.A(new_n488), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n307), .B2(new_n318), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n651), .A3(new_n714), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G116), .ZN(G18));
  NAND3_X1  g538(.A1(new_n713), .A2(new_n616), .A3(new_n608), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT106), .B1(new_n569), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT106), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n714), .A2(new_n727), .A3(new_n489), .A4(new_n700), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n665), .A2(new_n729), .A3(new_n450), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  AOI22_X1  g545(.A1(new_n276), .A2(KEYINPUT31), .B1(new_n277), .B2(new_n300), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n686), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n293), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n640), .A2(new_n734), .A3(new_n488), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n640), .A2(new_n734), .A3(new_n737), .A4(new_n488), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n567), .A2(new_n568), .ZN(new_n740));
  AOI211_X1 g554(.A(new_n691), .B(new_n740), .C1(new_n635), .C2(new_n636), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n725), .A2(new_n648), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n739), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  AND3_X1   g558(.A1(new_n640), .A2(new_n660), .A3(new_n734), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n705), .A2(new_n729), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n698), .A2(new_n748), .A3(new_n489), .A4(new_n699), .ZN(new_n749));
  INV_X1    g563(.A(new_n489), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT109), .B1(new_n700), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n637), .A2(new_n669), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n614), .A2(new_n609), .ZN(new_n753));
  AOI211_X1 g567(.A(G469), .B(G902), .C1(new_n710), .C2(new_n599), .ZN(new_n754));
  OAI211_X1 g568(.A(KEYINPUT108), .B(new_n616), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT108), .B1(new_n615), .B2(new_n616), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n759), .B1(new_n687), .B2(KEYINPUT32), .ZN(new_n760));
  OAI211_X1 g574(.A(KEYINPUT110), .B(new_n317), .C1(new_n313), .C2(new_n314), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n758), .B(new_n488), .C1(new_n762), .C2(new_n716), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT42), .B1(new_n752), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n757), .ZN(new_n765));
  AND4_X1   g579(.A1(new_n749), .A2(new_n751), .A3(new_n765), .A4(new_n755), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n767), .A3(new_n722), .A4(new_n705), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(new_n210), .ZN(G33));
  AND2_X1   g584(.A1(new_n751), .A2(new_n749), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n722), .A2(new_n771), .A3(new_n672), .A4(new_n758), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  NAND2_X1  g587(.A1(new_n642), .A2(new_n660), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT43), .B1(new_n690), .B2(KEYINPUT112), .ZN(new_n775));
  INV_X1    g589(.A(new_n628), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n690), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n690), .B(new_n776), .C1(KEYINPUT112), .C2(KEYINPUT43), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n774), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT44), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(KEYINPUT44), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n612), .A2(new_n613), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n612), .A2(KEYINPUT45), .A3(new_n613), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(G469), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n609), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(KEYINPUT111), .A3(new_n608), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n787), .A2(new_n609), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n789), .B1(KEYINPUT46), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT111), .B1(new_n788), .B2(new_n608), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n616), .A3(new_n677), .ZN(new_n794));
  INV_X1    g608(.A(new_n771), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n781), .A2(new_n782), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  NAND2_X1  g612(.A1(new_n793), .A2(new_n616), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(KEYINPUT113), .B2(KEYINPUT47), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n752), .A2(new_n319), .A3(new_n488), .ZN(new_n801));
  XNOR2_X1  g615(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n793), .A2(new_n616), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT114), .B(G140), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(G42));
  NOR2_X1   g620(.A1(new_n777), .A2(new_n702), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n688), .A2(new_n318), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n713), .A2(new_n608), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT49), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n488), .A2(new_n489), .A3(new_n616), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(KEYINPUT49), .B2(new_n810), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n807), .A2(new_n809), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n743), .A2(new_n730), .A3(new_n723), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n409), .A2(new_n410), .A3(new_n437), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n569), .A2(new_n648), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n641), .A3(new_n652), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n661), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n718), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n637), .A2(new_n641), .A3(new_n652), .A4(new_n818), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n619), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n488), .B1(new_n715), .B2(new_n716), .ZN(new_n825));
  INV_X1    g639(.A(new_n449), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n690), .A2(new_n826), .A3(new_n618), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n823), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT115), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n816), .A2(new_n821), .A3(new_n824), .A4(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n436), .B1(new_n407), .B2(new_n404), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n616), .A3(new_n615), .A4(new_n671), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n664), .B(new_n832), .C1(new_n307), .C2(new_n318), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n637), .A2(new_n669), .A3(new_n745), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n771), .A2(new_n833), .B1(new_n834), .B2(new_n766), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n764), .A3(new_n768), .A4(new_n772), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT116), .B1(new_n830), .B2(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n619), .A2(new_n822), .A3(new_n823), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n822), .B1(new_n619), .B2(new_n823), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n661), .B(new_n819), .C1(new_n717), .C2(new_n639), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n838), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n766), .A2(new_n705), .A3(new_n745), .ZN(new_n842));
  INV_X1    g656(.A(new_n832), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n665), .A2(new_n771), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n772), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n769), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n841), .A2(new_n846), .A3(new_n847), .A4(new_n816), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n837), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n741), .A2(new_n689), .A3(new_n675), .A4(new_n669), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(new_n706), .A3(new_n673), .A4(new_n746), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT52), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n849), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  XOR2_X1   g669(.A(KEYINPUT118), .B(KEYINPUT52), .Z(new_n856));
  NAND2_X1  g670(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n673), .A2(new_n746), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n673), .A2(new_n746), .A3(KEYINPUT117), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n850), .A2(new_n706), .A3(KEYINPUT52), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n857), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n849), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n855), .A2(KEYINPUT120), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n852), .B1(new_n837), .B2(new_n848), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n854), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n815), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n830), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n864), .A2(KEYINPUT53), .A3(new_n872), .A4(new_n846), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n815), .B(new_n873), .C1(new_n868), .C2(new_n854), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n444), .B1(new_n778), .B2(new_n779), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n702), .A2(new_n489), .A3(new_n725), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n739), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT50), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n810), .A2(new_n616), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n800), .B2(new_n803), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n876), .A2(new_n739), .A3(new_n771), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n795), .A2(new_n725), .ZN(new_n885));
  AND4_X1   g699(.A1(new_n488), .A2(new_n885), .A3(new_n443), .A4(new_n809), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n690), .A3(new_n628), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n876), .A2(new_n745), .A3(new_n885), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n880), .A2(new_n884), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT51), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n880), .A2(new_n884), .A3(KEYINPUT51), .A4(new_n889), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n321), .A2(G952), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n886), .B2(new_n637), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT121), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n876), .A2(new_n729), .A3(new_n739), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n488), .B1(new_n762), .B2(new_n716), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n876), .A2(new_n900), .A3(new_n885), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT48), .Z(new_n902));
  AOI21_X1  g716(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n898), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n892), .A2(new_n893), .A3(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n871), .A2(new_n875), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(G952), .A2(G953), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n814), .B1(new_n906), .B2(new_n907), .ZN(G75));
  OAI21_X1  g722(.A(new_n873), .B1(new_n868), .B2(new_n854), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(G210), .A3(G902), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT56), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n539), .A2(new_n541), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(new_n547), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT55), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n910), .B2(new_n911), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n321), .A2(G952), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(G51));
  NAND2_X1  g732(.A1(new_n909), .A2(KEYINPUT54), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n874), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n609), .B(KEYINPUT57), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n711), .B(KEYINPUT122), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n787), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n909), .A2(G902), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n917), .B1(new_n924), .B2(new_n926), .ZN(G54));
  NAND4_X1  g741(.A1(new_n909), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n928), .A2(new_n393), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n393), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n917), .ZN(G60));
  INV_X1    g745(.A(new_n626), .ZN(new_n932));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT59), .Z(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n920), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n917), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n934), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n871), .B2(new_n875), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n932), .B2(new_n940), .ZN(G63));
  XNOR2_X1  g755(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n429), .A2(new_n298), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n909), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n475), .A2(new_n478), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n909), .A2(new_n658), .A3(new_n944), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n937), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n947), .A2(KEYINPUT61), .A3(new_n937), .A4(new_n948), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(G66));
  OAI21_X1  g767(.A(G953), .B1(new_n446), .B2(new_n545), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n872), .B2(G953), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n912), .B1(G898), .B2(new_n321), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(G69));
  AOI21_X1  g771(.A(new_n321), .B1(G227), .B2(G900), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n860), .A2(new_n706), .A3(new_n861), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n703), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT62), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT62), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n962), .A3(new_n703), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n825), .A2(new_n678), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n964), .B(new_n771), .C1(new_n637), .C2(new_n817), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n804), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n961), .A2(new_n797), .A3(new_n963), .A4(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n321), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n270), .A2(new_n265), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT124), .Z(new_n970));
  OAI21_X1  g784(.A(new_n375), .B1(new_n334), .B2(new_n374), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n972), .ZN(new_n974));
  INV_X1    g788(.A(G900), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n321), .ZN(new_n976));
  INV_X1    g790(.A(new_n769), .ZN(new_n977));
  INV_X1    g791(.A(new_n794), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n741), .A3(new_n900), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n804), .A2(new_n977), .A3(new_n979), .A4(new_n772), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n797), .A2(new_n959), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n797), .A2(new_n983), .A3(new_n959), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n980), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n976), .B1(new_n985), .B2(new_n321), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n973), .B1(new_n986), .B2(KEYINPUT127), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n988));
  AOI211_X1 g802(.A(new_n988), .B(new_n976), .C1(new_n985), .C2(new_n321), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n958), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n986), .A2(new_n958), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n973), .A2(KEYINPUT125), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n968), .A2(new_n993), .A3(new_n972), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n991), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n990), .A2(new_n995), .ZN(G72));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n967), .B2(new_n830), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n268), .A2(new_n275), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n277), .B1(new_n1001), .B2(new_n250), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n998), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n985), .B2(new_n872), .ZN(new_n1005));
  OAI211_X1 g819(.A(new_n1003), .B(new_n937), .C1(new_n295), .C2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n867), .A2(new_n870), .ZN(new_n1007));
  INV_X1    g821(.A(new_n295), .ZN(new_n1008));
  NOR3_X1   g822(.A1(new_n1002), .A2(new_n1008), .A3(new_n1004), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1006), .B1(new_n1007), .B2(new_n1009), .ZN(G57));
endmodule


