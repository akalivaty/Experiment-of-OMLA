//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n580, new_n581, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n634, new_n635, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204, new_n1206, new_n1207, new_n1208, new_n1209;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT3), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  INV_X1    g044(.A(G101), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT67), .B(G2104), .ZN(new_n471));
  OAI22_X1  g046(.A1(new_n468), .A2(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G125), .ZN(new_n476));
  INV_X1    g051(.A(G113), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(new_n465), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n468), .A2(new_n473), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n466), .B1(new_n471), .B2(KEYINPUT3), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(new_n473), .ZN(new_n486));
  NOR2_X1   g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(new_n473), .B2(G112), .ZN(new_n488));
  OAI221_X1 g063(.A(new_n483), .B1(new_n484), .B2(new_n486), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT69), .B1(new_n473), .B2(G114), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(new_n495), .A3(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT70), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n492), .A2(new_n493), .A3(new_n496), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n475), .A2(G138), .A3(new_n473), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT4), .A2(G138), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n464), .A2(new_n473), .A3(new_n467), .A4(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n501), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n485), .A2(KEYINPUT68), .A3(G126), .A4(G2105), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n464), .A2(G126), .A3(G2105), .A4(new_n467), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n507), .A2(new_n512), .ZN(G164));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n517), .A2(KEYINPUT5), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT5), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G543), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n514), .A2(new_n515), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n519), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT71), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n519), .B(new_n529), .C1(new_n520), .C2(new_n526), .ZN(new_n530));
  NAND2_X1  g105(.A1(G75), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n521), .A2(new_n523), .ZN(new_n532));
  INV_X1    g107(.A(G62), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n528), .A2(new_n530), .B1(G651), .B2(new_n534), .ZN(G166));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  INV_X1    g111(.A(G89), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n516), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n538), .A2(new_n524), .B1(new_n518), .B2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  INV_X1    g119(.A(G77), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n532), .A2(new_n544), .B1(new_n545), .B2(new_n517), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT72), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n548));
  OAI221_X1 g123(.A(new_n548), .B1(new_n545), .B2(new_n517), .C1(new_n532), .C2(new_n544), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n547), .A2(G651), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n547), .A2(KEYINPUT73), .A3(new_n549), .A4(G651), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n526), .ZN(new_n555));
  XNOR2_X1  g130(.A(KEYINPUT74), .B(G90), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n518), .A2(G52), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT75), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n552), .A2(new_n553), .B1(G52), .B2(new_n518), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(new_n562), .A3(new_n557), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G171));
  NAND2_X1  g139(.A1(G68), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G56), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n532), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT76), .ZN(new_n569));
  INV_X1    g144(.A(G81), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n525), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G43), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n526), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G860), .ZN(G153));
  AND3_X1   g152(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G36), .ZN(G176));
  NAND2_X1  g154(.A1(G1), .A2(G3), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT8), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(new_n581), .ZN(G188));
  INV_X1    g157(.A(G91), .ZN(new_n583));
  OR4_X1    g158(.A1(KEYINPUT77), .A2(new_n532), .A3(new_n516), .A4(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT77), .B1(new_n526), .B2(new_n583), .ZN(new_n585));
  NAND2_X1  g160(.A1(G78), .A2(G543), .ZN(new_n586));
  XOR2_X1   g161(.A(KEYINPUT78), .B(G65), .Z(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n587), .B2(new_n532), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n584), .A2(new_n585), .B1(G651), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n518), .A2(G53), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT9), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(G299));
  INV_X1    g167(.A(G171), .ZN(G301));
  INV_X1    g168(.A(G166), .ZN(G303));
  NAND2_X1  g169(.A1(new_n555), .A2(G87), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n518), .A2(G49), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(G288));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  INV_X1    g174(.A(G48), .ZN(new_n600));
  OAI22_X1  g175(.A1(new_n526), .A2(new_n599), .B1(new_n571), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n524), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G651), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G305));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  INV_X1    g182(.A(G47), .ZN(new_n608));
  OAI22_X1  g183(.A1(new_n526), .A2(new_n607), .B1(new_n571), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(G72), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G60), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n532), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G651), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n609), .A2(new_n614), .ZN(G290));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n555), .A2(new_n616), .A3(G92), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n518), .A2(G54), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  INV_X1    g194(.A(G66), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n532), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G651), .ZN(new_n622));
  INV_X1    g197(.A(G92), .ZN(new_n623));
  OAI21_X1  g198(.A(KEYINPUT10), .B1(new_n526), .B2(new_n623), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n617), .A2(new_n618), .A3(new_n622), .A4(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G171), .B2(new_n626), .ZN(G284));
  OAI21_X1  g203(.A(new_n627), .B1(G171), .B2(new_n626), .ZN(G321));
  NAND2_X1  g204(.A1(G286), .A2(G868), .ZN(new_n630));
  INV_X1    g205(.A(G299), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G297));
  OAI21_X1  g207(.A(new_n630), .B1(new_n631), .B2(G868), .ZN(G280));
  INV_X1    g208(.A(new_n625), .ZN(new_n634));
  INV_X1    g209(.A(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(G860), .ZN(G148));
  NAND2_X1  g211(.A1(new_n575), .A2(new_n626), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n625), .A2(G559), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n626), .B2(new_n638), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n482), .A2(G123), .ZN(new_n641));
  INV_X1    g216(.A(G135), .ZN(new_n642));
  NOR2_X1   g217(.A1(G99), .A2(G2105), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(new_n473), .B2(G111), .ZN(new_n644));
  OAI221_X1 g219(.A(new_n641), .B1(new_n642), .B2(new_n486), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT80), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n475), .A2(new_n473), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n648), .A2(new_n471), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT13), .B(G2100), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n647), .A2(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2435), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2438), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT14), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2443), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2446), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(G14), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(G401));
  XOR2_X1   g245(.A(G2072), .B(G2078), .Z(new_n671));
  XOR2_X1   g246(.A(G2067), .B(G2678), .Z(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n671), .B1(new_n675), .B2(KEYINPUT18), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G2096), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n673), .A2(new_n674), .ZN(new_n680));
  AOI21_X1  g255(.A(KEYINPUT18), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n678), .B(new_n681), .Z(G227));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT83), .Z(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n683), .A2(new_n684), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT84), .ZN(new_n694));
  INV_X1    g269(.A(new_n692), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n695), .A2(new_n688), .A3(new_n685), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n691), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT21), .B(G1986), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1991), .B(G1996), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT22), .B(G1981), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n701), .B(new_n702), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  INV_X1    g279(.A(G1976), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n595), .A2(G16), .A3(new_n596), .A4(new_n597), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT33), .ZN(new_n707));
  OR2_X1    g282(.A1(G16), .A2(G23), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n707), .B1(new_n706), .B2(new_n708), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n705), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n711), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n713), .A2(G1976), .A3(new_n709), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G22), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G166), .B2(new_n716), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT87), .B(G1971), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n718), .A2(new_n720), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n715), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g298(.A(G16), .B1(new_n601), .B2(new_n604), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n716), .A2(G6), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT32), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n724), .A2(KEYINPUT32), .A3(new_n725), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT86), .B(G1981), .Z(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n728), .A2(new_n731), .A3(new_n729), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(KEYINPUT34), .B1(new_n723), .B2(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n733), .A2(new_n734), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n718), .B(new_n719), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT34), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n737), .A2(new_n738), .A3(new_n739), .A4(new_n715), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n736), .A2(new_n740), .A3(KEYINPUT88), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT36), .ZN(new_n742));
  INV_X1    g317(.A(new_n486), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G131), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n482), .A2(G119), .ZN(new_n745));
  OR2_X1    g320(.A1(G95), .A2(G2105), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n746), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  MUX2_X1   g323(.A(G25), .B(new_n748), .S(G29), .Z(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(KEYINPUT85), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT35), .B(G1991), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(KEYINPUT85), .ZN(new_n752));
  AND3_X1   g327(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n751), .B1(new_n750), .B2(new_n752), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G16), .A2(G24), .ZN(new_n756));
  INV_X1    g331(.A(G290), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1986), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n741), .A2(new_n742), .A3(new_n755), .A4(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n755), .A2(new_n736), .A3(KEYINPUT88), .A4(new_n740), .ZN(new_n762));
  OAI21_X1  g337(.A(KEYINPUT36), .B1(new_n762), .B2(new_n759), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT89), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G4), .B2(G16), .ZN(new_n766));
  OR3_X1    g341(.A1(new_n765), .A2(G4), .A3(G16), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n766), .B(new_n767), .C1(new_n625), .C2(new_n716), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1348), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OR2_X1    g346(.A1(G29), .A2(G33), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT94), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT25), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n743), .A2(G139), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n777));
  OAI211_X1 g352(.A(new_n775), .B(new_n776), .C1(new_n473), .C2(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G29), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n772), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G2072), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n716), .A2(G5), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G171), .B2(new_n716), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(G1961), .ZN(new_n785));
  AND2_X1   g360(.A1(KEYINPUT24), .A2(G34), .ZN(new_n786));
  NOR2_X1   g361(.A1(KEYINPUT24), .A2(G34), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n779), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n480), .B2(new_n779), .ZN(new_n789));
  INV_X1    g364(.A(G2084), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G29), .A2(G32), .ZN(new_n792));
  INV_X1    g367(.A(G141), .ZN(new_n793));
  INV_X1    g368(.A(G105), .ZN(new_n794));
  OAI22_X1  g369(.A1(new_n468), .A2(new_n793), .B1(new_n794), .B2(new_n471), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n795), .A2(new_n473), .B1(new_n482), .B2(G129), .ZN(new_n796));
  NAND3_X1  g371(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n797));
  XOR2_X1   g372(.A(new_n797), .B(KEYINPUT26), .Z(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n792), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT27), .B(G1996), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n785), .A2(new_n791), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT95), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n785), .A2(KEYINPUT95), .A3(new_n791), .A4(new_n803), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n806), .A2(new_n807), .B1(G1961), .B2(new_n784), .ZN(new_n808));
  NAND4_X1  g383(.A1(new_n764), .A2(new_n771), .A3(new_n782), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n716), .A2(KEYINPUT23), .A3(G20), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT23), .ZN(new_n811));
  INV_X1    g386(.A(G20), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(G16), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n810), .B(new_n813), .C1(new_n631), .C2(new_n716), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G1956), .ZN(new_n815));
  NOR2_X1   g390(.A1(G27), .A2(G29), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G164), .B2(G29), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n815), .B1(G2078), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n780), .A2(new_n781), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT31), .B(G11), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n716), .A2(G19), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n576), .B2(new_n716), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT92), .B(G1341), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n482), .A2(G128), .ZN(new_n826));
  INV_X1    g401(.A(G140), .ZN(new_n827));
  NOR2_X1   g402(.A1(G104), .A2(G2105), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(new_n473), .B2(G116), .ZN(new_n829));
  OAI221_X1 g404(.A(new_n826), .B1(new_n827), .B2(new_n486), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(G29), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT93), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n779), .A2(G26), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT28), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G2067), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n779), .A2(G35), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(G162), .B2(new_n779), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT29), .Z(new_n839));
  INV_X1    g414(.A(G2090), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n817), .A2(G2078), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n840), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT30), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n844), .A2(G28), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(G28), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n846), .A3(new_n779), .ZN(new_n847));
  NAND2_X1  g422(.A1(G168), .A2(G16), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(G16), .B2(G21), .ZN(new_n849));
  INV_X1    g424(.A(G1966), .ZN(new_n850));
  OAI221_X1 g425(.A(new_n847), .B1(new_n790), .B2(new_n789), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n801), .A2(new_n802), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n853), .ZN(new_n854));
  NOR4_X1   g429(.A1(new_n809), .A2(new_n825), .A3(new_n836), .A4(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n645), .A2(new_n779), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n849), .A2(new_n850), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(G150));
  INV_X1    g433(.A(KEYINPUT96), .ZN(new_n859));
  NAND2_X1  g434(.A1(G150), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n855), .A2(KEYINPUT96), .A3(new_n856), .A4(new_n857), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(G311));
  INV_X1    g437(.A(G93), .ZN(new_n863));
  INV_X1    g438(.A(G55), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n526), .A2(new_n863), .B1(new_n571), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n866), .A2(new_n603), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(G860), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT37), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n576), .A2(new_n869), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n575), .A2(new_n868), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n625), .A2(new_n635), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n871), .B1(new_n878), .B2(G860), .ZN(G145));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n498), .A2(new_n500), .B1(new_n503), .B2(new_n502), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n881), .A2(new_n506), .A3(new_n511), .A4(new_n508), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n508), .A2(new_n511), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n885), .A2(KEYINPUT97), .A3(new_n881), .A4(new_n506), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(new_n778), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n482), .A2(G130), .ZN(new_n889));
  INV_X1    g464(.A(G142), .ZN(new_n890));
  NOR2_X1   g465(.A1(G106), .A2(G2105), .ZN(new_n891));
  OAI21_X1  g466(.A(G2104), .B1(new_n473), .B2(G118), .ZN(new_n892));
  OAI221_X1 g467(.A(new_n889), .B1(new_n890), .B2(new_n486), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n651), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n888), .B(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n830), .B(new_n748), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n800), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n897), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n645), .B(G160), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(G162), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n880), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  AOI211_X1 g479(.A(KEYINPUT98), .B(new_n904), .C1(new_n898), .C2(new_n899), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n900), .ZN(new_n907));
  AOI21_X1  g482(.A(G37), .B1(new_n907), .B2(new_n904), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g485(.A1(new_n869), .A2(new_n626), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n912));
  NAND2_X1  g487(.A1(G299), .A2(new_n634), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n625), .A2(new_n589), .A3(new_n591), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n912), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT99), .ZN(new_n919));
  INV_X1    g494(.A(new_n914), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n625), .B1(new_n589), .B2(new_n591), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n914), .A2(KEYINPUT99), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n918), .B1(new_n924), .B2(new_n916), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n917), .B1(new_n925), .B2(new_n912), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n874), .B(new_n638), .ZN(new_n927));
  MUX2_X1   g502(.A(new_n926), .B(new_n915), .S(new_n927), .Z(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(KEYINPUT42), .ZN(new_n929));
  XNOR2_X1  g504(.A(G166), .B(new_n605), .ZN(new_n930));
  XNOR2_X1  g505(.A(G290), .B(G288), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n930), .B1(KEYINPUT101), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(KEYINPUT101), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n932), .B(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n929), .B(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n911), .B1(new_n935), .B2(new_n626), .ZN(G295));
  OAI21_X1  g511(.A(new_n911), .B1(new_n935), .B2(new_n626), .ZN(G331));
  NOR2_X1   g512(.A1(new_n559), .A2(KEYINPUT75), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n562), .B1(new_n561), .B2(new_n557), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n938), .A2(new_n939), .A3(G286), .ZN(new_n940));
  AOI21_X1  g515(.A(G168), .B1(new_n560), .B2(new_n563), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n874), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(G286), .B1(new_n938), .B2(new_n939), .ZN(new_n943));
  INV_X1    g518(.A(new_n874), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n560), .A2(G168), .A3(new_n563), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(KEYINPUT102), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n943), .A2(new_n944), .A3(new_n948), .A4(new_n945), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n947), .A2(new_n926), .A3(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n920), .A2(new_n921), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT103), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n942), .A2(new_n952), .A3(new_n946), .ZN(new_n953));
  OAI211_X1 g528(.A(KEYINPUT103), .B(new_n874), .C1(new_n940), .C2(new_n941), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n956), .B2(new_n934), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n959));
  OR3_X1    g534(.A1(new_n951), .A2(KEYINPUT104), .A3(KEYINPUT41), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT104), .B1(new_n951), .B2(KEYINPUT41), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n960), .B(new_n961), .C1(new_n916), .C2(new_n924), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n953), .A2(new_n962), .A3(new_n954), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n947), .A2(new_n949), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n951), .ZN(new_n965));
  INV_X1    g540(.A(new_n934), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n959), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n953), .A2(new_n954), .A3(new_n962), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n951), .B1(new_n947), .B2(new_n949), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n959), .B(new_n966), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n957), .B(new_n958), .C1(new_n967), .C2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n966), .B1(new_n950), .B2(new_n955), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n947), .A2(new_n926), .A3(new_n949), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n953), .A2(new_n954), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n934), .B(new_n974), .C1(new_n975), .C2(new_n951), .ZN(new_n976));
  INV_X1    g551(.A(G37), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n973), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n958), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n957), .B1(new_n967), .B2(new_n971), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(new_n982), .B2(new_n958), .ZN(new_n983));
  MUX2_X1   g558(.A(new_n980), .B(new_n983), .S(KEYINPUT44), .Z(G397));
  INV_X1    g559(.A(KEYINPUT62), .ZN(new_n985));
  XOR2_X1   g560(.A(KEYINPUT110), .B(G8), .Z(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(G168), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(new_n507), .B2(new_n512), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI211_X1 g567(.A(KEYINPUT108), .B(new_n989), .C1(new_n507), .C2(new_n512), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT50), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT106), .B(G40), .Z(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n474), .A2(new_n479), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n990), .B2(KEYINPUT50), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n994), .A2(new_n999), .A3(G2084), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n992), .A2(new_n1001), .A3(new_n993), .ZN(new_n1002));
  INV_X1    g577(.A(new_n997), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT45), .B(new_n989), .C1(new_n507), .C2(new_n512), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(G1966), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n988), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT120), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT51), .ZN(new_n1010));
  INV_X1    g585(.A(G8), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n850), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT50), .ZN(new_n1014));
  INV_X1    g589(.A(new_n993), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT108), .B1(new_n882), .B2(new_n989), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1017), .A2(new_n790), .A3(new_n998), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1011), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n988), .B1(new_n1019), .B2(KEYINPUT121), .ZN(new_n1020));
  OAI21_X1  g595(.A(G8), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT121), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1010), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n987), .B1(new_n1013), .B2(new_n1018), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n1025), .A2(KEYINPUT51), .A3(new_n988), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n985), .B(new_n1009), .C1(new_n1024), .C2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1028), .A2(KEYINPUT109), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(KEYINPUT109), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1029), .B(new_n1030), .C1(G166), .C2(new_n1011), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G303), .A2(G8), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1031), .B1(new_n1032), .B2(new_n1030), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT107), .B(G1971), .Z(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AOI211_X1 g610(.A(new_n1001), .B(G1384), .C1(new_n884), .C2(new_n886), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n997), .B1(new_n990), .B2(new_n1001), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1035), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1017), .A2(new_n840), .A3(new_n998), .ZN(new_n1040));
  AOI211_X1 g615(.A(new_n1011), .B(new_n1033), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n1042));
  INV_X1    g617(.A(G1981), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1042), .B1(new_n605), .B2(new_n1043), .ZN(new_n1044));
  NOR4_X1   g619(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT111), .A4(G1981), .ZN(new_n1045));
  OAI22_X1  g620(.A1(new_n1044), .A2(new_n1045), .B1(new_n1043), .B2(new_n605), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT49), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT112), .ZN(new_n1050));
  OAI221_X1 g625(.A(new_n1050), .B1(new_n1043), .B2(new_n605), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1003), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1048), .A2(new_n1051), .A3(new_n986), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(G288), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G1976), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(G288), .B2(new_n705), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1052), .A2(new_n986), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1052), .A2(new_n986), .A3(new_n1055), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1053), .B(new_n1057), .C1(new_n1058), .C2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1041), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1062), .B1(new_n994), .B2(new_n999), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1017), .A2(KEYINPUT115), .A3(new_n998), .ZN(new_n1064));
  INV_X1    g639(.A(G1961), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n887), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n1067));
  INV_X1    g642(.A(G2078), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n1037), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1002), .A2(new_n1005), .A3(new_n1068), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1070), .B1(new_n1073), .B2(KEYINPUT122), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1074), .B1(KEYINPUT122), .B2(new_n1073), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n990), .B2(KEYINPUT50), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n882), .A2(KEYINPUT114), .A3(new_n1014), .A4(new_n989), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n992), .A2(KEYINPUT50), .A3(new_n993), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n1003), .A3(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1039), .B1(G2090), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(new_n986), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1033), .ZN(new_n1085));
  AND4_X1   g660(.A1(G171), .A2(new_n1061), .A3(new_n1076), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1027), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT124), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1009), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT62), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1027), .A2(new_n1091), .A3(new_n1086), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT125), .ZN(new_n1094));
  INV_X1    g669(.A(G1956), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1082), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT56), .B(G2072), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1067), .A2(new_n1037), .A3(new_n1097), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(G299), .B(KEYINPUT57), .Z(new_n1100));
  NOR2_X1   g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(G1348), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1063), .A2(new_n1064), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n997), .B1(new_n992), .B2(new_n993), .ZN(new_n1104));
  INV_X1    g679(.A(G2067), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1096), .A2(new_n1100), .A3(new_n1098), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1101), .B1(new_n1109), .B2(new_n634), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n625), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1103), .A2(new_n634), .A3(new_n1106), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(KEYINPUT60), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1099), .A2(KEYINPUT119), .A3(new_n1100), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT119), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1108), .A2(new_n1115), .A3(KEYINPUT61), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1108), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1103), .A2(new_n1122), .A3(new_n634), .A4(new_n1106), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT58), .B(G1341), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1124), .B1(new_n1104), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1996), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1067), .A2(new_n1127), .A3(new_n1037), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1125), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1052), .A2(KEYINPUT116), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1126), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n575), .A2(KEYINPUT117), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1133), .A2(KEYINPUT59), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(KEYINPUT59), .ZN(new_n1135));
  OAI211_X1 g710(.A(new_n1121), .B(new_n1123), .C1(new_n1134), .C2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1110), .B1(new_n1117), .B2(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(G171), .B(KEYINPUT54), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1076), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1061), .A2(new_n1085), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n478), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(G2105), .B1(new_n478), .B2(new_n1142), .ZN(new_n1144));
  OAI21_X1  g719(.A(G40), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1145), .B1(new_n473), .B2(new_n472), .ZN(new_n1146));
  AOI21_X1  g721(.A(G1384), .B1(new_n884), .B2(new_n886), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1147), .A2(KEYINPUT45), .ZN(new_n1148));
  NOR4_X1   g723(.A1(new_n1148), .A2(new_n1036), .A3(new_n1070), .A4(G2078), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1139), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1141), .B1(new_n1072), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1137), .A2(new_n1140), .A3(new_n1151), .A4(new_n1089), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(G8), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1060), .A2(new_n1154), .A3(new_n1033), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1053), .A2(new_n705), .A3(new_n1054), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT113), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1157), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1052), .A2(new_n986), .ZN(new_n1161));
  NOR3_X1   g736(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT63), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1025), .A2(G168), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1163), .B1(new_n1141), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1163), .B1(new_n1154), .B2(new_n1033), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1061), .A2(new_n1166), .A3(G168), .A4(new_n1025), .ZN(new_n1167));
  AOI211_X1 g742(.A(new_n1155), .B(new_n1162), .C1(new_n1165), .C2(new_n1167), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1152), .A2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1088), .A2(new_n1170), .A3(new_n1090), .A4(new_n1092), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1094), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1147), .A2(KEYINPUT45), .A3(new_n997), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n830), .B(new_n1105), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n799), .B(new_n1127), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n748), .A2(new_n751), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n748), .A2(new_n751), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(G1986), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1181), .B1(new_n1182), .B2(new_n757), .ZN(new_n1183));
  NOR2_X1   g758(.A1(G290), .A2(G1986), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1173), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1172), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1173), .A2(new_n1184), .ZN(new_n1187));
  XOR2_X1   g762(.A(new_n1187), .B(KEYINPUT48), .Z(new_n1188));
  AOI21_X1  g763(.A(new_n1188), .B1(new_n1173), .B2(new_n1180), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1173), .A2(new_n1127), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT46), .ZN(new_n1191));
  OR3_X1    g766(.A1(new_n1190), .A2(KEYINPUT126), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1174), .A2(new_n800), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1193), .A2(new_n1173), .B1(KEYINPUT126), .B2(new_n1191), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1190), .B1(KEYINPUT126), .B2(new_n1191), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1192), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT47), .Z(new_n1197));
  OAI22_X1  g772(.A1(new_n1176), .A2(new_n1179), .B1(G2067), .B2(new_n830), .ZN(new_n1198));
  AOI211_X1 g773(.A(new_n1189), .B(new_n1197), .C1(new_n1173), .C2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1186), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g775(.A(G227), .ZN(new_n1202));
  OAI21_X1  g776(.A(new_n1202), .B1(new_n668), .B2(new_n669), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n1203), .B1(new_n906), .B2(new_n908), .ZN(new_n1204));
  NAND4_X1  g778(.A1(new_n980), .A2(G319), .A3(new_n703), .A4(new_n1204), .ZN(G225));
  NAND2_X1  g779(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1206));
  AOI21_X1  g780(.A(new_n460), .B1(new_n972), .B2(new_n979), .ZN(new_n1207));
  INV_X1    g781(.A(KEYINPUT127), .ZN(new_n1208));
  NAND4_X1  g782(.A1(new_n1207), .A2(new_n1208), .A3(new_n703), .A4(new_n1204), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n1206), .A2(new_n1209), .ZN(G308));
endmodule


