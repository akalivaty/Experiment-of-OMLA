//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT30), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(KEYINPUT22), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT25), .ZN(new_n213));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G169gat), .ZN(new_n222));
  INV_X1    g021(.A(G176gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT23), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n213), .B1(new_n221), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(KEYINPUT64), .B(new_n213), .C1(new_n221), .C2(new_n228), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n219), .A2(new_n220), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(G183gat), .A3(G190gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n236), .A3(new_n215), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  AND4_X1   g037(.A1(KEYINPUT25), .A2(new_n224), .A3(new_n226), .A4(new_n227), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n231), .A2(new_n232), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT27), .B(G183gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT28), .A3(new_n218), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT27), .B1(new_n217), .B2(KEYINPUT66), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT66), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT27), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(G183gat), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n244), .A2(new_n247), .A3(new_n218), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n243), .B1(new_n248), .B2(KEYINPUT28), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n222), .A2(new_n223), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT26), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n250), .A2(new_n251), .A3(new_n227), .ZN(new_n252));
  NOR2_X1   g051(.A1(G169gat), .A2(G176gat), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n253), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n252), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n255), .B1(new_n252), .B2(new_n254), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n249), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT29), .B1(new_n241), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G226gat), .A2(G233gat), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n261), .B(KEYINPUT71), .Z(new_n262));
  OAI21_X1  g061(.A(KEYINPUT73), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n262), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n264), .B1(new_n241), .B2(new_n259), .ZN(new_n265));
  AND3_X1   g064(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT25), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n240), .B1(new_n268), .B2(KEYINPUT64), .ZN(new_n269));
  INV_X1    g068(.A(new_n232), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n259), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT29), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n265), .B1(new_n273), .B2(new_n264), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n212), .B(new_n263), .C1(new_n274), .C2(KEYINPUT73), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n276));
  AOI22_X1  g075(.A1(new_n229), .A2(new_n230), .B1(new_n238), .B2(new_n239), .ZN(new_n277));
  INV_X1    g076(.A(new_n258), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n256), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n277), .A2(new_n232), .B1(new_n249), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n264), .B1(new_n280), .B2(KEYINPUT29), .ZN(new_n281));
  INV_X1    g080(.A(new_n265), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n212), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n276), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI211_X1 g084(.A(KEYINPUT72), .B(new_n212), .C1(new_n281), .C2(new_n282), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n205), .B(new_n275), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n204), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT72), .B1(new_n274), .B2(new_n212), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n283), .A2(new_n276), .A3(new_n284), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n289), .B1(new_n292), .B2(new_n275), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT74), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G1gat), .B(G29gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT0), .ZN(new_n296));
  XNOR2_X1  g095(.A(G57gat), .B(G85gat), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n296), .B(new_n297), .Z(new_n298));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n299));
  XOR2_X1   g098(.A(G127gat), .B(G134gat), .Z(new_n300));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n300), .B1(KEYINPUT1), .B2(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G113gat), .B(G120gat), .Z(new_n303));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304));
  XNOR2_X1  g103(.A(G127gat), .B(G134gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(G155gat), .B(G162gat), .Z(new_n308));
  OR2_X1    g107(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n309));
  NAND2_X1  g108(.A1(KEYINPUT76), .A2(KEYINPUT2), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G141gat), .B(G148gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n308), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314));
  INV_X1    g113(.A(G141gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(new_n315), .B2(G148gat), .ZN(new_n316));
  INV_X1    g115(.A(G148gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(KEYINPUT77), .A3(G141gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(G148gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  INV_X1    g120(.A(G155gat), .ZN(new_n322));
  INV_X1    g121(.A(G162gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(new_n324), .B2(KEYINPUT2), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n313), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n307), .A2(new_n327), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n313), .A2(new_n326), .A3(KEYINPUT78), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT78), .B1(new_n313), .B2(new_n326), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n328), .B1(new_n331), .B2(new_n307), .ZN(new_n332));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT79), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n327), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n315), .A2(G148gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n317), .A2(G141gat), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n309), .B(new_n310), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n339), .A2(new_n308), .B1(new_n320), .B2(new_n325), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT78), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n336), .A2(new_n341), .A3(KEYINPUT3), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n302), .A2(new_n306), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(new_n340), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n343), .A2(new_n347), .A3(new_n340), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT4), .B1(new_n307), .B2(new_n327), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n333), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n299), .B1(new_n334), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n341), .A3(new_n307), .ZN(new_n353));
  INV_X1    g152(.A(new_n328), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n356));
  INV_X1    g155(.A(new_n333), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n342), .A2(new_n345), .B1(new_n349), .B2(new_n348), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n358), .A2(KEYINPUT5), .B1(new_n359), .B2(new_n333), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n298), .B1(new_n352), .B2(new_n360), .ZN(new_n361));
  AOI211_X1 g160(.A(KEYINPUT79), .B(new_n333), .C1(new_n353), .C2(new_n354), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n351), .B1(new_n362), .B2(new_n299), .ZN(new_n363));
  INV_X1    g162(.A(new_n298), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n355), .A2(new_n357), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n365), .A2(KEYINPUT79), .B1(new_n359), .B2(new_n333), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n363), .B(new_n364), .C1(new_n366), .C2(new_n299), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n361), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n352), .A2(new_n360), .ZN(new_n370));
  INV_X1    g169(.A(new_n368), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n364), .A3(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n204), .B(new_n275), .C1(new_n285), .C2(new_n286), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT75), .B(KEYINPUT30), .ZN(new_n374));
  AOI22_X1  g173(.A1(new_n369), .A2(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n275), .B1(new_n285), .B2(new_n286), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n204), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT74), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n287), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n294), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT81), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT69), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n343), .B(new_n259), .C1(new_n269), .C2(new_n270), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT68), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n271), .A2(new_n307), .ZN(new_n385));
  NAND2_X1  g184(.A1(G227gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT68), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n241), .A2(new_n387), .A3(new_n343), .A4(new_n259), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n384), .A2(new_n385), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT34), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT32), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n384), .A2(new_n388), .A3(new_n385), .ZN(new_n394));
  INV_X1    g193(.A(new_n386), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT33), .B1(new_n394), .B2(new_n395), .ZN(new_n397));
  XOR2_X1   g196(.A(G15gat), .B(G43gat), .Z(new_n398));
  XNOR2_X1  g197(.A(G71gat), .B(G99gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n396), .A2(new_n397), .A3(new_n401), .ZN(new_n402));
  AOI221_X4 g201(.A(new_n393), .B1(KEYINPUT33), .B2(new_n400), .C1(new_n394), .C2(new_n395), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n382), .B(new_n392), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n394), .A2(new_n395), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT32), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT33), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(new_n408), .A3(new_n400), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n396), .B1(new_n397), .B2(new_n401), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n391), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n410), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n382), .B1(new_n413), .B2(new_n392), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n415), .B(G22gat), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  XOR2_X1   g216(.A(G78gat), .B(G106gat), .Z(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(G50gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT83), .ZN(new_n420));
  INV_X1    g219(.A(G228gat), .ZN(new_n421));
  INV_X1    g220(.A(G233gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT3), .B1(new_n212), .B2(new_n272), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n336), .A2(new_n341), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n340), .A2(new_n344), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n212), .B1(new_n427), .B2(new_n272), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n423), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n424), .A2(new_n340), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n431), .A2(new_n423), .A3(new_n428), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n420), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n430), .A2(new_n432), .A3(new_n420), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n417), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n435), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(new_n416), .A3(new_n433), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n412), .A2(new_n414), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT81), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n294), .A2(new_n375), .A3(new_n379), .A4(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n381), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n377), .A2(new_n287), .B1(new_n373), .B2(new_n374), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n369), .A2(new_n372), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT86), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT86), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n448), .A3(new_n445), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n392), .B1(new_n402), .B2(new_n403), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT70), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n411), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n413), .A2(KEYINPUT70), .A3(new_n392), .ZN(new_n454));
  AOI211_X1 g253(.A(KEYINPUT35), .B(new_n439), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n443), .A2(KEYINPUT35), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n369), .A2(new_n372), .A3(new_n373), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT37), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n292), .A2(new_n458), .A3(new_n275), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n284), .B(new_n263), .C1(new_n274), .C2(KEYINPUT73), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n460), .B(KEYINPUT37), .C1(new_n284), .C2(new_n274), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n461), .A3(new_n289), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT38), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n376), .B2(KEYINPUT37), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(new_n289), .A3(new_n459), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n457), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n439), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n359), .A2(new_n333), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT39), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n364), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n332), .A2(new_n333), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n472), .A2(KEYINPUT85), .A3(KEYINPUT39), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(new_n333), .B2(new_n359), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT85), .B1(new_n472), .B2(KEYINPUT39), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI211_X1 g277(.A(KEYINPUT40), .B(new_n471), .C1(new_n474), .C2(new_n475), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n478), .A2(new_n367), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n468), .B1(new_n444), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n467), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n381), .A2(new_n442), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n439), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n453), .A2(new_n454), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT36), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT36), .B1(new_n412), .B2(new_n414), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n482), .B1(new_n490), .B2(KEYINPUT84), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT84), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n484), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n456), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OR3_X1    g293(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(KEYINPUT91), .A3(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT88), .B(G29gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(G36gat), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n497), .B1(new_n499), .B2(KEYINPUT92), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT91), .B1(new_n495), .B2(new_n496), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT15), .ZN(new_n503));
  XOR2_X1   g302(.A(KEYINPUT89), .B(G43gat), .Z(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(G50gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT90), .B(G50gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(G43gat), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  OR2_X1    g307(.A1(G43gat), .A2(G50gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(G43gat), .A2(G50gat), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n511), .B1(new_n499), .B2(KEYINPUT92), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n502), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT87), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n496), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n496), .A2(new_n514), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n495), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n499), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n511), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT17), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT16), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n523), .B1(new_n524), .B2(G1gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT94), .ZN(new_n526));
  AOI21_X1  g325(.A(G8gat), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(new_n526), .B2(new_n525), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n523), .A2(G1gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n525), .A2(KEYINPUT93), .A3(G8gat), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n528), .B(new_n531), .C1(new_n529), .C2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n520), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n522), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n521), .A2(new_n533), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n536), .A2(KEYINPUT18), .A3(new_n537), .A4(new_n538), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n520), .B(new_n533), .Z(new_n543));
  XOR2_X1   g342(.A(new_n537), .B(KEYINPUT13), .Z(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n541), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(G197gat), .ZN(new_n548));
  XOR2_X1   g347(.A(KEYINPUT11), .B(G169gat), .Z(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT12), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n546), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n541), .A2(new_n553), .A3(new_n542), .A4(new_n545), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n494), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT96), .B(G57gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(G64gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT97), .ZN(new_n560));
  INV_X1    g359(.A(G64gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(G57gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G71gat), .B(G78gat), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n560), .B1(new_n559), .B2(new_n562), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n564), .A2(new_n569), .ZN(new_n571));
  XNOR2_X1  g370(.A(G57gat), .B(G64gat), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n571), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  OAI22_X1  g372(.A1(new_n567), .A2(new_n568), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT21), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G127gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n574), .B(KEYINPUT98), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n533), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n580), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G155gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n584), .A2(new_n588), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT7), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G99gat), .B(G106gat), .Z(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n522), .A2(new_n535), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  AND2_X1   g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n520), .A2(new_n602), .B1(KEYINPUT41), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT100), .ZN(new_n606));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT99), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n605), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G134gat), .B(G162gat), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n606), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n611), .A2(new_n616), .A3(new_n612), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n591), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g421(.A1(new_n574), .A2(KEYINPUT101), .A3(new_n600), .ZN(new_n623));
  AOI21_X1  g422(.A(KEYINPUT101), .B1(new_n574), .B2(new_n600), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n599), .A2(KEYINPUT102), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n598), .B(new_n626), .Z(new_n627));
  OR2_X1    g426(.A1(new_n574), .A2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT105), .ZN(new_n634));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n581), .A2(KEYINPUT10), .A3(new_n602), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n639), .B(new_n628), .C1(new_n623), .C2(new_n624), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n641), .A2(new_n642), .B1(G230gat), .B2(G233gat), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n638), .A2(KEYINPUT103), .A3(new_n640), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n643), .A2(KEYINPUT104), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT104), .B1(new_n643), .B2(new_n644), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n632), .B(new_n637), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n641), .A2(new_n630), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n637), .B1(new_n632), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n622), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT106), .Z(new_n654));
  NAND2_X1  g453(.A1(new_n557), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n445), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(G1gat), .Z(G1324gat));
  INV_X1    g456(.A(KEYINPUT42), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n655), .A2(new_n444), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  AOI21_X1  g459(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(G8gat), .B1(new_n655), .B2(new_n444), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(KEYINPUT107), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n664), .B1(new_n660), .B2(new_n665), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n661), .A2(new_n662), .B1(new_n659), .B2(new_n666), .ZN(G1325gat));
  OAI21_X1  g466(.A(G15gat), .B1(new_n655), .B2(new_n489), .ZN(new_n668));
  INV_X1    g467(.A(new_n485), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n669), .A2(G15gat), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n668), .B1(new_n655), .B2(new_n670), .ZN(G1326gat));
  NOR3_X1   g470(.A1(new_n494), .A2(new_n556), .A3(new_n468), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n654), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  AOI21_X1  g474(.A(new_n468), .B1(new_n381), .B2(new_n442), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n487), .A2(new_n488), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT84), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n482), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n493), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n443), .A2(KEYINPUT35), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n450), .A2(new_n455), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n620), .B1(new_n680), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n589), .A2(new_n590), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n651), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n556), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n445), .ZN(new_n690));
  INV_X1    g489(.A(new_n498), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT45), .ZN(new_n693));
  INV_X1    g492(.A(new_n688), .ZN(new_n694));
  OAI21_X1  g493(.A(KEYINPUT44), .B1(new_n494), .B2(new_n620), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n676), .A2(new_n677), .A3(new_n482), .ZN(new_n697));
  OAI211_X1 g496(.A(new_n696), .B(new_n621), .C1(new_n697), .C2(new_n456), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n484), .A2(new_n489), .A3(new_n679), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n683), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n702), .A2(KEYINPUT108), .A3(new_n696), .A4(new_n621), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n694), .B1(new_n695), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n498), .B1(new_n706), .B2(new_n445), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n693), .A2(new_n707), .ZN(G1328gat));
  INV_X1    g507(.A(G36gat), .ZN(new_n709));
  INV_X1    g508(.A(new_n444), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n689), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT46), .Z(new_n712));
  OAI21_X1  g511(.A(G36gat), .B1(new_n706), .B2(new_n444), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1329gat));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n689), .A2(new_n504), .A3(new_n485), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n504), .B1(new_n705), .B2(new_n677), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n717), .B2(KEYINPUT109), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n700), .A2(new_n703), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n684), .A2(new_n696), .ZN(new_n720));
  OAI211_X1 g519(.A(new_n677), .B(new_n688), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n504), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n721), .A2(KEYINPUT109), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n715), .B1(new_n718), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n716), .A2(KEYINPUT47), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n504), .B1(new_n721), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n704), .B1(new_n696), .B2(new_n684), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n728), .A2(KEYINPUT110), .A3(new_n677), .A4(new_n688), .ZN(new_n729));
  AOI211_X1 g528(.A(KEYINPUT111), .B(new_n725), .C1(new_n727), .C2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n721), .A2(new_n726), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(new_n722), .A3(new_n729), .ZN(new_n733));
  INV_X1    g532(.A(new_n725), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n724), .B1(new_n730), .B2(new_n735), .ZN(G1330gat));
  NAND4_X1  g535(.A1(new_n672), .A2(new_n506), .A3(new_n621), .A4(new_n686), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n706), .A2(new_n468), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(new_n506), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT48), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g540(.A(KEYINPUT48), .B(new_n737), .C1(new_n738), .C2(new_n506), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1331gat));
  AND4_X1   g542(.A1(new_n556), .A2(new_n702), .A3(new_n622), .A4(new_n651), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n690), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(new_n558), .Z(G1332gat));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n710), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT49), .B(G64gat), .Z(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(G1333gat));
  NAND2_X1  g549(.A1(new_n744), .A2(new_n677), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n669), .A2(G71gat), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n751), .A2(G71gat), .B1(new_n744), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g553(.A1(new_n744), .A2(new_n439), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g555(.A1(new_n685), .A2(new_n555), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n702), .A2(new_n621), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n758), .A2(new_n759), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n652), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n595), .A3(new_n690), .ZN(new_n764));
  INV_X1    g563(.A(new_n728), .ZN(new_n765));
  INV_X1    g564(.A(new_n757), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n652), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n765), .A2(new_n445), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n764), .B1(new_n769), .B2(new_n595), .ZN(G1336gat));
  NAND3_X1  g569(.A1(new_n728), .A2(new_n710), .A3(new_n767), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n771), .A2(new_n772), .A3(G92gat), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n771), .B2(G92gat), .ZN(new_n774));
  NOR4_X1   g573(.A1(new_n762), .A2(G92gat), .A3(new_n444), .A4(new_n652), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777));
  XNOR2_X1  g576(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n771), .A2(G92gat), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n776), .A2(new_n777), .B1(new_n779), .B2(new_n780), .ZN(G1337gat));
  INV_X1    g580(.A(G99gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n782), .A3(new_n485), .ZN(new_n783));
  NOR3_X1   g582(.A1(new_n765), .A2(new_n489), .A3(new_n768), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n782), .ZN(G1338gat));
  OAI211_X1 g584(.A(new_n439), .B(new_n651), .C1(new_n760), .C2(new_n761), .ZN(new_n786));
  INV_X1    g585(.A(G106gat), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n765), .A2(new_n768), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n468), .A2(new_n787), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(KEYINPUT53), .B1(new_n791), .B2(KEYINPUT114), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n789), .A2(new_n790), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n793), .B(new_n794), .C1(new_n795), .C2(new_n788), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n792), .A2(new_n796), .ZN(G1339gat));
  OAI21_X1  g596(.A(new_n636), .B1(new_n648), .B2(KEYINPUT54), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n798), .B(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT54), .B1(new_n641), .B2(new_n630), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n645), .B2(new_n646), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n800), .A2(new_n803), .A3(KEYINPUT55), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(new_n647), .A3(new_n555), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  INV_X1    g605(.A(new_n646), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n643), .A2(KEYINPUT104), .A3(new_n644), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n801), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n798), .B(KEYINPUT115), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(KEYINPUT116), .B(new_n806), .C1(new_n809), .C2(new_n810), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n805), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n543), .A2(new_n544), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n550), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n554), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n632), .A2(new_n637), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n807), .B2(new_n808), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n821), .B2(new_n649), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n620), .B1(new_n815), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n813), .A2(new_n814), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n621), .A2(new_n819), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n825), .A2(new_n826), .A3(new_n647), .A4(new_n804), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n685), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n653), .A2(new_n555), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(new_n439), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n444), .A2(new_n690), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n669), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(G113gat), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n834), .A2(new_n835), .A3(new_n556), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n830), .A2(new_n445), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n440), .A2(new_n444), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n555), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n836), .B1(new_n835), .B2(new_n841), .ZN(G1340gat));
  INV_X1    g641(.A(G120gat), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n834), .A2(new_n843), .A3(new_n652), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n651), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n843), .B2(new_n845), .ZN(G1341gat));
  OAI21_X1  g645(.A(new_n579), .B1(new_n839), .B2(new_n591), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n685), .A2(G127gat), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT117), .B1(new_n834), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n834), .A2(KEYINPUT117), .A3(new_n848), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(G1342gat));
  NOR2_X1   g651(.A1(new_n620), .A2(G134gat), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT56), .B1(new_n839), .B2(new_n854), .ZN(new_n855));
  OR3_X1    g654(.A1(new_n839), .A2(KEYINPUT56), .A3(new_n854), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n831), .A2(new_n621), .A3(new_n833), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(KEYINPUT118), .A3(G134gat), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT118), .B1(new_n857), .B2(G134gat), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n855), .B(new_n856), .C1(new_n859), .C2(new_n860), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n677), .A2(new_n468), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n710), .ZN(new_n864));
  AND4_X1   g663(.A1(new_n315), .A2(new_n837), .A3(new_n555), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(KEYINPUT58), .ZN(new_n866));
  AND4_X1   g665(.A1(new_n555), .A2(new_n811), .A3(new_n647), .A4(new_n804), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n822), .A2(KEYINPUT119), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n651), .A2(new_n869), .A3(new_n819), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n620), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n685), .B1(new_n872), .B2(new_n827), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n439), .B1(new_n873), .B2(new_n829), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(KEYINPUT57), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n876), .B(new_n439), .C1(new_n828), .C2(new_n829), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n677), .A2(new_n832), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n875), .A2(new_n877), .A3(new_n555), .A4(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G141gat), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n879), .A2(new_n880), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n866), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n879), .A2(new_n885), .A3(G141gat), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n885), .B1(new_n879), .B2(G141gat), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n886), .A2(new_n887), .A3(new_n865), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(G1344gat));
  NAND2_X1  g689(.A1(new_n837), .A2(new_n864), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n317), .A3(new_n651), .ZN(new_n893));
  XNOR2_X1  g692(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n654), .A2(new_n556), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n876), .B(new_n439), .C1(new_n895), .C2(new_n873), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT57), .B1(new_n830), .B2(new_n468), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n896), .A2(new_n651), .A3(new_n878), .A4(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n894), .B1(new_n898), .B2(G148gat), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n652), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(KEYINPUT59), .A3(new_n317), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n893), .B1(new_n899), .B2(new_n902), .ZN(G1345gat));
  OAI21_X1  g702(.A(G155gat), .B1(new_n900), .B2(new_n591), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n685), .A2(new_n322), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n891), .B2(new_n905), .ZN(G1346gat));
  NOR3_X1   g705(.A1(new_n891), .A2(G162gat), .A3(new_n620), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n907), .B(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G162gat), .B1(new_n900), .B2(new_n620), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1347gat));
  NAND2_X1  g710(.A1(new_n710), .A2(new_n445), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n669), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n468), .B(new_n913), .C1(new_n828), .C2(new_n829), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n914), .A2(new_n222), .A3(new_n556), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n830), .A2(new_n690), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n440), .A2(new_n710), .ZN(new_n917));
  XOR2_X1   g716(.A(new_n917), .B(KEYINPUT124), .Z(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n555), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n915), .B1(new_n921), .B2(new_n222), .ZN(G1348gat));
  OAI21_X1  g721(.A(G176gat), .B1(new_n914), .B2(new_n652), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n651), .A2(new_n223), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n919), .B2(new_n924), .ZN(G1349gat));
  OAI21_X1  g724(.A(G183gat), .B1(new_n914), .B2(new_n591), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n685), .A2(new_n242), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n919), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n914), .B2(new_n620), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n930), .B(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n920), .A2(new_n218), .A3(new_n621), .ZN(new_n935));
  XNOR2_X1  g734(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n934), .B(new_n935), .C1(new_n932), .C2(new_n936), .ZN(G1351gat));
  NOR2_X1   g736(.A1(new_n863), .A2(new_n444), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n916), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g739(.A(G197gat), .B1(new_n940), .B2(new_n555), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n896), .A2(new_n897), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n677), .A2(new_n912), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n555), .A2(G197gat), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n941), .B1(new_n945), .B2(new_n946), .ZN(G1352gat));
  OAI21_X1  g746(.A(G204gat), .B1(new_n944), .B2(new_n652), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n652), .A2(G204gat), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n939), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT62), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n948), .A2(new_n951), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n940), .A2(new_n207), .A3(new_n685), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n896), .A2(new_n685), .A3(new_n897), .A4(new_n943), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1354gat));
  AOI21_X1  g756(.A(G218gat), .B1(new_n940), .B2(new_n621), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n620), .A2(new_n208), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT127), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n958), .B1(new_n945), .B2(new_n960), .ZN(G1355gat));
endmodule


