//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n565, new_n566, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n458), .A2(KEYINPUT66), .ZN(new_n459));
  AOI22_X1  g034(.A1(new_n458), .A2(KEYINPUT66), .B1(G567), .B2(new_n454), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT67), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n478), .B1(new_n466), .B2(G2104), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n464), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n479), .A2(new_n467), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(G137), .A3(new_n475), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n464), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G101), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n483), .A2(KEYINPUT69), .A3(G101), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n477), .A2(new_n482), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G160));
  NAND3_X1  g065(.A1(new_n479), .A2(new_n467), .A3(new_n480), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G136), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n475), .A2(G112), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n476), .A2(new_n481), .ZN(new_n497));
  INV_X1    g072(.A(G124), .ZN(new_n498));
  OR3_X1    g073(.A1(new_n497), .A2(KEYINPUT70), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT70), .B1(new_n497), .B2(new_n498), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n499), .B2(new_n500), .ZN(G162));
  AND2_X1   g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n479), .A2(new_n480), .A3(new_n467), .A4(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT71), .B1(new_n471), .B2(G114), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  INV_X1    g082(.A(G114), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(G2105), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n506), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT72), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n505), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n507), .B1(new_n508), .B2(G2105), .ZN(new_n513));
  NOR3_X1   g088(.A1(new_n471), .A2(KEYINPUT71), .A3(G114), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(new_n503), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n472), .A2(new_n474), .A3(G138), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT4), .B1(new_n491), .B2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT3), .B(G2104), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n475), .A2(new_n520), .A3(new_n521), .A4(G138), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n511), .A2(new_n517), .B1(new_n519), .B2(new_n522), .ZN(G164));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(G50), .A3(G543), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT73), .ZN(new_n526));
  INV_X1    g101(.A(G88), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT74), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n529), .B2(KEYINPUT5), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT5), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n531), .A2(KEYINPUT74), .A3(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n529), .A2(KEYINPUT5), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(new_n524), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n526), .B1(new_n527), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n535), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G651), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n537), .A2(new_n540), .ZN(G166));
  INV_X1    g116(.A(new_n536), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n542), .A2(G89), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n535), .A2(G63), .A3(G651), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT7), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n524), .A2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G51), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n543), .A2(new_n549), .ZN(G168));
  AOI22_X1  g125(.A1(new_n535), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n539), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n547), .A2(G52), .ZN(new_n553));
  INV_X1    g128(.A(G90), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n536), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(G171));
  AOI22_X1  g131(.A1(new_n535), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n539), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n547), .A2(G43), .ZN(new_n559));
  INV_X1    g134(.A(G81), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n536), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  AOI22_X1  g142(.A1(new_n535), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n539), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n542), .A2(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n547), .A2(G53), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT9), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  OR2_X1    g150(.A1(new_n537), .A2(new_n540), .ZN(G303));
  NAND3_X1  g151(.A1(new_n547), .A2(KEYINPUT75), .A3(G49), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n524), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n535), .A2(G87), .A3(new_n524), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n535), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  NAND3_X1  g160(.A1(new_n533), .A2(G61), .A3(new_n534), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(KEYINPUT76), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n588));
  NAND4_X1  g163(.A1(new_n533), .A2(new_n588), .A3(G61), .A4(new_n534), .ZN(new_n589));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n535), .A2(G86), .A3(new_n524), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n547), .A2(G48), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n592), .A2(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n542), .A2(G85), .B1(G47), .B2(new_n547), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n535), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n539), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n535), .A2(G92), .A3(new_n524), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n535), .A2(G66), .ZN(new_n604));
  INV_X1    g179(.A(G79), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n529), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n606), .A2(G651), .B1(new_n547), .B2(G54), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G868), .ZN(G284));
  XNOR2_X1  g185(.A(G284), .B(KEYINPUT77), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT78), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n614));
  AOI21_X1  g189(.A(G868), .B1(G299), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n614), .B2(G299), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n613), .A2(new_n616), .ZN(G297));
  XNOR2_X1  g192(.A(G297), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n609), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n609), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(KEYINPUT81), .A2(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n520), .A2(new_n483), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  NOR2_X1   g203(.A1(KEYINPUT81), .A2(G2100), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n625), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n492), .A2(G135), .ZN(new_n631));
  OAI221_X1 g206(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n475), .C2(G111), .ZN(new_n632));
  INV_X1    g207(.A(G123), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n497), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT82), .B(G2096), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n630), .B(new_n636), .C1(new_n628), .C2(new_n625), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2438), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2430), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(KEYINPUT14), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT84), .Z(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n639), .B2(new_n641), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n651), .A2(new_n654), .A3(new_n652), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(new_n657), .A3(G14), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT85), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT17), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2084), .B(G2090), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n664), .B1(new_n661), .B2(new_n663), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n662), .B2(new_n663), .ZN(new_n667));
  INV_X1    g242(.A(new_n663), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n668), .A2(new_n664), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n661), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n665), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2096), .B(G2100), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  AND2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  NOR3_X1   g258(.A1(new_n677), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n677), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT86), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1981), .B(G1986), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G35), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT101), .Z(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G162), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT102), .B(KEYINPUT29), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G2090), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT31), .B(G11), .Z(new_n701));
  NOR2_X1   g276(.A1(new_n634), .A2(new_n694), .ZN(new_n702));
  INV_X1    g277(.A(G28), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(KEYINPUT30), .ZN(new_n704));
  AOI21_X1  g279(.A(G29), .B1(new_n703), .B2(KEYINPUT30), .ZN(new_n705));
  AOI211_X1 g280(.A(new_n701), .B(new_n702), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G16), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G21), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G168), .B2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT99), .B(G1966), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n708), .B(new_n710), .C1(G168), .C2(new_n707), .ZN(new_n713));
  AND4_X1   g288(.A1(new_n700), .A2(new_n706), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n707), .A2(G5), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G301), .B2(G16), .ZN(new_n716));
  INV_X1    g291(.A(G1961), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(G16), .A2(G19), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n562), .B2(G16), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT90), .B(G1341), .Z(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n718), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n694), .A2(G26), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT28), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n492), .A2(G140), .ZN(new_n727));
  OAI221_X1 g302(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n475), .C2(G116), .ZN(new_n728));
  INV_X1    g303(.A(G128), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n727), .B(new_n728), .C1(new_n729), .C2(new_n497), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n726), .B1(new_n730), .B2(G29), .ZN(new_n731));
  INV_X1    g306(.A(G2067), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n699), .B2(new_n697), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n694), .A2(G27), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G164), .B2(new_n694), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(G2078), .Z(new_n737));
  NAND4_X1  g312(.A1(new_n714), .A2(new_n724), .A3(new_n734), .A4(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G34), .ZN(new_n739));
  AND2_X1   g314(.A1(new_n739), .A2(KEYINPUT24), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n739), .A2(KEYINPUT24), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n694), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G160), .B2(new_n694), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT95), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G2084), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT96), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  INV_X1    g323(.A(G2072), .ZN(new_n749));
  OR2_X1    g324(.A1(G29), .A2(G33), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT91), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(KEYINPUT25), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n751), .A2(KEYINPUT91), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT25), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n751), .A2(KEYINPUT91), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n753), .A2(new_n757), .B1(G139), .B2(new_n492), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n520), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT92), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n476), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n760), .B2(new_n759), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(KEYINPUT93), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(KEYINPUT93), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n758), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n750), .B1(new_n765), .B2(new_n694), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n748), .B1(new_n749), .B2(new_n766), .ZN(new_n767));
  NOR3_X1   g342(.A1(new_n738), .A2(new_n747), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n749), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT94), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(KEYINPUT94), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT100), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n716), .A2(new_n717), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n694), .A2(G32), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n492), .A2(G141), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT26), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n778), .A2(new_n779), .B1(G105), .B2(new_n483), .ZN(new_n780));
  INV_X1    g355(.A(G129), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n775), .B(new_n780), .C1(new_n781), .C2(new_n497), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n774), .B1(new_n783), .B2(new_n694), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT97), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT27), .B(G1996), .ZN(new_n786));
  OAI221_X1 g361(.A(new_n773), .B1(new_n744), .B2(G2084), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n770), .A2(new_n771), .B1(new_n772), .B2(new_n787), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n787), .A2(new_n772), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT103), .B(KEYINPUT23), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n707), .A2(G20), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G299), .B2(G16), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1956), .ZN(new_n794));
  OR2_X1    g369(.A1(G4), .A2(G16), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n608), .B2(new_n707), .ZN(new_n796));
  INV_X1    g371(.A(G1348), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n794), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT98), .ZN(new_n801));
  AND3_X1   g376(.A1(new_n785), .A2(new_n801), .A3(new_n786), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n801), .B1(new_n785), .B2(new_n786), .ZN(new_n803));
  NOR3_X1   g378(.A1(new_n800), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n768), .A2(new_n788), .A3(new_n789), .A4(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(G1971), .ZN(new_n806));
  NAND2_X1  g381(.A1(G303), .A2(G16), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT89), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n707), .A2(G22), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n807), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n808), .B1(new_n807), .B2(new_n809), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n806), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n812), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n814), .A2(G1971), .A3(new_n810), .ZN(new_n815));
  INV_X1    g390(.A(G305), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(G16), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G6), .B2(G16), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT32), .B(G1981), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n813), .A2(new_n815), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n707), .A2(G23), .ZN(new_n823));
  INV_X1    g398(.A(G288), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(new_n707), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT33), .B(G1976), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n825), .B(new_n826), .Z(new_n827));
  NOR2_X1   g402(.A1(new_n818), .A2(new_n820), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(KEYINPUT34), .B1(new_n822), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n814), .A2(new_n810), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n832), .A2(new_n806), .B1(new_n818), .B2(new_n820), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT34), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n833), .A2(new_n829), .A3(new_n834), .A4(new_n815), .ZN(new_n835));
  MUX2_X1   g410(.A(G24), .B(G290), .S(G16), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1986), .ZN(new_n837));
  INV_X1    g412(.A(G25), .ZN(new_n838));
  OR3_X1    g413(.A1(new_n838), .A2(KEYINPUT87), .A3(G29), .ZN(new_n839));
  OAI21_X1  g414(.A(KEYINPUT87), .B1(new_n838), .B2(G29), .ZN(new_n840));
  OAI221_X1 g415(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n475), .C2(G107), .ZN(new_n841));
  INV_X1    g416(.A(G119), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n497), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(G131), .B2(new_n492), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n839), .B(new_n840), .C1(new_n844), .C2(new_n694), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT35), .B(G1991), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT88), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n837), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n831), .A2(new_n835), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT36), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT36), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n831), .A2(new_n835), .A3(new_n852), .A4(new_n849), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n805), .B1(new_n851), .B2(new_n853), .ZN(G311));
  NOR2_X1   g429(.A1(G311), .A2(KEYINPUT104), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n856));
  AOI211_X1 g431(.A(new_n856), .B(new_n805), .C1(new_n851), .C2(new_n853), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n857), .ZN(G150));
  NAND2_X1  g433(.A1(new_n547), .A2(G55), .ZN(new_n859));
  INV_X1    g434(.A(G93), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(new_n536), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n535), .A2(G67), .ZN(new_n862));
  NAND2_X1  g437(.A1(G80), .A2(G543), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n539), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G860), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT37), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n609), .A2(G559), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n562), .A2(new_n865), .ZN(new_n871));
  OAI22_X1  g446(.A1(new_n558), .A2(new_n561), .B1(new_n861), .B2(new_n864), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n870), .B(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT105), .Z(new_n877));
  OAI21_X1  g452(.A(new_n866), .B1(new_n874), .B2(new_n875), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n868), .B1(new_n877), .B2(new_n878), .ZN(G145));
  XNOR2_X1  g454(.A(G160), .B(new_n634), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(G162), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT106), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n765), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n883), .B1(new_n765), .B2(new_n884), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n730), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  INV_X1    g464(.A(new_n730), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n885), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n891), .A3(new_n782), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n782), .B1(new_n888), .B2(new_n891), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n492), .A2(G142), .ZN(new_n895));
  OAI221_X1 g470(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n475), .C2(G118), .ZN(new_n896));
  INV_X1    g471(.A(G130), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n497), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(new_n627), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(new_n844), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n519), .A2(new_n522), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n504), .A2(new_n510), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n900), .B(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n893), .A2(new_n894), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n888), .A2(new_n891), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n783), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n904), .B1(new_n908), .B2(new_n892), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n882), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G37), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n905), .B1(new_n893), .B2(new_n894), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n908), .A2(new_n904), .A3(new_n892), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n913), .A3(new_n881), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n910), .A2(new_n911), .A3(new_n914), .A4(new_n916), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(G395));
  INV_X1    g495(.A(G868), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n861), .B2(new_n864), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n621), .B(new_n873), .Z(new_n923));
  NAND2_X1  g498(.A1(new_n608), .A2(G299), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n572), .A2(new_n570), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n925), .A2(new_n569), .A3(new_n603), .A4(new_n607), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT41), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n924), .A2(KEYINPUT41), .A3(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n926), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n816), .B(G166), .ZN(new_n932));
  XNOR2_X1  g507(.A(G290), .B(new_n824), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n932), .B(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n934), .B(KEYINPUT42), .Z(new_n935));
  OAI221_X1 g510(.A(new_n929), .B1(new_n931), .B2(new_n923), .C1(new_n935), .C2(KEYINPUT109), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(KEYINPUT109), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n929), .B1(new_n931), .B2(new_n923), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n936), .A2(new_n939), .B1(KEYINPUT109), .B2(new_n935), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n922), .B1(new_n940), .B2(new_n921), .ZN(G295));
  OAI21_X1  g516(.A(new_n922), .B1(new_n940), .B2(new_n921), .ZN(G331));
  AOI21_X1  g517(.A(G301), .B1(new_n871), .B2(new_n872), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n871), .A2(G301), .A3(new_n872), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(G168), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n945), .ZN(new_n947));
  OAI21_X1  g522(.A(G286), .B1(new_n947), .B2(new_n943), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n931), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n928), .A2(new_n927), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n946), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n934), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT43), .ZN(new_n955));
  INV_X1    g530(.A(new_n934), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n950), .A2(new_n952), .A3(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n911), .A4(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT110), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT44), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n954), .A2(new_n911), .A3(new_n957), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n958), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n959), .A2(new_n962), .A3(KEYINPUT44), .A4(new_n958), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(G397));
  INV_X1    g541(.A(KEYINPUT122), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT111), .B(G40), .Z(new_n968));
  AND4_X1   g543(.A1(new_n477), .A2(new_n482), .A3(new_n488), .A4(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n901), .B2(new_n902), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT119), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n515), .A2(new_n516), .A3(new_n503), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n516), .B1(new_n515), .B2(new_n503), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n901), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1384), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n977), .A2(new_n971), .A3(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT119), .B(new_n969), .C1(new_n970), .C2(new_n971), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n974), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1956), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(G164), .B2(G1384), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n477), .A2(new_n482), .A3(new_n488), .A4(new_n968), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(new_n970), .B2(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT56), .B(G2072), .ZN(new_n989));
  AOI22_X1  g564(.A1(new_n981), .A2(new_n982), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT57), .ZN(new_n991));
  XNOR2_X1  g566(.A(G299), .B(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n967), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT61), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n990), .B2(new_n992), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n980), .A2(new_n979), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n515), .A2(new_n503), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n519), .B2(new_n522), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT50), .B1(new_n998), .B2(G1384), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT119), .B1(new_n999), .B2(new_n969), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n982), .B1(new_n996), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n984), .A2(new_n986), .A3(new_n989), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(G299), .B(KEYINPUT57), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(KEYINPUT122), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n993), .A2(new_n995), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n992), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n994), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n969), .A2(new_n970), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT58), .B(G1341), .Z(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n987), .B2(G1996), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n562), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT59), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1006), .A2(new_n1009), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1017), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n465), .A2(new_n467), .A3(new_n521), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n518), .A2(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n472), .A2(new_n474), .A3(G138), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n480), .A2(new_n467), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(new_n479), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n1023), .B2(KEYINPUT4), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n971), .B(new_n978), .C1(new_n1024), .C2(new_n997), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT116), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n971), .B1(new_n977), .B2(new_n978), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1018), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n969), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n797), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n969), .A2(new_n970), .A3(new_n732), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT60), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n609), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1030), .A2(KEYINPUT60), .A3(new_n608), .A4(new_n1031), .ZN(new_n1035));
  AOI22_X1  g610(.A1(new_n1034), .A2(new_n1035), .B1(new_n1033), .B2(new_n1032), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1032), .A2(new_n609), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1037), .A2(new_n993), .A3(new_n1005), .ZN(new_n1038));
  OAI22_X1  g613(.A1(new_n1016), .A2(new_n1036), .B1(new_n1038), .B2(new_n1007), .ZN(new_n1039));
  INV_X1    g614(.A(G2084), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1028), .A2(new_n1040), .A3(new_n969), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT120), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n977), .A2(new_n1042), .A3(KEYINPUT45), .A4(new_n978), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n983), .B1(new_n998), .B2(G1384), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n969), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n511), .A2(new_n517), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1384), .B1(new_n1046), .B2(new_n901), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1042), .B1(new_n1047), .B2(KEYINPUT45), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n710), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1041), .A2(G168), .A3(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(G8), .ZN(new_n1051));
  AOI21_X1  g626(.A(G168), .B1(new_n1041), .B2(new_n1049), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT51), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1050), .A2(new_n1054), .A3(G8), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1029), .A2(new_n717), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n987), .B2(G2078), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  XOR2_X1   g636(.A(G171), .B(KEYINPUT54), .Z(new_n1062));
  NAND3_X1  g637(.A1(new_n903), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1044), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT124), .B(G2078), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1064), .A2(new_n489), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1062), .B1(new_n1063), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1061), .A2(new_n1068), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1045), .A2(new_n1048), .A3(G2078), .ZN(new_n1070));
  OR2_X1    g645(.A1(new_n1070), .A2(KEYINPUT123), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1058), .B1(new_n1070), .B2(KEYINPUT123), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1060), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1062), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1069), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1056), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n1078));
  INV_X1    g653(.A(G8), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1078), .B1(G166), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1063), .A2(new_n969), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT45), .B1(new_n977), .B2(new_n978), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n806), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1971), .B1(new_n984), .B2(new_n986), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT115), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G2090), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1028), .A2(new_n1090), .A3(new_n969), .ZN(new_n1091));
  OAI211_X1 g666(.A(G8), .B(new_n1081), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n996), .A2(new_n1000), .A3(G2090), .ZN(new_n1093));
  OAI21_X1  g668(.A(G8), .B1(new_n1093), .B2(new_n1087), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1081), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1010), .A2(G8), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n592), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(G305), .A2(new_n1099), .A3(G1981), .ZN(new_n1100));
  INV_X1    g675(.A(G1981), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n592), .B(new_n595), .C1(new_n1098), .C2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT49), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1097), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1100), .A2(KEYINPUT49), .A3(new_n1102), .ZN(new_n1106));
  INV_X1    g681(.A(G1976), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1010), .B(G8), .C1(new_n1107), .C2(G288), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT52), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1108), .A2(new_n1110), .B1(G288), .B2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g688(.A1(new_n1105), .A2(new_n1106), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1092), .A2(new_n1096), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1092), .A2(new_n1096), .A3(new_n1114), .A4(KEYINPUT125), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1039), .A2(new_n1076), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1053), .A2(new_n1121), .A3(new_n1055), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1121), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1125));
  AOI21_X1  g700(.A(G301), .B1(new_n1125), .B2(new_n1061), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1117), .A2(new_n1118), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1041), .A2(new_n1049), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(G8), .A3(G168), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1115), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(KEYINPUT121), .B(new_n1129), .C1(new_n1115), .C2(new_n1131), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1114), .A2(KEYINPUT63), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1136), .A2(new_n1131), .ZN(new_n1137));
  OAI21_X1  g712(.A(G8), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1095), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1137), .A2(new_n1092), .A3(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1134), .A2(new_n1135), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1142), .A2(new_n1107), .A3(new_n824), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(G1981), .B2(G305), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1097), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1092), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1144), .A2(new_n1145), .B1(new_n1146), .B2(new_n1114), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1120), .A2(new_n1128), .A3(new_n1141), .A4(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1044), .A2(new_n985), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(G290), .A2(G1986), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT112), .ZN(new_n1152));
  NAND2_X1  g727(.A1(G290), .A2(G1986), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1150), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT113), .Z(new_n1155));
  XNOR2_X1  g730(.A(new_n730), .B(new_n732), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n782), .B(G1996), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1149), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(new_n1159), .B(KEYINPUT114), .Z(new_n1160));
  INV_X1    g735(.A(new_n847), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n844), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n844), .A2(new_n1161), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1150), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1155), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1148), .A2(new_n1166), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1165), .A2(KEYINPUT126), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1165), .A2(KEYINPUT126), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1152), .A2(new_n1150), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1170), .B(KEYINPUT48), .Z(new_n1171));
  NAND3_X1  g746(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1149), .B1(new_n1157), .B2(new_n782), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1150), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT46), .ZN(new_n1175));
  INV_X1    g750(.A(G1996), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1175), .B1(new_n1149), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1173), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT47), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n730), .A2(G2067), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1149), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1172), .A2(new_n1179), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1167), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g759(.A1(G229), .A2(new_n461), .A3(G227), .ZN(new_n1186));
  AND2_X1   g760(.A1(new_n658), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g761(.A1(new_n1187), .A2(new_n915), .A3(new_n963), .ZN(G225));
  INV_X1    g762(.A(G225), .ZN(G308));
endmodule


