//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n563, new_n564,
    new_n565, new_n566, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1227, new_n1228;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT65), .Z(G319));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n464));
  AND3_X1   g039(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n465), .A2(KEYINPUT68), .A3(G137), .A4(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n461), .A2(new_n463), .A3(new_n466), .A4(new_n464), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n460), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n467), .A2(new_n471), .B1(G101), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n475), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n476), .B2(new_n466), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n462), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n464), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n473), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT69), .ZN(G160));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n461), .A2(new_n463), .A3(G2105), .A4(new_n464), .ZN(new_n489));
  INV_X1    g064(.A(G124), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n469), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G136), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT70), .ZN(G162));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n461), .A2(new_n463), .A3(new_n496), .A4(new_n464), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n495), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n497), .A2(KEYINPUT4), .B1(new_n475), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(G114), .B2(new_n466), .ZN(new_n502));
  INV_X1    g077(.A(G126), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n489), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n499), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  XOR2_X1   g085(.A(new_n510), .B(KEYINPUT71), .Z(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  OAI21_X1  g088(.A(G543), .B1(new_n513), .B2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(KEYINPUT72), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n517), .A2(new_n513), .A3(KEYINPUT5), .A4(G543), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(new_n518), .B1(new_n507), .B2(new_n508), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n511), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n516), .A2(new_n518), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n521), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT75), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT75), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n507), .A2(new_n508), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G543), .B1(new_n517), .B2(KEYINPUT5), .ZN(new_n536));
  INV_X1    g111(.A(new_n518), .ZN(new_n537));
  OAI211_X1 g112(.A(G89), .B(new_n534), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n529), .A2(KEYINPUT7), .A3(new_n530), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n533), .A2(new_n538), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n509), .A2(G51), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(G63), .A2(G651), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n516), .B2(new_n518), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n542), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n536), .A2(new_n537), .ZN(new_n548));
  OAI211_X1 g123(.A(KEYINPUT74), .B(new_n543), .C1(new_n548), .C2(new_n545), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n541), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n540), .ZN(new_n551));
  AOI21_X1  g126(.A(KEYINPUT7), .B1(new_n529), .B2(new_n530), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n539), .B1(new_n553), .B2(new_n538), .ZN(new_n554));
  OR2_X1    g129(.A1(new_n550), .A2(new_n554), .ZN(G286));
  INV_X1    g130(.A(G286), .ZN(G168));
  NAND2_X1  g131(.A1(new_n509), .A2(G52), .ZN(new_n557));
  INV_X1    g132(.A(G90), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n520), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n522), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(new_n524), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n559), .A2(new_n561), .ZN(G171));
  AOI22_X1  g137(.A1(new_n522), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(new_n524), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n519), .A2(G81), .B1(G43), .B2(new_n509), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT77), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  XOR2_X1   g147(.A(KEYINPUT78), .B(KEYINPUT9), .Z(new_n573));
  NAND3_X1  g148(.A1(new_n509), .A2(new_n573), .A3(G53), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT79), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n509), .A2(G53), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n509), .A2(new_n573), .A3(new_n578), .A4(G53), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n575), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G65), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n516), .B2(new_n518), .ZN(new_n582));
  AND2_X1   g157(.A1(G78), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n519), .A2(G91), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n580), .A2(new_n584), .A3(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  NAND2_X1  g162(.A1(new_n519), .A2(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n509), .A2(G49), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  AND2_X1   g166(.A1(new_n522), .A2(G61), .ZN(new_n592));
  AND2_X1   g167(.A1(G73), .A2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n519), .A2(G86), .B1(G48), .B2(new_n509), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(new_n509), .A2(G47), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n520), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n524), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n519), .A2(G92), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT10), .Z(new_n606));
  AOI22_X1  g181(.A1(new_n522), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n524), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G54), .B2(new_n509), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n604), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(G868), .B2(new_n615), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n475), .A2(new_n472), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT80), .B(G2100), .Z(new_n627));
  OAI22_X1  g202(.A1(new_n625), .A2(KEYINPUT13), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(KEYINPUT13), .B2(new_n625), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n626), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G111), .C2(new_n466), .ZN(new_n633));
  INV_X1    g208(.A(G123), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n489), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n492), .B2(G135), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n631), .A2(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2430), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT83), .ZN(new_n640));
  XOR2_X1   g215(.A(KEYINPUT82), .B(G2438), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT14), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n646), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2443), .B(G2446), .Z(new_n652));
  OR2_X1    g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n660), .B2(KEYINPUT18), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT84), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2100), .ZN(new_n663));
  INV_X1    g238(.A(KEYINPUT18), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n658), .A2(new_n659), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(G2096), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n663), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n671), .A2(new_n676), .A3(new_n674), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n671), .A2(new_n676), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n679));
  AOI211_X1 g254(.A(new_n675), .B(new_n677), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n678), .B2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT86), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(G229));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n689), .A2(G22), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(G303), .B2(G16), .ZN(new_n691));
  INV_X1    g266(.A(G1971), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(G288), .A2(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n689), .A2(G23), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT33), .B(G1976), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT89), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n696), .B(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(KEYINPUT90), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(KEYINPUT90), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n691), .A2(new_n692), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n693), .A2(new_n701), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT91), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n594), .A2(G16), .A3(new_n595), .ZN(new_n707));
  OR2_X1    g282(.A1(G6), .A2(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT32), .B(G1981), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n707), .A2(new_n708), .A3(new_n710), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n712), .A2(KEYINPUT88), .A3(new_n713), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n705), .A2(new_n706), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n718), .ZN(new_n720));
  OAI21_X1  g295(.A(KEYINPUT91), .B1(new_n704), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n719), .A2(KEYINPUT34), .A3(new_n721), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n689), .A2(G24), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n602), .B2(new_n689), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(G1986), .Z(new_n728));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G25), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n492), .A2(G131), .ZN(new_n731));
  INV_X1    g306(.A(G119), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n466), .A2(G107), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n489), .A2(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n730), .B1(new_n736), .B2(new_n729), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT35), .B(G1991), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT87), .Z(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n737), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n728), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n724), .A2(KEYINPUT93), .A3(new_n725), .A4(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT36), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n742), .B1(new_n722), .B2(new_n723), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(new_n725), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G29), .A2(G35), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G162), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT29), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(G2090), .Z(new_n754));
  NOR2_X1   g329(.A1(G16), .A2(G19), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n566), .B2(G16), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT95), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(G1341), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n729), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT97), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT28), .ZN(new_n761));
  INV_X1    g336(.A(G128), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n466), .A2(G116), .ZN(new_n763));
  OAI21_X1  g338(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n764));
  OAI22_X1  g339(.A1(new_n489), .A2(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(new_n492), .B2(G140), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(new_n729), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT96), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n767), .A2(new_n768), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n761), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2067), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n729), .A2(G32), .ZN(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT26), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g352(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n777), .A2(new_n778), .B1(new_n472), .B2(G105), .ZN(new_n779));
  INV_X1    g354(.A(G141), .ZN(new_n780));
  INV_X1    g355(.A(G129), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n779), .B1(new_n469), .B2(new_n780), .C1(new_n781), .C2(new_n489), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(KEYINPUT99), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n774), .B1(new_n786), .B2(new_n729), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT27), .B(G1996), .Z(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n773), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n689), .A2(G20), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT23), .Z(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G299), .B2(G16), .ZN(new_n793));
  INV_X1    g368(.A(G1956), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n689), .A2(G5), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G171), .B2(new_n689), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n797), .A2(G1961), .ZN(new_n798));
  NOR2_X1   g373(.A1(G164), .A2(new_n729), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G27), .B2(new_n729), .ZN(new_n800));
  INV_X1    g375(.A(G2078), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  NOR4_X1   g378(.A1(new_n795), .A2(new_n798), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n754), .A2(new_n758), .A3(new_n790), .A4(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n610), .A2(G16), .ZN(new_n807));
  INV_X1    g382(.A(G4), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G16), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT94), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT94), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n807), .B(new_n811), .C1(new_n808), .C2(G16), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G1348), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n729), .A2(G33), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT25), .Z(new_n818));
  INV_X1    g393(.A(G139), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(new_n469), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g398(.A1(G115), .A2(G2104), .ZN(new_n824));
  INV_X1    g399(.A(G127), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n480), .B2(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n822), .A2(new_n823), .B1(G2105), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n816), .B1(new_n827), .B2(new_n729), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G2072), .ZN(new_n829));
  AOI21_X1  g404(.A(G1348), .B1(new_n810), .B2(new_n812), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n815), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G34), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n832), .A2(KEYINPUT24), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(KEYINPUT24), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n729), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(G160), .B2(new_n729), .ZN(new_n836));
  INV_X1    g411(.A(G2084), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n831), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT102), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n689), .A2(G21), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G168), .B2(new_n689), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(G1966), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(G1966), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n636), .A2(G29), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT31), .B(G11), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT100), .B(G28), .Z(new_n847));
  AND2_X1   g422(.A1(new_n847), .A2(KEYINPUT30), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n729), .B1(new_n847), .B2(KEYINPUT30), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n845), .B(new_n846), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n850), .B1(new_n797), .B2(G1961), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n843), .A2(new_n844), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n806), .A2(new_n839), .A3(new_n840), .A4(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(new_n831), .A3(new_n838), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT102), .B1(new_n856), .B2(new_n805), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n749), .A2(new_n745), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n747), .A2(KEYINPUT93), .A3(new_n725), .A4(new_n859), .ZN(new_n860));
  AND4_X1   g435(.A1(new_n746), .A2(new_n750), .A3(new_n858), .A4(new_n860), .ZN(G311));
  NAND4_X1  g436(.A1(new_n750), .A2(new_n746), .A3(new_n858), .A4(new_n860), .ZN(G150));
  NAND2_X1  g437(.A1(new_n611), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT38), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n865), .A2(new_n524), .ZN(new_n866));
  AOI22_X1  g441(.A1(new_n519), .A2(G93), .B1(G55), .B2(new_n509), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n566), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n564), .A2(new_n565), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n864), .B(new_n873), .Z(new_n874));
  AND2_X1   g449(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n876));
  NOR3_X1   g451(.A1(new_n875), .A2(new_n876), .A3(G860), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n868), .A2(G860), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n879));
  XOR2_X1   g454(.A(new_n878), .B(new_n879), .Z(new_n880));
  OR2_X1    g455(.A1(new_n877), .A2(new_n880), .ZN(G145));
  XNOR2_X1  g456(.A(G160), .B(new_n636), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(G162), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n785), .B(new_n766), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n475), .A2(new_n498), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT104), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n499), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n504), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n884), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n884), .A2(new_n891), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n827), .A2(KEYINPUT105), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n492), .A2(G142), .ZN(new_n896));
  AND4_X1   g471(.A1(G2105), .A2(new_n461), .A3(new_n463), .A4(new_n464), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(G130), .ZN(new_n898));
  OAI21_X1  g473(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT106), .ZN(new_n900));
  INV_X1    g475(.A(G118), .ZN(new_n901));
  AOI22_X1  g476(.A1(new_n899), .A2(new_n900), .B1(new_n901), .B2(G2105), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n900), .B2(new_n899), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n896), .A2(new_n898), .A3(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n625), .B(new_n904), .Z(new_n905));
  NAND2_X1  g480(.A1(new_n895), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n827), .A2(KEYINPUT105), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(new_n736), .ZN(new_n908));
  INV_X1    g483(.A(new_n905), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n892), .A2(new_n893), .A3(new_n894), .A4(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n908), .B1(new_n906), .B2(new_n910), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n883), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n913), .ZN(new_n915));
  INV_X1    g490(.A(new_n883), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(new_n916), .A3(new_n911), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g495(.A(new_n620), .B(new_n873), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n611), .A2(new_n615), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n610), .A2(G299), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n922), .A2(new_n923), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(KEYINPUT41), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT41), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n925), .B1(new_n930), .B2(new_n921), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n931), .A2(KEYINPUT42), .ZN(new_n932));
  XNOR2_X1  g507(.A(G303), .B(new_n602), .ZN(new_n933));
  XOR2_X1   g508(.A(G305), .B(G288), .Z(new_n934));
  XNOR2_X1  g509(.A(new_n933), .B(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(KEYINPUT42), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n932), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n936), .B1(new_n932), .B2(new_n937), .ZN(new_n939));
  OAI21_X1  g514(.A(G868), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(G868), .B2(new_n869), .ZN(G295));
  OAI21_X1  g516(.A(new_n940), .B1(G868), .B2(new_n869), .ZN(G331));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n870), .A2(G301), .A3(new_n872), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(G301), .B1(new_n870), .B2(new_n872), .ZN(new_n946));
  OAI21_X1  g521(.A(G286), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n946), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(G168), .A3(new_n944), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n926), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n927), .A2(new_n947), .A3(new_n929), .A4(new_n949), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(new_n935), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n918), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n935), .B1(new_n951), .B2(new_n952), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n943), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n953), .A2(new_n918), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n955), .A2(KEYINPUT107), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  AOI211_X1 g534(.A(new_n959), .B(new_n935), .C1(new_n951), .C2(new_n952), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n957), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n956), .B1(new_n961), .B2(new_n943), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT44), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT43), .B1(new_n954), .B2(new_n955), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n964), .B1(new_n961), .B2(KEYINPUT43), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n963), .A2(new_n967), .ZN(G397));
  INV_X1    g543(.A(G114), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n500), .B1(new_n969), .B2(G2105), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n897), .B2(G126), .ZN(new_n971));
  AOI221_X4 g546(.A(KEYINPUT104), .B1(new_n475), .B2(new_n498), .C1(new_n497), .C2(KEYINPUT4), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n889), .B1(new_n885), .B2(new_n886), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT45), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n473), .A2(G40), .A3(new_n484), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n766), .B(G2067), .ZN(new_n981));
  INV_X1    g556(.A(G1996), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(new_n786), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n982), .B2(new_n786), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n736), .A2(new_n740), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n731), .A2(new_n739), .A3(new_n735), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n980), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(G290), .A2(G1986), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(KEYINPUT108), .ZN(new_n990));
  NAND2_X1  g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n990), .B(new_n991), .Z(new_n992));
  AOI21_X1  g567(.A(new_n988), .B1(new_n992), .B2(new_n979), .ZN(new_n993));
  INV_X1    g568(.A(G1976), .ZN(new_n994));
  NOR2_X1   g569(.A1(G288), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g570(.A(KEYINPUT111), .B(G8), .Z(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n974), .A2(new_n975), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(new_n978), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT112), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(new_n997), .C1(new_n998), .C2(new_n978), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n995), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT52), .B1(G288), .B2(new_n994), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1003), .A2(KEYINPUT114), .A3(new_n1004), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n1003), .B2(KEYINPUT113), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(KEYINPUT113), .B2(new_n1003), .ZN(new_n1012));
  NOR2_X1   g587(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G305), .A2(G1981), .ZN(new_n1015));
  INV_X1    g590(.A(G1981), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n594), .A2(new_n1016), .A3(new_n595), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  AND2_X1   g593(.A1(KEYINPUT115), .A2(KEYINPUT49), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1014), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1020), .B(new_n1021), .C1(new_n1018), .C2(new_n1014), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1009), .A2(new_n1012), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1025), .A2(G1384), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n974), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1384), .B1(new_n971), .B2(new_n887), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT109), .B1(new_n1028), .B2(KEYINPUT45), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n975), .B1(new_n499), .B2(new_n504), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1032), .A3(new_n1025), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1033), .A2(G40), .A3(new_n473), .A4(new_n484), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT110), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1031), .A2(new_n1032), .A3(new_n1025), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(new_n978), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1031), .A2(new_n1025), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n974), .A2(new_n1026), .B1(new_n1038), .B2(KEYINPUT109), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT110), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1035), .A2(new_n1041), .A3(new_n692), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1031), .A2(KEYINPUT50), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1044), .A2(new_n978), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n974), .A2(new_n1046), .A3(new_n975), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n1048), .A2(G2090), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1024), .B1(new_n1042), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(G303), .A2(G8), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n1051), .B(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1021), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1017), .ZN(new_n1056));
  NOR2_X1   g631(.A1(G288), .A2(G1976), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n1022), .B2(new_n1057), .ZN(new_n1058));
  OAI22_X1  g633(.A1(new_n1023), .A2(new_n1054), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1046), .B1(new_n974), .B2(new_n975), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1046), .B(new_n975), .C1(new_n499), .C2(new_n504), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1061), .A2(new_n473), .A3(G40), .A4(new_n484), .ZN(new_n1062));
  OR3_X1    g637(.A1(new_n1060), .A2(G2090), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n996), .B1(new_n1042), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1054), .B1(new_n1053), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n995), .ZN(new_n1066));
  AND4_X1   g641(.A1(KEYINPUT114), .A2(new_n1021), .A3(new_n1066), .A4(new_n1004), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT114), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1022), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n473), .A2(G40), .A3(new_n484), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(new_n975), .A3(new_n974), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1001), .B1(new_n1071), .B2(new_n997), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1002), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT113), .B(new_n1066), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT52), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1003), .A2(KEYINPUT113), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT116), .B1(new_n1069), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1009), .A2(new_n1012), .A3(new_n1079), .A4(new_n1022), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1065), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1070), .A2(new_n1027), .A3(new_n1029), .A4(new_n1033), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(KEYINPUT110), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1040), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n801), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1085), .A2(KEYINPUT125), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n1088));
  AOI21_X1  g663(.A(G2078), .B1(new_n1035), .B2(new_n1041), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(KEYINPUT53), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1961), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1026), .B1(new_n499), .B2(new_n504), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n473), .A2(new_n1093), .A3(new_n484), .A4(G40), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n976), .A2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1086), .A2(G2078), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1048), .A2(new_n1092), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1091), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1966), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n976), .B2(new_n1094), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1047), .A2(new_n1070), .A3(new_n837), .A4(new_n1043), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n997), .B1(new_n550), .B2(new_n554), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT123), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1105), .B(new_n997), .C1(new_n550), .C2(new_n554), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1024), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1108), .B(KEYINPUT51), .C1(new_n1107), .C2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1102), .A2(new_n997), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1107), .A2(KEYINPUT51), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1110), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1111), .B1(new_n1110), .B2(new_n1114), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1098), .B(G171), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1059), .B1(new_n1081), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1048), .A2(new_n1092), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n482), .A2(G2105), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1122), .A2(G40), .A3(new_n1096), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n977), .A2(new_n473), .A3(new_n1027), .A4(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT125), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1089), .A2(new_n1088), .A3(KEYINPUT53), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(G171), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1097), .A2(G301), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1131), .B1(new_n1091), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1120), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1135));
  AOI21_X1  g710(.A(G301), .B1(new_n1091), .B2(new_n1097), .ZN(new_n1136));
  AOI211_X1 g711(.A(G171), .B(new_n1125), .C1(new_n1087), .C2(new_n1090), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(G1348), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n998), .A2(G2067), .A3(new_n978), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT120), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1047), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1043), .A2(G40), .A3(new_n473), .A4(new_n484), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n814), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n998), .A2(new_n978), .ZN(new_n1145));
  INV_X1    g720(.A(G2067), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(new_n1147), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1141), .A2(new_n1149), .A3(new_n611), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT121), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1141), .A2(new_n1149), .A3(new_n1152), .A4(new_n611), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT56), .B(G2072), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1037), .A2(new_n1039), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n794), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n580), .A2(new_n584), .A3(new_n585), .A4(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1163), .A2(new_n1164), .A3(KEYINPUT122), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1157), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1151), .A2(new_n1153), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1155), .A2(new_n1165), .A3(new_n1156), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1155), .A2(new_n1165), .A3(KEYINPUT119), .A4(new_n1156), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1170), .A2(new_n1175), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1139), .A2(KEYINPUT120), .A3(new_n1140), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1148), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1177), .A2(new_n1178), .A3(KEYINPUT60), .ZN(new_n1179));
  OAI21_X1  g754(.A(KEYINPUT60), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n611), .ZN(new_n1181));
  OAI211_X1 g756(.A(KEYINPUT60), .B(new_n610), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1179), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(KEYINPUT58), .B(G1341), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1082), .A2(G1996), .B1(new_n1145), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n566), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT59), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1185), .A2(new_n1188), .A3(new_n566), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1169), .A2(KEYINPUT61), .A3(new_n1171), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1165), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1192), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1193));
  OAI211_X1 g768(.A(new_n1190), .B(new_n1191), .C1(new_n1193), .C2(KEYINPUT61), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1176), .B1(new_n1183), .B2(new_n1194), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1081), .A2(new_n1134), .A3(new_n1138), .A4(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1119), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1112), .A2(G286), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1054), .A2(KEYINPUT63), .A3(new_n1199), .ZN(new_n1200));
  NOR3_X1   g775(.A1(new_n1023), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1065), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1202), .A2(new_n1203), .A3(new_n1199), .ZN(new_n1204));
  XOR2_X1   g779(.A(KEYINPUT117), .B(KEYINPUT63), .Z(new_n1205));
  AOI21_X1  g780(.A(new_n1201), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n993), .B1(new_n1197), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n979), .A2(new_n982), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT46), .ZN(new_n1209));
  AND2_X1   g784(.A1(new_n786), .A2(new_n981), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1209), .B1(new_n980), .B2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(new_n1211), .B(KEYINPUT126), .ZN(new_n1212));
  OR2_X1    g787(.A1(new_n1212), .A2(KEYINPUT47), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1212), .A2(KEYINPUT47), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n984), .A2(new_n986), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n766), .A2(new_n1146), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n980), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n979), .A2(new_n989), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1218), .B(KEYINPUT127), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT48), .ZN(new_n1220));
  OR2_X1    g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n988), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1217), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AND3_X1   g798(.A1(new_n1213), .A2(new_n1214), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g799(.A1(new_n1207), .A2(new_n1224), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g800(.A(G319), .ZN(new_n1227));
  NOR4_X1   g801(.A1(G229), .A2(new_n1227), .A3(G401), .A4(G227), .ZN(new_n1228));
  NAND3_X1  g802(.A1(new_n965), .A2(new_n1228), .A3(new_n919), .ZN(G225));
  INV_X1    g803(.A(G225), .ZN(G308));
endmodule


