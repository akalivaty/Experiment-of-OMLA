//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n528,
    new_n529, new_n530, new_n531, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n542, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(new_n453), .B(KEYINPUT68), .Z(G261));
  INV_X1    g030(.A(new_n451), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n456), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT69), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n463), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n465), .A2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(new_n468), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n462), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NOR3_X1   g053(.A1(new_n471), .A2(new_n475), .A3(new_n478), .ZN(G160));
  NAND4_X1  g054(.A1(new_n463), .A2(new_n466), .A3(G2105), .A4(new_n468), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n467), .A2(G112), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  OAI22_X1  g058(.A1(new_n480), .A2(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n469), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(G136), .ZN(G162));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n463), .A2(new_n466), .A3(new_n468), .A4(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n472), .A2(new_n468), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n487), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n489), .A2(KEYINPUT4), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G114), .C2(new_n467), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n480), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n492), .A2(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n498), .A2(KEYINPUT6), .A3(G651), .ZN(new_n499));
  AOI21_X1  g074(.A(KEYINPUT6), .B1(new_n498), .B2(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G543), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G88), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n499), .A2(new_n500), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n505), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n509), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT72), .ZN(new_n516));
  XOR2_X1   g091(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n516), .A2(new_n517), .ZN(new_n519));
  INV_X1    g094(.A(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n501), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(G51), .B2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n507), .A2(G89), .ZN(new_n523));
  AND2_X1   g098(.A1(G63), .A2(G651), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n502), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  AOI22_X1  g102(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n511), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n529), .B1(G90), .B2(new_n504), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n521), .A2(G52), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  AOI22_X1  g108(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n511), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n521), .A2(G43), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n504), .A2(G81), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  NAND4_X1  g115(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND4_X1  g118(.A1(G319), .A2(G483), .A3(G661), .A4(new_n543), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT73), .ZN(G188));
  INV_X1    g120(.A(G53), .ZN(new_n546));
  OAI21_X1  g121(.A(KEYINPUT9), .B1(new_n508), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT9), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n521), .A2(new_n548), .A3(G53), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g125(.A(KEYINPUT75), .B(G65), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n502), .A2(KEYINPUT74), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n502), .A2(KEYINPUT74), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g129(.A1(G78), .A2(G543), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n504), .A2(G91), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n550), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(KEYINPUT76), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n550), .A2(new_n560), .A3(new_n556), .A4(new_n557), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G299));
  NAND2_X1  g138(.A1(new_n521), .A2(G49), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n504), .A2(G87), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n568), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G288));
  AOI21_X1  g147(.A(KEYINPUT78), .B1(new_n504), .B2(G86), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n504), .A2(KEYINPUT78), .A3(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n503), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(G651), .A2(new_n579), .B1(new_n521), .B2(G48), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n511), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT79), .ZN(new_n584));
  AOI22_X1  g159(.A1(G47), .A2(new_n521), .B1(new_n504), .B2(G85), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT80), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n585), .A2(KEYINPUT80), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n504), .A2(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT10), .Z(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n552), .B2(new_n553), .ZN(new_n595));
  AND2_X1   g170(.A1(G79), .A2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(G651), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n521), .A2(G54), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n591), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n591), .B1(new_n599), .B2(G868), .ZN(G321));
  XNOR2_X1  g176(.A(new_n562), .B(KEYINPUT81), .ZN(new_n602));
  MUX2_X1   g177(.A(new_n602), .B(G286), .S(G868), .Z(G297));
  XNOR2_X1  g178(.A(G297), .B(KEYINPUT82), .ZN(G280));
  XOR2_X1   g179(.A(KEYINPUT83), .B(G559), .Z(new_n605));
  OAI21_X1  g180(.A(new_n599), .B1(G860), .B2(new_n605), .ZN(G148));
  NAND2_X1  g181(.A1(new_n599), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n539), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n490), .A2(new_n476), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT84), .B(KEYINPUT12), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  INV_X1    g189(.A(G2100), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n485), .A2(G135), .ZN(new_n617));
  INV_X1    g192(.A(G123), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n467), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI22_X1  g195(.A1(new_n480), .A2(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(G2096), .B1(new_n617), .B2(new_n621), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n616), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT85), .Z(G156));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT88), .B(G2438), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n628), .B(new_n629), .Z(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2430), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(KEYINPUT14), .A3(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G1341), .B(G1348), .Z(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n634), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT86), .B(KEYINPUT16), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT87), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n642), .ZN(new_n644));
  AND3_X1   g219(.A1(new_n643), .A2(G14), .A3(new_n644), .ZN(G401));
  INV_X1    g220(.A(KEYINPUT18), .ZN(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT17), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(new_n615), .ZN(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  AOI21_X1  g229(.A(new_n654), .B1(new_n649), .B2(KEYINPUT18), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(new_n623), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n653), .B(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT20), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  OR3_X1    g241(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT89), .ZN(new_n669));
  XOR2_X1   g244(.A(G1981), .B(G1986), .Z(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n669), .B(new_n674), .ZN(G229));
  NOR2_X1   g250(.A1(G4), .A2(G16), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n599), .B2(G16), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT93), .B(G1348), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n677), .B(new_n678), .Z(new_n679));
  NOR2_X1   g254(.A1(G29), .A2(G35), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(G162), .B2(G29), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT29), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G2090), .ZN(new_n683));
  NAND3_X1  g258(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT26), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  AOI22_X1  g262(.A1(new_n686), .A2(new_n687), .B1(G105), .B2(new_n476), .ZN(new_n688));
  INV_X1    g263(.A(G129), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n480), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n485), .B2(G141), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G29), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT95), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n692), .B(new_n693), .C1(G29), .C2(G32), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(new_n693), .B2(new_n692), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT27), .B(G1996), .Z(new_n696));
  AND2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n698));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G26), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G128), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n467), .A2(G116), .ZN(new_n703));
  OAI21_X1  g278(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n704));
  OAI22_X1  g279(.A1(new_n480), .A2(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n485), .B2(G140), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n701), .B1(new_n706), .B2(new_n699), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G2067), .ZN(new_n708));
  NOR4_X1   g283(.A1(new_n679), .A2(new_n683), .A3(new_n697), .A4(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NOR2_X1   g285(.A1(G171), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G5), .B2(new_n710), .ZN(new_n712));
  INV_X1    g287(.A(G1961), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G1341), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n539), .A2(G16), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G16), .B2(G19), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n714), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(G160), .A2(G29), .ZN(new_n719));
  INV_X1    g294(.A(G34), .ZN(new_n720));
  AOI21_X1  g295(.A(G29), .B1(new_n720), .B2(KEYINPUT24), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(KEYINPUT24), .B2(new_n720), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n717), .A2(new_n715), .B1(G2084), .B2(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n699), .A2(G33), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT25), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n490), .A2(G127), .ZN(new_n728));
  INV_X1    g303(.A(G115), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n462), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n727), .B1(new_n730), .B2(G2105), .ZN(new_n731));
  INV_X1    g306(.A(G139), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(new_n469), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n725), .B1(new_n733), .B2(G29), .ZN(new_n734));
  INV_X1    g309(.A(G2072), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n724), .B(new_n736), .C1(new_n695), .C2(new_n696), .ZN(new_n737));
  OAI22_X1  g312(.A1(new_n712), .A2(new_n713), .B1(new_n735), .B2(new_n734), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT30), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT96), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n740), .A2(new_n739), .A3(G28), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n740), .B1(new_n739), .B2(G28), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n699), .B1(new_n739), .B2(G28), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT31), .B(G11), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n622), .B2(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n710), .A2(G21), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G168), .B2(new_n710), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n746), .B1(G2084), .B2(new_n723), .C1(new_n748), .C2(G1966), .ZN(new_n749));
  NOR4_X1   g324(.A1(new_n718), .A2(new_n737), .A3(new_n738), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n710), .A2(G20), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT23), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n562), .B2(new_n710), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT97), .B(G1956), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n748), .A2(G1966), .ZN(new_n756));
  NOR2_X1   g331(.A1(G27), .A2(G29), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G164), .B2(G29), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n756), .B1(G2078), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G2078), .B2(new_n758), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n709), .A2(new_n750), .A3(new_n755), .A4(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n589), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G16), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G16), .B2(G24), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G1986), .ZN(new_n766));
  INV_X1    g341(.A(G1986), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n764), .B(new_n767), .C1(G16), .C2(G24), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(KEYINPUT91), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n699), .A2(G25), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n485), .A2(G131), .ZN(new_n772));
  INV_X1    g347(.A(G119), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n467), .A2(G107), .ZN(new_n774));
  OAI21_X1  g349(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n480), .A2(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n771), .B1(new_n777), .B2(new_n699), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT35), .B(G1991), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n710), .A2(G22), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G166), .B2(new_n710), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(G1971), .Z(new_n783));
  MUX2_X1   g358(.A(G6), .B(G305), .S(G16), .Z(new_n784));
  XOR2_X1   g359(.A(KEYINPUT32), .B(G1981), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  MUX2_X1   g361(.A(G23), .B(new_n567), .S(G16), .Z(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT33), .B(G1976), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n783), .A2(new_n786), .A3(new_n789), .ZN(new_n790));
  AOI211_X1 g365(.A(KEYINPUT92), .B(new_n780), .C1(new_n790), .C2(KEYINPUT34), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT91), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n766), .A2(new_n792), .A3(new_n768), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n790), .A2(KEYINPUT34), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n770), .A2(new_n791), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n761), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n791), .A2(new_n794), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n798), .A2(KEYINPUT36), .A3(new_n793), .A4(new_n770), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT98), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n797), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n800), .B1(new_n797), .B2(new_n799), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(G311));
  NAND2_X1  g378(.A1(new_n797), .A2(new_n799), .ZN(G150));
  NAND2_X1  g379(.A1(new_n599), .A2(G559), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT38), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n521), .A2(G55), .ZN(new_n807));
  NAND2_X1  g382(.A1(G80), .A2(G543), .ZN(new_n808));
  INV_X1    g383(.A(G67), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n503), .B2(new_n809), .ZN(new_n810));
  AOI22_X1  g385(.A1(G651), .A2(new_n810), .B1(new_n504), .B2(G93), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n539), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n807), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(new_n538), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n806), .B(new_n815), .Z(new_n816));
  AND2_X1   g391(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n816), .A2(KEYINPUT39), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n817), .A2(new_n818), .A3(G860), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n813), .A2(G860), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT37), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n819), .A2(new_n821), .ZN(G145));
  XOR2_X1   g397(.A(new_n622), .B(G160), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G162), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n492), .A2(new_n496), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n706), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n691), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n827), .A2(new_n733), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT100), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n777), .B(new_n613), .ZN(new_n830));
  INV_X1    g405(.A(G130), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n467), .A2(G118), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n833));
  OAI22_X1  g408(.A1(new_n480), .A2(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(new_n485), .B2(G142), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n830), .B(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n827), .A2(new_n733), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT99), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n829), .A2(new_n836), .A3(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n836), .B1(new_n829), .B2(new_n838), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n824), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G37), .ZN(new_n843));
  INV_X1    g418(.A(new_n824), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n839), .B(new_n844), .C1(new_n841), .C2(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n841), .A2(new_n845), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n842), .B(new_n843), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g424(.A1(new_n813), .A2(G868), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n599), .A2(new_n561), .A3(new_n559), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n562), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n853), .A3(KEYINPUT102), .ZN(new_n854));
  OR3_X1    g429(.A1(new_n562), .A2(KEYINPUT102), .A3(new_n852), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n851), .A2(new_n853), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n857), .A2(KEYINPUT41), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n854), .A2(KEYINPUT41), .A3(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n607), .B(new_n815), .Z(new_n861));
  MUX2_X1   g436(.A(new_n856), .B(new_n860), .S(new_n861), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT104), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n567), .B(KEYINPUT103), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(new_n589), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n588), .B2(new_n587), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G305), .B(G303), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n866), .A3(new_n867), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT42), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n863), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n862), .A2(KEYINPUT104), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n850), .B1(new_n877), .B2(G868), .ZN(G295));
  AOI21_X1  g453(.A(new_n850), .B1(new_n877), .B2(G868), .ZN(G331));
  NAND3_X1  g454(.A1(new_n812), .A2(new_n814), .A3(G301), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(G301), .B1(new_n812), .B2(new_n814), .ZN(new_n882));
  OAI21_X1  g457(.A(G286), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n882), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n884), .A2(G168), .A3(new_n880), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n885), .A3(KEYINPUT41), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n856), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n857), .A2(new_n883), .A3(new_n885), .A4(KEYINPUT41), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n873), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT105), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n887), .A2(new_n891), .A3(new_n873), .A4(new_n888), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n894));
  INV_X1    g469(.A(new_n873), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n883), .A2(new_n885), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(new_n858), .B2(new_n859), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n856), .A2(new_n896), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n895), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n893), .A2(new_n894), .A3(new_n843), .A4(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n843), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n897), .A2(new_n899), .A3(new_n895), .ZN(new_n904));
  OAI21_X1  g479(.A(KEYINPUT43), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n900), .A2(new_n890), .A3(new_n843), .A4(new_n892), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n911));
  OR3_X1    g486(.A1(new_n903), .A2(KEYINPUT43), .A3(new_n904), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n906), .B1(new_n913), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g489(.A(G1384), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(new_n492), .B2(new_n496), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n466), .A2(new_n468), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n919), .A2(G137), .A3(new_n467), .A4(new_n463), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n473), .A2(new_n474), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(G2105), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n920), .A2(new_n922), .A3(G40), .A4(new_n477), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G1996), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n925), .A3(new_n691), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n926), .B(KEYINPUT107), .Z(new_n927));
  XNOR2_X1  g502(.A(new_n706), .B(G2067), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n925), .B2(new_n691), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n924), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g506(.A(new_n777), .B(new_n779), .Z(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n924), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n589), .B(new_n767), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n934), .B1(new_n924), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n916), .A2(new_n923), .ZN(new_n937));
  INV_X1    g512(.A(G8), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G1981), .ZN(new_n940));
  INV_X1    g515(.A(new_n575), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n940), .B(new_n580), .C1(new_n941), .C2(new_n573), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT113), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT113), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n576), .A2(new_n944), .A3(new_n940), .A4(new_n580), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(KEYINPUT114), .B(G86), .Z(new_n947));
  NAND2_X1  g522(.A1(new_n504), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n940), .B1(new_n580), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n946), .A2(KEYINPUT49), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT49), .B1(new_n946), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n953), .A2(G1976), .A3(G288), .ZN(new_n954));
  INV_X1    g529(.A(new_n946), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n939), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n923), .ZN(new_n957));
  OAI211_X1 g532(.A(KEYINPUT45), .B(new_n915), .C1(new_n492), .C2(new_n496), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n918), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n923), .B1(new_n916), .B2(new_n917), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(KEYINPUT108), .A3(new_n958), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT109), .B(G1971), .Z(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n916), .A2(KEYINPUT50), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n968), .B1(new_n492), .B2(new_n496), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n957), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(KEYINPUT110), .B(G2090), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n965), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(G303), .A2(G8), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT55), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n965), .A2(new_n973), .A3(KEYINPUT111), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n976), .A2(new_n979), .A3(G8), .A4(new_n980), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n564), .A2(new_n565), .A3(G1976), .A4(new_n566), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT112), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n939), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT52), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n986), .B1(new_n571), .B2(G1976), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n953), .B2(new_n939), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n956), .B1(new_n981), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT63), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n971), .A2(KEYINPUT115), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n972), .B1(new_n971), .B2(KEYINPUT115), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n965), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G8), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n978), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n989), .A2(new_n997), .A3(new_n981), .ZN(new_n998));
  INV_X1    g573(.A(G2084), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n966), .A2(new_n999), .A3(new_n957), .A4(new_n969), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT116), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1966), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n959), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n923), .B1(new_n825), .B2(new_n968), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1005), .A2(KEYINPUT116), .A3(new_n999), .A4(new_n966), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1007), .A2(G8), .A3(G168), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n992), .B1(new_n998), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n976), .A2(G8), .A3(new_n980), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(new_n978), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1009), .A2(new_n992), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1012), .A2(new_n1013), .A3(new_n981), .A4(new_n989), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n991), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G2078), .B1(new_n961), .B2(new_n963), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT124), .B1(new_n1016), .B2(KEYINPUT53), .ZN(new_n1017));
  INV_X1    g592(.A(G2078), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n962), .A2(KEYINPUT108), .A3(new_n958), .ZN(new_n1019));
  AOI21_X1  g594(.A(KEYINPUT108), .B1(new_n962), .B2(new_n958), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT124), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1017), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n967), .B2(new_n970), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1005), .A2(KEYINPUT117), .A3(new_n966), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(new_n713), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n962), .A2(KEYINPUT53), .A3(new_n1018), .A4(new_n958), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G171), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1025), .A2(G301), .A3(new_n1032), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n998), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1007), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1002), .A2(new_n1004), .A3(new_n1006), .A4(KEYINPUT121), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G168), .ZN(new_n1043));
  AND2_X1   g618(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT122), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n1007), .B2(G8), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1007), .A2(new_n1046), .A3(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G168), .A2(new_n938), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(KEYINPUT51), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1048), .A2(KEYINPUT123), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n1047), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1045), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1040), .A2(new_n1050), .A3(new_n1041), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT125), .ZN(new_n1059));
  AOI21_X1  g634(.A(G301), .B1(new_n1025), .B2(new_n1032), .ZN(new_n1060));
  AOI211_X1 g635(.A(G171), .B(new_n1031), .C1(new_n1017), .C2(new_n1024), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1059), .B1(new_n1062), .B2(KEYINPUT54), .ZN(new_n1063));
  NOR4_X1   g638(.A1(new_n1060), .A2(new_n1061), .A3(KEYINPUT125), .A4(new_n1037), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1038), .B(new_n1058), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT61), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n558), .A2(KEYINPUT57), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n558), .A2(KEYINPUT57), .ZN(new_n1068));
  INV_X1    g643(.A(G1956), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n967), .B2(new_n970), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT56), .B(G2072), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n962), .A2(new_n958), .A3(new_n1071), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1067), .A2(new_n1068), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1066), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT58), .B(G1341), .ZN(new_n1077));
  OAI22_X1  g652(.A1(new_n959), .A2(G1996), .B1(new_n937), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n538), .B1(new_n1079), .B2(KEYINPUT59), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1079), .A2(KEYINPUT59), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1081), .B(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1075), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(KEYINPUT61), .A3(new_n1073), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1076), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1348), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1027), .A2(new_n1028), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G2067), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n937), .A2(new_n1089), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(KEYINPUT119), .A3(KEYINPUT60), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(KEYINPUT60), .A3(new_n1090), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1093), .A2(new_n1094), .A3(new_n852), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n852), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1092), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1091), .A2(KEYINPUT60), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1086), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1091), .A2(new_n852), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1073), .B1(new_n1101), .B2(new_n1075), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT120), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n599), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1093), .A2(new_n1094), .A3(new_n852), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1098), .B1(new_n1109), .B2(new_n1092), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1105), .B(new_n1102), .C1(new_n1110), .C2(new_n1086), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1104), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1015), .B1(new_n1065), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1056), .A2(new_n1114), .A3(new_n1057), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n998), .A2(new_n1034), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(KEYINPUT126), .A3(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1058), .A2(KEYINPUT62), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT126), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n936), .B1(new_n1113), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n924), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n691), .B2(new_n928), .ZN(new_n1124));
  XOR2_X1   g699(.A(new_n1124), .B(KEYINPUT127), .Z(new_n1125));
  NAND2_X1  g700(.A1(new_n924), .A2(new_n925), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT46), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(new_n1128), .B(KEYINPUT47), .Z(new_n1129));
  OR4_X1    g704(.A1(new_n779), .A2(new_n931), .A3(new_n772), .A4(new_n776), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n706), .A2(new_n1089), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1123), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n589), .A2(new_n767), .A3(new_n924), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT48), .ZN(new_n1134));
  AOI211_X1 g709(.A(new_n1129), .B(new_n1132), .C1(new_n933), .C2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1122), .A2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g711(.A1(new_n901), .A2(new_n905), .ZN(new_n1138));
  NOR4_X1   g712(.A1(G229), .A2(G401), .A3(new_n460), .A4(G227), .ZN(new_n1139));
  NAND3_X1  g713(.A1(new_n848), .A2(new_n1138), .A3(new_n1139), .ZN(G225));
  INV_X1    g714(.A(G225), .ZN(G308));
endmodule


