//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n554, new_n555, new_n556, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT68), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n460), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT69), .ZN(G160));
  AOI21_X1  g054(.A(new_n460), .B1(new_n466), .B2(new_n468), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT70), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OAI21_X1  g057(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G112), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n475), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G136), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n490), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n463), .A2(new_n469), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT71), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n495), .A2(new_n498), .A3(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n463), .A2(new_n469), .A3(KEYINPUT72), .A4(new_n491), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n494), .A2(new_n497), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G2105), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n480), .B2(G126), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  AND2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g088(.A(new_n513), .B(KEYINPUT74), .Z(new_n514));
  NOR2_X1   g089(.A1(new_n508), .A2(new_n509), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OR3_X1    g093(.A1(new_n515), .A2(new_n518), .A3(KEYINPUT73), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT73), .B1(new_n515), .B2(new_n518), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n521), .A2(G88), .B1(G50), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n514), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XOR2_X1   g101(.A(new_n526), .B(KEYINPUT7), .Z(new_n527));
  AND3_X1   g102(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n528));
  AOI211_X1 g103(.A(new_n527), .B(new_n528), .C1(G51), .C2(new_n523), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n521), .A2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n515), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G651), .B1(new_n523), .B2(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n519), .A2(new_n520), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  NAND2_X1  g115(.A1(new_n521), .A2(G81), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n515), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n512), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n546), .B1(new_n545), .B2(new_n544), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n523), .A2(G43), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n541), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n521), .A2(new_n558), .A3(G91), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT77), .B1(new_n537), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n523), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OR3_X1    g139(.A1(new_n563), .A2(KEYINPUT9), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT9), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n515), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n565), .A2(new_n566), .B1(G651), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n562), .A2(new_n570), .ZN(G299));
  NAND2_X1  g146(.A1(new_n514), .A2(new_n524), .ZN(G303));
  NAND2_X1  g147(.A1(new_n521), .A2(G87), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n510), .A2(G74), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(G49), .B2(new_n523), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(G288));
  NAND3_X1  g151(.A1(new_n519), .A2(G86), .A3(new_n520), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n515), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n523), .B2(G48), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT78), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n577), .A2(new_n584), .A3(new_n581), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(new_n523), .A2(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI221_X1 g165(.A(new_n588), .B1(new_n512), .B2(new_n589), .C1(new_n537), .C2(new_n590), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(KEYINPUT79), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(KEYINPUT79), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT80), .Z(new_n596));
  INV_X1    g171(.A(G92), .ZN(new_n597));
  XNOR2_X1  g172(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n598));
  OR3_X1    g173(.A1(new_n537), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n537), .B2(new_n597), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n515), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(new_n523), .B2(G54), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n599), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n596), .B1(G868), .B2(new_n606), .ZN(G321));
  XNOR2_X1  g182(.A(G321), .B(KEYINPUT82), .ZN(G284));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n562), .A2(new_n570), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g193(.A1(new_n463), .A2(new_n469), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n473), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n481), .A2(G123), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n486), .A2(G135), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n460), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2096), .Z(new_n631));
  NAND3_X1  g206(.A1(new_n624), .A2(new_n625), .A3(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT83), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2427), .B(G2430), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n635), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT16), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n642), .B(new_n643), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n640), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(G14), .B1(new_n645), .B2(new_n647), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(G401));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT84), .ZN(new_n652));
  NOR2_X1   g227(.A1(G2072), .A2(G2078), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n442), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n654), .B(KEYINPUT17), .Z(new_n659));
  OAI211_X1 g234(.A(new_n656), .B(new_n658), .C1(new_n659), .C2(new_n652), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n654), .A2(new_n657), .A3(new_n651), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n652), .A3(new_n657), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n623), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT85), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT19), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT86), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  OR3_X1    g255(.A1(new_n673), .A2(new_n680), .A3(new_n676), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n673), .A2(new_n680), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT20), .Z(new_n684));
  OAI21_X1  g259(.A(new_n670), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n682), .A2(new_n684), .A3(new_n670), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n669), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n687), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n689), .A2(new_n685), .A3(new_n668), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n688), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  AND3_X1   g271(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n693), .B2(new_n695), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(G229));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G32), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n481), .A2(G129), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT92), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n486), .A2(G141), .ZN(new_n705));
  NAND3_X1  g280(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT26), .Z(new_n707));
  NAND4_X1  g282(.A1(new_n702), .A2(new_n704), .A3(new_n705), .A4(new_n707), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n708), .A2(KEYINPUT93), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(KEYINPUT93), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n701), .B1(new_n712), .B2(new_n700), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT27), .B(G1996), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n700), .A2(G35), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G162), .B2(new_n700), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT29), .ZN(new_n717));
  OAI22_X1  g292(.A1(new_n713), .A2(new_n714), .B1(G2090), .B2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NOR2_X1   g294(.A1(G168), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n719), .B2(G21), .ZN(new_n721));
  INV_X1    g296(.A(G1966), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n606), .A2(G16), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G4), .B2(G16), .ZN(new_n725));
  INV_X1    g300(.A(G1348), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n721), .A2(new_n722), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n700), .A2(G26), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n481), .A2(G128), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n732));
  INV_X1    g307(.A(G116), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G2105), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n486), .B2(G140), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n730), .B1(new_n737), .B2(new_n700), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT91), .B(G2067), .Z(new_n739));
  NOR2_X1   g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR4_X1   g315(.A1(new_n723), .A2(new_n727), .A3(new_n728), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n719), .A2(G5), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G171), .B2(new_n719), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT94), .Z(new_n744));
  AOI22_X1  g319(.A1(new_n744), .A2(G1961), .B1(new_n725), .B2(new_n726), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n718), .B(new_n746), .C1(G2090), .C2(new_n717), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n713), .A2(new_n714), .ZN(new_n748));
  NAND2_X1  g323(.A1(G160), .A2(G29), .ZN(new_n749));
  INV_X1    g324(.A(G34), .ZN(new_n750));
  AOI21_X1  g325(.A(G29), .B1(new_n750), .B2(KEYINPUT24), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(KEYINPUT24), .B2(new_n750), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  OAI221_X1 g328(.A(new_n748), .B1(G1961), .B2(new_n744), .C1(G2084), .C2(new_n753), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT95), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n719), .A2(G20), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT23), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n610), .B2(new_n719), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1956), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT31), .B(G11), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n630), .A2(new_n700), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT30), .B(G28), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n760), .B(new_n761), .C1(new_n700), .C2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n700), .A2(G33), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n619), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(new_n460), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT25), .Z(new_n768));
  INV_X1    g343(.A(G139), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n475), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(new_n700), .ZN(new_n772));
  INV_X1    g347(.A(new_n739), .ZN(new_n773));
  INV_X1    g348(.A(new_n738), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n763), .B1(G2072), .B2(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G2072), .B2(new_n772), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n700), .A2(G27), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G164), .B2(new_n700), .ZN(new_n778));
  INV_X1    g353(.A(G2078), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  AOI211_X1 g356(.A(new_n759), .B(new_n781), .C1(G2084), .C2(new_n753), .ZN(new_n782));
  NOR2_X1   g357(.A1(G16), .A2(G19), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(new_n550), .B2(G16), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT90), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1341), .Z(new_n786));
  NAND4_X1  g361(.A1(new_n747), .A2(new_n755), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT36), .ZN(new_n788));
  OR2_X1    g363(.A1(G16), .A2(G24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G290), .B2(new_n719), .ZN(new_n790));
  INV_X1    g365(.A(G1986), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n700), .A2(G25), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n481), .A2(G119), .ZN(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n796));
  INV_X1    g371(.A(G107), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(G2105), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n486), .B2(G131), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n794), .B1(new_n801), .B2(new_n700), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT35), .B(G1991), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n792), .A2(new_n793), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n719), .A2(G22), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G166), .B2(new_n719), .ZN(new_n807));
  INV_X1    g382(.A(G1971), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n719), .A2(G23), .ZN(new_n810));
  INV_X1    g385(.A(G288), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n719), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT33), .B(G1976), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT88), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n812), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n809), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g391(.A1(G6), .A2(G16), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n586), .B2(G16), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT32), .B(G1981), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT34), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n805), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(KEYINPUT89), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(KEYINPUT89), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n821), .A2(new_n822), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n788), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n826), .A2(new_n788), .A3(new_n828), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n787), .B1(new_n830), .B2(new_n831), .ZN(G311));
  INV_X1    g407(.A(new_n787), .ZN(new_n833));
  INV_X1    g408(.A(new_n831), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n829), .ZN(G150));
  AOI22_X1  g410(.A1(new_n521), .A2(G93), .B1(G55), .B2(new_n523), .ZN(new_n836));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  INV_X1    g412(.A(G67), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n515), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n512), .B1(new_n839), .B2(KEYINPUT97), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(KEYINPUT97), .B2(new_n839), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n613), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT98), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n550), .A2(new_n841), .A3(new_n836), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n842), .A2(new_n549), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n848), .B(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT99), .Z(new_n854));
  AOI21_X1  g429(.A(G860), .B1(new_n852), .B2(KEYINPUT39), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n854), .A2(KEYINPUT100), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT100), .B1(new_n854), .B2(new_n855), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n844), .B1(new_n856), .B2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(G160), .B(new_n630), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n488), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n711), .A2(new_n736), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n709), .A2(new_n710), .A3(new_n737), .ZN(new_n863));
  AND3_X1   g438(.A1(new_n862), .A2(new_n506), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n506), .B1(new_n862), .B2(new_n863), .ZN(new_n865));
  OAI22_X1  g440(.A1(new_n864), .A2(new_n865), .B1(new_n766), .B2(new_n770), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(G164), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n862), .A2(new_n506), .A3(new_n863), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n868), .A2(new_n771), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n486), .A2(G142), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n460), .A2(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(G130), .B2(new_n481), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n621), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n801), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n871), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n866), .A2(new_n870), .A3(new_n878), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(KEYINPUT101), .B2(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n881), .A2(KEYINPUT101), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n861), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n881), .A2(new_n860), .ZN(new_n885));
  AOI21_X1  g460(.A(G37), .B1(new_n885), .B2(new_n880), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(G395));
  INV_X1    g464(.A(G868), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n842), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n610), .A2(new_n606), .ZN(new_n892));
  NAND2_X1  g467(.A1(G299), .A2(new_n605), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT41), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n892), .A2(new_n896), .A3(new_n893), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(KEYINPUT103), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(new_n899), .A3(KEYINPUT41), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n851), .B(new_n615), .ZN(new_n902));
  MUX2_X1   g477(.A(new_n901), .B(new_n894), .S(new_n902), .Z(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(G166), .A2(G305), .ZN(new_n906));
  NAND2_X1  g481(.A1(G303), .A2(new_n586), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT104), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(G290), .A2(G288), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n592), .A2(new_n811), .A3(new_n593), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n909), .A2(new_n911), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(KEYINPUT104), .A3(new_n908), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n905), .B(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n891), .B1(new_n918), .B2(new_n890), .ZN(G295));
  OAI21_X1  g494(.A(new_n891), .B1(new_n918), .B2(new_n890), .ZN(G331));
  INV_X1    g495(.A(new_n917), .ZN(new_n921));
  XNOR2_X1  g496(.A(G286), .B(G301), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n851), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(G286), .B(G171), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(new_n850), .A3(new_n849), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n923), .A2(new_n925), .A3(new_n893), .A4(new_n892), .ZN(new_n926));
  INV_X1    g501(.A(new_n925), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n851), .A2(KEYINPUT106), .A3(new_n922), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n921), .B(new_n926), .C1(new_n901), .C2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  INV_X1    g508(.A(G37), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n925), .A2(new_n893), .A3(new_n892), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n935), .B1(new_n929), .B2(new_n930), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n895), .A2(new_n897), .B1(new_n923), .B2(new_n925), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n917), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n926), .B1(new_n901), .B2(new_n931), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n917), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n932), .A2(new_n941), .A3(new_n934), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n939), .B1(new_n942), .B2(new_n933), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n932), .A2(new_n941), .A3(new_n933), .A4(new_n934), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n946), .A2(KEYINPUT44), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n938), .B(new_n934), .C1(new_n940), .C2(new_n917), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT107), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n932), .A2(new_n950), .A3(new_n934), .A4(new_n938), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n951), .A3(KEYINPUT43), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n947), .A2(new_n952), .A3(KEYINPUT108), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT108), .B1(new_n947), .B2(new_n952), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n945), .B1(new_n953), .B2(new_n954), .ZN(G397));
  XNOR2_X1  g530(.A(G299), .B(KEYINPUT57), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1956), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n959));
  XNOR2_X1  g534(.A(KEYINPUT109), .B(G40), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n959), .B1(new_n478), .B2(new_n961), .ZN(new_n962));
  NOR4_X1   g537(.A1(new_n472), .A2(new_n477), .A3(KEYINPUT110), .A4(new_n960), .ZN(new_n963));
  AOI21_X1  g538(.A(G1384), .B1(new_n501), .B2(new_n505), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n965));
  OAI22_X1  g540(.A1(new_n962), .A2(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n964), .A2(KEYINPUT116), .A3(new_n965), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT116), .B1(new_n964), .B2(new_n965), .ZN(new_n968));
  OAI22_X1  g543(.A1(new_n966), .A2(KEYINPUT115), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n506), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n470), .A2(new_n471), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(G2105), .ZN(new_n973));
  INV_X1    g548(.A(new_n477), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n974), .A3(new_n961), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT110), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n478), .A2(new_n959), .A3(new_n961), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n971), .A2(KEYINPUT50), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n958), .B1(new_n969), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n971), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n976), .A2(new_n977), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n964), .A2(KEYINPUT45), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  XOR2_X1   g561(.A(KEYINPUT56), .B(G2072), .Z(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n957), .B1(new_n981), .B2(new_n989), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n977), .A2(new_n976), .B1(new_n964), .B2(new_n965), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n971), .A2(new_n992), .A3(KEYINPUT50), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT112), .B1(new_n964), .B2(new_n965), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n991), .A2(new_n993), .A3(KEYINPUT117), .A4(new_n994), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n726), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n984), .A2(new_n964), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G2067), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n605), .B1(new_n999), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n981), .A2(new_n957), .A3(new_n989), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n990), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n506), .A2(new_n965), .A3(new_n970), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n964), .A2(KEYINPUT116), .A3(new_n965), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n978), .A2(new_n979), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n966), .A2(KEYINPUT115), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1956), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n956), .B1(new_n1013), .B2(new_n988), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(KEYINPUT61), .A3(new_n1005), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT118), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1014), .A2(new_n1017), .A3(KEYINPUT61), .A4(new_n1005), .ZN(new_n1018));
  AND2_X1   g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  AND3_X1   g594(.A1(new_n999), .A2(new_n605), .A3(new_n1003), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT60), .B1(new_n1020), .B2(new_n1004), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT61), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1005), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(new_n990), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n605), .A2(KEYINPUT60), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n999), .A2(new_n1003), .A3(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT58), .B(G1341), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1001), .A2(new_n1027), .B1(new_n986), .B2(G1996), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n550), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT59), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1021), .A2(new_n1024), .A3(new_n1026), .A4(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1006), .B1(new_n1019), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n986), .A2(new_n722), .ZN(new_n1033));
  INV_X1    g608(.A(G2084), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n991), .A2(new_n993), .A3(new_n1034), .A4(new_n994), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(G168), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  AOI21_X1  g612(.A(G168), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT51), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1040), .A3(G8), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT119), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT111), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n962), .A2(new_n963), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT45), .B1(new_n506), .B2(new_n970), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n982), .B(G1384), .C1(new_n501), .C2(new_n505), .ZN(new_n1047));
  NOR3_X1   g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1044), .B1(new_n1048), .B2(G1971), .ZN(new_n1049));
  INV_X1    g624(.A(G2090), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n991), .A2(new_n993), .A3(new_n1050), .A4(new_n994), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n986), .A2(KEYINPUT111), .A3(new_n808), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n1056), .B(new_n1057), .C1(G303), .C2(G8), .ZN(new_n1058));
  AND4_X1   g633(.A1(new_n1054), .A2(G303), .A3(new_n1055), .A4(G8), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1053), .A2(G8), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n582), .A2(G1981), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n582), .A2(G1981), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT49), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1062), .B(new_n1067), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1066), .A2(G8), .A3(new_n1000), .A4(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n811), .A2(G1976), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1000), .A2(new_n1070), .A3(G8), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT52), .ZN(new_n1072));
  INV_X1    g647(.A(G1976), .ZN(new_n1073));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(G288), .B2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1000), .A2(new_n1070), .A3(new_n1074), .A4(G8), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1069), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1061), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1011), .A2(new_n1050), .A3(new_n1012), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n986), .A2(new_n808), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1060), .B1(new_n1081), .B2(G8), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1039), .A2(new_n1084), .A3(new_n1041), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1043), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1961), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n997), .A2(new_n1087), .A3(new_n998), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n986), .B2(G2078), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n478), .A2(G40), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT121), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1091), .B(new_n1092), .C1(new_n964), .C2(KEYINPUT45), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1093), .A2(KEYINPUT53), .A3(new_n779), .A4(new_n985), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1092), .B1(new_n983), .B2(new_n1091), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1088), .A2(new_n1090), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(G171), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT54), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1048), .A2(KEYINPUT53), .A3(new_n779), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1088), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1090), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1088), .B2(new_n1101), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1099), .B1(new_n1105), .B2(G301), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1086), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(G171), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(G171), .B2(new_n1097), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1032), .A2(new_n1107), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1043), .A2(KEYINPUT62), .A3(new_n1085), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1043), .A2(new_n1085), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1043), .A2(KEYINPUT122), .A3(KEYINPUT62), .A4(new_n1085), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1083), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(new_n1108), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1115), .A2(new_n1118), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1069), .A2(new_n1073), .A3(new_n811), .ZN(new_n1123));
  OAI211_X1 g698(.A(G8), .B(new_n1000), .C1(new_n1123), .C2(new_n1064), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1061), .B2(new_n1076), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1127), .A2(G8), .A3(G168), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1120), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1060), .B1(new_n1053), .B2(G8), .ZN(new_n1130));
  OR4_X1    g705(.A1(new_n1126), .A2(new_n1078), .A3(new_n1128), .A4(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1125), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1112), .A2(new_n1122), .A3(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n983), .A2(new_n1045), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n736), .B(new_n1002), .ZN(new_n1135));
  INV_X1    g710(.A(G1996), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1135), .B1(new_n712), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1136), .B2(new_n712), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n801), .A2(new_n803), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n801), .A2(new_n803), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g716(.A(G290), .B(G1986), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1134), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1133), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1134), .A2(new_n791), .A3(new_n593), .A4(new_n592), .ZN(new_n1145));
  XOR2_X1   g720(.A(new_n1145), .B(KEYINPUT48), .Z(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1134), .B2(new_n1141), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1148));
  NOR2_X1   g723(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1148), .B(new_n1149), .Z(new_n1150));
  NAND2_X1  g725(.A1(new_n712), .A2(new_n1135), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1151), .A2(new_n1134), .B1(KEYINPUT124), .B2(KEYINPUT46), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1139), .B(KEYINPUT123), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1138), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(G2067), .B2(new_n736), .ZN(new_n1158));
  AOI211_X1 g733(.A(new_n1147), .B(new_n1155), .C1(new_n1134), .C2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1144), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g735(.A(G319), .B1(new_n648), .B2(new_n649), .ZN(new_n1162));
  NOR2_X1   g736(.A1(G227), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g737(.A(new_n1163), .B1(new_n697), .B2(new_n698), .ZN(new_n1164));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g740(.A(KEYINPUT126), .B(new_n1163), .C1(new_n697), .C2(new_n698), .ZN(new_n1167));
  AOI22_X1  g741(.A1(new_n884), .A2(new_n886), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AND3_X1   g742(.A1(new_n943), .A2(new_n1168), .A3(KEYINPUT127), .ZN(new_n1169));
  AOI21_X1  g743(.A(KEYINPUT127), .B1(new_n943), .B2(new_n1168), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n1169), .A2(new_n1170), .ZN(G308));
  NAND2_X1  g745(.A1(new_n943), .A2(new_n1168), .ZN(G225));
endmodule


