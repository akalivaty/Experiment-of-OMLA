//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n770, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981;
  AND2_X1   g000(.A1(G71gat), .A2(G78gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(G57gat), .B(G64gat), .Z(new_n205));
  AOI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(KEYINPUT92), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(KEYINPUT9), .B2(new_n202), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OAI221_X1 g007(.A(new_n205), .B1(KEYINPUT9), .B2(new_n202), .C1(new_n204), .C2(KEYINPUT92), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G231gat), .A2(G233gat), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n213), .B(new_n214), .Z(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(G127gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n217), .A2(G1gat), .ZN(new_n218));
  OAI21_X1  g017(.A(G8gat), .B1(new_n218), .B2(KEYINPUT89), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n217), .B1(new_n220), .B2(G1gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G1gat), .B2(new_n217), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n219), .B(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(KEYINPUT21), .B2(new_n210), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n216), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G127gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n215), .B(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n225), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G183gat), .B(G211gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT94), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n233));
  INV_X1    g032(.A(G155gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n232), .B(new_n235), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n226), .A2(new_n230), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n226), .B2(new_n230), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n240));
  OR3_X1    g039(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n241), .A2(KEYINPUT87), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(KEYINPUT87), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G43gat), .B(G50gat), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n245), .A2(KEYINPUT15), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n245), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT88), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n244), .A2(KEYINPUT88), .A3(new_n246), .A4(new_n247), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n241), .A2(new_n240), .ZN(new_n253));
  NAND2_X1  g052(.A1(G29gat), .A2(G36gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n255), .A2(KEYINPUT15), .A3(new_n245), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT17), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G85gat), .A2(G92gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT7), .ZN(new_n262));
  INV_X1    g061(.A(G99gat), .ZN(new_n263));
  INV_X1    g062(.A(G106gat), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT8), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XOR2_X1   g064(.A(KEYINPUT95), .B(G85gat), .Z(new_n266));
  OAI211_X1 g065(.A(new_n262), .B(new_n265), .C1(G92gat), .C2(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G99gat), .B(G106gat), .Z(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n267), .B(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT96), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n267), .B(new_n268), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT96), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n256), .B1(new_n250), .B2(new_n251), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT17), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  AND3_X1   g078(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n275), .B2(new_n258), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g081(.A(G190gat), .B(G218gat), .Z(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n283), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n279), .A2(new_n285), .A3(new_n281), .ZN(new_n286));
  XOR2_X1   g085(.A(G134gat), .B(G162gat), .Z(new_n287));
  AOI21_X1  g086(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n289), .A2(KEYINPUT97), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n284), .A2(new_n286), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(KEYINPUT97), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n292), .B(KEYINPUT98), .Z(new_n293));
  XNOR2_X1  g092(.A(new_n291), .B(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n239), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n252), .A2(new_n257), .A3(new_n223), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT90), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n277), .A2(KEYINPUT90), .A3(new_n223), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n258), .A2(new_n224), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G229gat), .A2(G233gat), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n302), .B(KEYINPUT13), .Z(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(KEYINPUT91), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT91), .B1(new_n301), .B2(new_n303), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n223), .B1(new_n277), .B2(KEYINPUT17), .ZN(new_n308));
  AOI211_X1 g107(.A(new_n259), .B(new_n256), .C1(new_n250), .C2(new_n251), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n302), .B(new_n300), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT18), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G113gat), .B(G141gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G169gat), .B(G197gat), .Z(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(KEYINPUT86), .B(KEYINPUT12), .Z(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n307), .A2(new_n312), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n301), .A2(new_n303), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT91), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n304), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT18), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n319), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G230gat), .A2(G233gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n272), .A2(new_n210), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n270), .A2(new_n211), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT10), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n210), .A2(KEYINPUT10), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n274), .B2(new_n271), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n330), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n330), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n332), .A2(new_n331), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(G176gat), .B(G204gat), .Z(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT101), .ZN(new_n341));
  XNOR2_X1  g140(.A(G120gat), .B(G148gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n339), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n336), .A2(new_n338), .A3(new_n345), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n295), .A2(new_n329), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G226gat), .ZN(new_n352));
  INV_X1    g151(.A(G233gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(G169gat), .ZN(new_n357));
  INV_X1    g156(.A(G176gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT26), .ZN(new_n359));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT26), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n356), .B(new_n359), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G183gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT27), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT27), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G183gat), .ZN(new_n368));
  INV_X1    g167(.A(G190gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n366), .A2(new_n368), .A3(KEYINPUT28), .A4(new_n369), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n364), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT25), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT24), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n356), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT64), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(new_n365), .A3(new_n369), .ZN(new_n379));
  NAND3_X1  g178(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n381));
  AND4_X1   g180(.A1(new_n377), .A2(new_n379), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n363), .A2(KEYINPUT23), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(G169gat), .B2(G176gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n383), .A2(new_n360), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n375), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n383), .A2(new_n360), .A3(new_n385), .ZN(new_n388));
  NOR2_X1   g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n376), .A2(KEYINPUT65), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n356), .A3(new_n391), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n391), .A2(new_n356), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n388), .A2(KEYINPUT25), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n374), .B1(new_n387), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n355), .B1(new_n395), .B2(KEYINPUT29), .ZN(new_n396));
  NAND2_X1  g195(.A1(G211gat), .A2(G218gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(G211gat), .A2(G218gat), .ZN(new_n399));
  NOR3_X1   g198(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT70), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT22), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(G197gat), .A2(G204gat), .ZN(new_n403));
  AND2_X1   g202(.A1(G197gat), .A2(G204gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  OR2_X1    g205(.A1(G197gat), .A2(G204gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(G197gat), .A2(G204gat), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n407), .A2(new_n408), .B1(new_n401), .B2(new_n397), .ZN(new_n409));
  INV_X1    g208(.A(G211gat), .ZN(new_n410));
  INV_X1    g209(.A(G218gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT70), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n413), .A3(new_n397), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n406), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n372), .A2(new_n373), .ZN(new_n417));
  INV_X1    g216(.A(new_n364), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n379), .A2(new_n377), .A3(new_n380), .A4(new_n381), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT25), .B1(new_n388), .B2(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n390), .A2(new_n391), .A3(new_n356), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT25), .B1(new_n391), .B2(new_n356), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n422), .A2(new_n386), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n419), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n354), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n396), .A2(new_n416), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G8gat), .B(G36gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(G64gat), .B(G92gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n428), .B(new_n429), .Z(new_n430));
  INV_X1    g229(.A(KEYINPUT29), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n354), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT71), .B1(new_n395), .B2(new_n355), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT71), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n425), .A2(new_n434), .A3(new_n354), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n432), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n427), .B(new_n430), .C1(new_n436), .C2(new_n416), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT30), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n433), .A2(new_n435), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n416), .B1(new_n439), .B2(new_n396), .ZN(new_n440));
  INV_X1    g239(.A(new_n427), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT72), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT72), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n443), .B(new_n427), .C1(new_n436), .C2(new_n416), .ZN(new_n444));
  INV_X1    g243(.A(new_n430), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n442), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  OR2_X1    g245(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n447));
  NAND2_X1  g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(KEYINPUT74), .A2(KEYINPUT2), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AND2_X1   g249(.A1(G141gat), .A2(G148gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(G141gat), .A2(G148gat), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  OR2_X1    g253(.A1(G155gat), .A2(G162gat), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n455), .A2(KEYINPUT73), .A3(new_n448), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT73), .ZN(new_n457));
  AND2_X1   g256(.A1(G155gat), .A2(G162gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(G155gat), .A2(G162gat), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT2), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n234), .A2(KEYINPUT75), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT75), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G155gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT76), .B(G162gat), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n453), .B1(new_n458), .B2(new_n459), .ZN(new_n469));
  OAI22_X1  g268(.A1(new_n454), .A2(new_n461), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g270(.A(G134gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G127gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n227), .A2(G134gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G113gat), .B(G120gat), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n475), .B1(new_n476), .B2(KEYINPUT1), .ZN(new_n477));
  INV_X1    g276(.A(G120gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(G113gat), .ZN(new_n479));
  INV_X1    g278(.A(G113gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G120gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G127gat), .B(G134gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT1), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n477), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT77), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n477), .A2(new_n485), .A3(KEYINPUT77), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT75), .B(G155gat), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT2), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n458), .A2(new_n459), .ZN(new_n496));
  XNOR2_X1  g295(.A(G141gat), .B(G148gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n450), .A2(new_n453), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n460), .A3(new_n456), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n471), .A2(new_n490), .A3(new_n503), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n477), .A2(new_n485), .A3(KEYINPUT66), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT66), .B1(new_n477), .B2(new_n485), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n456), .A2(new_n460), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n508), .A2(new_n500), .B1(new_n495), .B2(new_n498), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(KEYINPUT4), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(G225gat), .A2(G233gat), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n499), .A2(new_n501), .A3(new_n485), .A4(new_n477), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n504), .A2(new_n510), .A3(new_n511), .A4(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT5), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n477), .A2(new_n485), .A3(KEYINPUT77), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT77), .B1(new_n477), .B2(new_n485), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n470), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n512), .ZN(new_n520));
  INV_X1    g319(.A(new_n511), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n516), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n470), .A2(new_n513), .A3(new_n486), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n477), .A2(new_n485), .A3(KEYINPUT66), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT66), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n486), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n524), .B1(new_n513), .B2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n529), .A2(new_n516), .A3(new_n511), .A4(new_n504), .ZN(new_n530));
  XOR2_X1   g329(.A(G1gat), .B(G29gat), .Z(new_n531));
  XNOR2_X1  g330(.A(G57gat), .B(G85gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n523), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT6), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n535), .B1(new_n523), .B2(new_n530), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n530), .ZN(new_n541));
  INV_X1    g340(.A(new_n535), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(KEYINPUT6), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n438), .B(new_n446), .C1(new_n540), .C2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G78gat), .B(G106gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT31), .B(G50gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n398), .A2(new_n399), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n409), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n431), .B1(new_n409), .B2(new_n550), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n502), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n470), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT29), .B1(new_n509), .B2(new_n502), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(new_n555), .B2(new_n416), .ZN(new_n556));
  INV_X1    g355(.A(G228gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(new_n353), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT3), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n405), .B(new_n414), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(new_n561), .B2(KEYINPUT29), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n559), .B1(new_n562), .B2(new_n470), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n503), .A2(new_n431), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n561), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n563), .A2(new_n565), .A3(KEYINPUT80), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT80), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT3), .B1(new_n416), .B2(new_n431), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n558), .B1(new_n568), .B2(new_n509), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n416), .B1(new_n503), .B2(new_n431), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  AOI221_X4 g370(.A(G22gat), .B1(new_n556), .B2(new_n559), .C1(new_n566), .C2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G22gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n566), .A2(new_n571), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n549), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT80), .B1(new_n563), .B2(new_n565), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n569), .A2(new_n570), .A3(new_n567), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(G22gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n574), .A2(new_n573), .A3(new_n575), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n582), .A3(new_n548), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n545), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n395), .B1(new_n505), .B2(new_n506), .ZN(new_n588));
  INV_X1    g387(.A(G227gat), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n589), .A2(new_n353), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n425), .A2(new_n507), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G15gat), .B(G43gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT68), .ZN(new_n594));
  XNOR2_X1  g393(.A(G71gat), .B(G99gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT67), .B(KEYINPUT33), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n592), .A2(KEYINPUT32), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT69), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT69), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n592), .A2(new_n602), .A3(KEYINPUT32), .A4(new_n599), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT34), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n591), .ZN(new_n606));
  INV_X1    g405(.A(new_n590), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI211_X1 g407(.A(KEYINPUT34), .B(new_n590), .C1(new_n588), .C2(new_n591), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n592), .A2(KEYINPUT32), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n592), .A2(new_n597), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n612), .A3(new_n596), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n604), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n610), .B1(new_n604), .B2(new_n613), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n587), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n604), .A2(new_n613), .ZN(new_n618));
  INV_X1    g417(.A(new_n610), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(KEYINPUT36), .A3(new_n614), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT30), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n437), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n440), .A2(new_n441), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(KEYINPUT30), .A3(new_n430), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n446), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n528), .A2(new_n513), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n509), .A2(KEYINPUT4), .A3(new_n485), .A4(new_n477), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n504), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n521), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n519), .A2(new_n512), .A3(new_n511), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT81), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n519), .A2(new_n512), .A3(KEYINPUT81), .A4(new_n511), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n631), .A2(new_n636), .A3(KEYINPUT39), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n630), .A2(new_n638), .A3(new_n521), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n637), .A2(KEYINPUT40), .A3(new_n535), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n541), .A2(new_n542), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n637), .A2(new_n535), .A3(new_n639), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT83), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT82), .B(KEYINPUT40), .ZN(new_n645));
  AND3_X1   g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n644), .B1(new_n643), .B2(new_n645), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n627), .B(new_n642), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n641), .A2(new_n537), .A3(new_n536), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n651), .B(new_n427), .C1(new_n436), .C2(new_n416), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n396), .A2(new_n561), .A3(new_n426), .ZN(new_n653));
  OAI211_X1 g452(.A(KEYINPUT37), .B(new_n653), .C1(new_n436), .C2(new_n561), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT38), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n652), .A2(new_n654), .A3(new_n655), .A4(new_n445), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n650), .A2(new_n543), .A3(new_n437), .A4(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n442), .A2(KEYINPUT37), .A3(new_n444), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n652), .A2(new_n445), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n584), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n586), .B(new_n622), .C1(new_n649), .C2(new_n661), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n584), .A2(new_n620), .A3(new_n614), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n627), .B1(new_n543), .B2(new_n650), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT35), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n584), .A2(new_n620), .A3(new_n614), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT35), .B1(new_n667), .B2(new_n545), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n662), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT84), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT84), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n662), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n351), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n540), .A2(new_n544), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n627), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n678), .A2(G8gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT102), .B(KEYINPUT16), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G8gat), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT42), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n683), .B1(KEYINPUT42), .B2(new_n682), .ZN(G1325gat));
  INV_X1    g483(.A(G15gat), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n620), .A2(new_n614), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n674), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n622), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n688), .B1(new_n691), .B2(new_n685), .ZN(G1326gat));
  NAND2_X1  g491(.A1(new_n674), .A2(new_n585), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT103), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT43), .B(G22gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  INV_X1    g495(.A(new_n294), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n697), .B1(new_n671), .B2(new_n673), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n237), .A2(new_n238), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n699), .A2(new_n328), .A3(new_n349), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n675), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n701), .A2(G29gat), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT45), .Z(new_n704));
  AND3_X1   g503(.A1(new_n662), .A2(new_n669), .A3(new_n672), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n672), .B1(new_n662), .B2(new_n669), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n294), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n670), .A2(new_n708), .A3(new_n294), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n697), .B1(new_n662), .B2(new_n669), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(KEYINPUT104), .A3(new_n708), .ZN(new_n713));
  AOI22_X1  g512(.A1(KEYINPUT44), .A2(new_n707), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n700), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT105), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AND3_X1   g515(.A1(new_n712), .A2(KEYINPUT104), .A3(new_n708), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT104), .B1(new_n712), .B2(new_n708), .ZN(new_n718));
  OAI22_X1  g517(.A1(new_n698), .A2(new_n708), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(new_n720), .A3(new_n700), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n716), .A2(new_n675), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(G29gat), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n723), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n716), .A2(new_n627), .A3(new_n721), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT106), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT106), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n716), .A2(new_n721), .A3(new_n727), .A4(new_n627), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(G36gat), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n627), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n701), .A2(G36gat), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT46), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(G1329gat));
  OR2_X1    g532(.A1(new_n686), .A2(G43gat), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n701), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n716), .A2(new_n689), .A3(new_n721), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(G43gat), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT47), .B1(new_n701), .B2(new_n734), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n719), .A2(new_n689), .A3(new_n700), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(G43gat), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI211_X1 g541(.A(KEYINPUT107), .B(new_n738), .C1(new_n739), .C2(G43gat), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n737), .A2(KEYINPUT47), .B1(new_n742), .B2(new_n743), .ZN(G1330gat));
  INV_X1    g543(.A(KEYINPUT48), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n584), .A2(G50gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n701), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n745), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n719), .A2(new_n585), .A3(new_n700), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G50gat), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n750), .B(new_n752), .C1(new_n749), .C2(new_n748), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n716), .A2(new_n585), .A3(new_n721), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n747), .B1(new_n754), .B2(G50gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n755), .B2(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g555(.A1(new_n670), .A2(new_n328), .A3(new_n295), .A4(new_n349), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n675), .ZN(new_n758));
  XOR2_X1   g557(.A(KEYINPUT109), .B(G57gat), .Z(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1332gat));
  AND2_X1   g559(.A1(new_n757), .A2(new_n627), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  AND2_X1   g561(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n761), .B2(new_n762), .ZN(G1333gat));
  NAND2_X1  g564(.A1(new_n757), .A2(new_n689), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n686), .A2(G71gat), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n766), .A2(G71gat), .B1(new_n757), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n757), .A2(new_n585), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT110), .B(G78gat), .Z(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1335gat));
  NAND2_X1  g571(.A1(new_n328), .A2(new_n239), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n773), .A2(new_n350), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n719), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(KEYINPUT111), .A3(new_n675), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n775), .B2(new_n702), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n777), .A2(new_n266), .A3(new_n779), .ZN(new_n780));
  AOI211_X1 g579(.A(new_n697), .B(new_n773), .C1(new_n662), .C2(new_n669), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(KEYINPUT51), .Z(new_n782));
  OR3_X1    g581(.A1(new_n702), .A2(new_n266), .A3(new_n350), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(G1336gat));
  NAND2_X1  g583(.A1(new_n776), .A2(new_n627), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n781), .A2(new_n786), .A3(KEYINPUT51), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n782), .B2(new_n786), .ZN(new_n788));
  INV_X1    g587(.A(G92gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n627), .A2(new_n349), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT112), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n785), .A2(G92gat), .B1(new_n788), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n789), .B1(new_n776), .B2(new_n627), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n782), .B2(new_n791), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n793), .A2(new_n794), .B1(new_n795), .B2(new_n796), .ZN(G1337gat));
  OAI21_X1  g596(.A(KEYINPUT114), .B1(new_n775), .B2(new_n622), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G99gat), .ZN(new_n799));
  NOR3_X1   g598(.A1(new_n775), .A2(KEYINPUT114), .A3(new_n622), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n687), .A2(new_n263), .A3(new_n349), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n799), .A2(new_n800), .B1(new_n782), .B2(new_n801), .ZN(G1338gat));
  NAND2_X1  g601(.A1(new_n776), .A2(new_n585), .ZN(new_n803));
  XOR2_X1   g602(.A(KEYINPUT115), .B(G106gat), .Z(new_n804));
  NOR3_X1   g603(.A1(new_n350), .A2(G106gat), .A3(new_n584), .ZN(new_n805));
  AOI22_X1  g604(.A1(new_n803), .A2(new_n804), .B1(new_n788), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807));
  INV_X1    g606(.A(new_n804), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n776), .B2(new_n585), .ZN(new_n809));
  INV_X1    g608(.A(new_n805), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n807), .B1(new_n782), .B2(new_n810), .ZN(new_n811));
  OAI22_X1  g610(.A1(new_n806), .A2(new_n807), .B1(new_n809), .B2(new_n811), .ZN(G1339gat));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n332), .A2(new_n331), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT10), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n334), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n272), .A2(new_n273), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n270), .A2(KEYINPUT96), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n816), .A2(new_n820), .A3(new_n337), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n336), .A2(new_n821), .A3(KEYINPUT54), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n346), .B1(new_n336), .B2(KEYINPUT54), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n813), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n337), .B1(new_n816), .B2(new_n820), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n345), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n336), .A2(new_n821), .A3(KEYINPUT54), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n827), .A2(KEYINPUT55), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n348), .A3(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n320), .B1(new_n307), .B2(new_n312), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n325), .A2(new_n326), .A3(new_n319), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n301), .A2(new_n303), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n260), .A2(new_n223), .A3(new_n278), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n302), .B1(new_n835), .B2(new_n300), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n317), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n832), .A2(new_n349), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n697), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n832), .A2(new_n837), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n824), .A2(new_n348), .A3(new_n829), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n294), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n699), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n295), .A2(new_n328), .A3(new_n350), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n730), .A2(new_n675), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n845), .A2(new_n667), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n329), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g648(.A1(new_n847), .A2(new_n349), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n699), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(G127gat), .ZN(G1342gat));
  AND2_X1   g652(.A1(new_n847), .A2(new_n294), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n845), .A2(new_n667), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n294), .A2(new_n730), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(G134gat), .A3(new_n702), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n855), .A2(KEYINPUT56), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT56), .B1(new_n855), .B2(new_n857), .ZN(new_n859));
  OAI22_X1  g658(.A1(new_n472), .A2(new_n854), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT116), .ZN(G1343gat));
  NOR2_X1   g660(.A1(new_n689), .A2(new_n846), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT117), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n584), .A2(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n841), .B1(new_n321), .B2(new_n327), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n832), .A2(new_n837), .A3(new_n349), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n294), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n842), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n839), .A2(KEYINPUT118), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n239), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n295), .A2(new_n328), .A3(new_n350), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n867), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n840), .A2(new_n294), .A3(new_n841), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n239), .B1(new_n870), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n875), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT57), .B1(new_n879), .B2(new_n585), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n329), .B(new_n864), .C1(new_n876), .C2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n877), .B1(new_n839), .B2(KEYINPUT118), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n870), .A2(new_n871), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n699), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n866), .B1(new_n886), .B2(new_n844), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n585), .B1(new_n843), .B2(new_n844), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n865), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n890), .A2(KEYINPUT120), .A3(new_n329), .A4(new_n864), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n883), .A2(G141gat), .A3(new_n891), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n888), .A2(new_n689), .A3(new_n846), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(G141gat), .A3(new_n328), .ZN(new_n895));
  XNOR2_X1  g694(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n892), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n881), .A2(G141gat), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT58), .B1(new_n899), .B2(new_n895), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1344gat));
  OAI211_X1 g700(.A(new_n349), .B(new_n864), .C1(new_n876), .C2(new_n880), .ZN(new_n902));
  INV_X1    g701(.A(G148gat), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n903), .A2(KEYINPUT59), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n888), .A2(new_n865), .B1(new_n879), .B2(new_n866), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n863), .A2(new_n350), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g706(.A(G148gat), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n902), .A2(new_n904), .B1(new_n908), .B2(KEYINPUT59), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n894), .A2(G148gat), .A3(new_n350), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT121), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n910), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n913));
  INV_X1    g712(.A(new_n904), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n863), .B1(new_n887), .B2(new_n889), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n349), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n879), .A2(new_n866), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n889), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n906), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n917), .B1(new_n920), .B2(G148gat), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n912), .B(new_n913), .C1(new_n916), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n911), .A2(new_n922), .ZN(G1345gat));
  AOI21_X1  g722(.A(new_n466), .B1(new_n893), .B2(new_n699), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n699), .A2(new_n466), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT122), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n924), .B1(new_n915), .B2(new_n926), .ZN(G1346gat));
  NAND2_X1  g726(.A1(new_n675), .A2(new_n493), .ZN(new_n928));
  OR4_X1    g727(.A1(new_n689), .A2(new_n888), .A3(new_n856), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n915), .A2(new_n294), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(KEYINPUT123), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n467), .B1(new_n930), .B2(KEYINPUT123), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n845), .A2(new_n675), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n667), .A2(new_n730), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n936), .A2(new_n357), .A3(new_n328), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n845), .A2(KEYINPUT124), .A3(new_n675), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(new_n329), .A3(new_n935), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n937), .B1(new_n942), .B2(new_n357), .ZN(G1348gat));
  OAI21_X1  g742(.A(G176gat), .B1(new_n936), .B2(new_n350), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n941), .A2(new_n935), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n349), .A2(new_n358), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(G1349gat));
  AND3_X1   g746(.A1(new_n699), .A2(new_n366), .A3(new_n368), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n935), .B(new_n948), .C1(new_n939), .C2(new_n940), .ZN(new_n949));
  OAI21_X1  g748(.A(G183gat), .B1(new_n936), .B2(new_n239), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n936), .B2(new_n697), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n294), .A2(new_n369), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n945), .B2(new_n955), .ZN(G1351gat));
  NOR3_X1   g755(.A1(new_n689), .A2(new_n675), .A3(new_n730), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT125), .Z(new_n958));
  NAND2_X1  g757(.A1(new_n919), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(G197gat), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n959), .A2(new_n960), .A3(new_n328), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n689), .A2(new_n730), .A3(new_n584), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n941), .A2(new_n329), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n961), .B1(new_n963), .B2(new_n960), .ZN(G1352gat));
  NOR2_X1   g763(.A1(new_n350), .A2(G204gat), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n962), .B(new_n965), .C1(new_n939), .C2(new_n940), .ZN(new_n966));
  XNOR2_X1  g765(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g768(.A(G204gat), .B1(new_n959), .B2(new_n350), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(G1353gat));
  AND2_X1   g770(.A1(new_n957), .A2(new_n699), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n410), .B1(new_n919), .B2(new_n972), .ZN(new_n973));
  OR3_X1    g772(.A1(new_n973), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n941), .A2(new_n410), .A3(new_n699), .A4(new_n962), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n973), .A2(KEYINPUT63), .ZN(new_n976));
  OAI21_X1  g775(.A(KEYINPUT127), .B1(new_n973), .B2(KEYINPUT63), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n974), .B(new_n975), .C1(new_n976), .C2(new_n977), .ZN(G1354gat));
  OAI21_X1  g777(.A(G218gat), .B1(new_n959), .B2(new_n697), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n941), .A2(new_n962), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n294), .A2(new_n411), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(G1355gat));
endmodule


