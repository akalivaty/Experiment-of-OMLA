//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT0), .A4(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n190), .A2(G146), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n188), .B2(G143), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n190), .A2(KEYINPUT64), .A3(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n192), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT67), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G134), .ZN(new_n202));
  NOR2_X1   g016(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n202), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n205), .B1(new_n207), .B2(G137), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(G137), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(G131), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n207), .A2(G137), .ZN(new_n212));
  INV_X1    g026(.A(new_n205), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(new_n203), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n214), .A2(new_n215), .A3(new_n209), .A4(new_n208), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n218), .B(new_n192), .C1(new_n197), .C2(new_n198), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n200), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(new_n189), .A3(new_n191), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n221), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n223), .B1(new_n197), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n202), .A2(new_n209), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G131), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n216), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n220), .A2(KEYINPUT30), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT30), .ZN(new_n230));
  INV_X1    g044(.A(new_n228), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n199), .B1(new_n216), .B2(new_n211), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  INV_X1    g048(.A(G119), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n234), .B1(new_n235), .B2(G116), .ZN(new_n236));
  INV_X1    g050(.A(G116), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT66), .A3(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n237), .A2(G119), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n240), .B1(new_n236), .B2(new_n238), .ZN(new_n245));
  INV_X1    g059(.A(new_n243), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n229), .A2(new_n233), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT31), .ZN(new_n250));
  NOR2_X1   g064(.A1(G237), .A2(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G210), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n252), .B(KEYINPUT27), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(G101), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n248), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n220), .A2(new_n256), .A3(new_n228), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n249), .A2(new_n250), .A3(new_n255), .A4(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT68), .ZN(new_n259));
  INV_X1    g073(.A(new_n257), .ZN(new_n260));
  INV_X1    g074(.A(new_n255), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n262), .A2(new_n263), .A3(new_n250), .A4(new_n249), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n257), .A2(KEYINPUT28), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n220), .A2(new_n267), .A3(new_n256), .A4(new_n228), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n248), .B1(new_n231), .B2(new_n232), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n249), .A2(new_n255), .A3(new_n257), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n271), .A2(new_n261), .B1(new_n272), .B2(KEYINPUT31), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(G472), .A2(G902), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n187), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n275), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n265), .B2(new_n273), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n187), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n281));
  NAND3_X1  g095(.A1(new_n277), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n220), .A2(new_n228), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n248), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n269), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n255), .A2(KEYINPUT29), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n271), .B2(new_n261), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n249), .A2(new_n257), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(new_n261), .ZN(new_n295));
  AOI211_X1 g109(.A(KEYINPUT71), .B(new_n255), .C1(new_n249), .C2(new_n257), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n289), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G472), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n283), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n291), .A2(new_n296), .A3(new_n295), .ZN(new_n301));
  OAI211_X1 g115(.A(KEYINPUT72), .B(G472), .C1(new_n301), .C2(new_n289), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n279), .A2(KEYINPUT32), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n282), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G214), .B1(G237), .B2(G902), .ZN(new_n306));
  OAI21_X1  g120(.A(G210), .B1(G237), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(G107), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT79), .B1(new_n308), .B2(G104), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT79), .ZN(new_n310));
  INV_X1    g124(.A(G104), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(G107), .ZN(new_n312));
  INV_X1    g126(.A(G101), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n308), .A2(KEYINPUT78), .A3(G104), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT3), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n308), .A2(KEYINPUT78), .A3(KEYINPUT3), .A4(G104), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n314), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n308), .A2(G104), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n311), .A2(G107), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n313), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT80), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n317), .A2(new_n318), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n309), .A2(new_n312), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(new_n313), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT80), .ZN(new_n327));
  INV_X1    g141(.A(new_n322), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n330));
  INV_X1    g144(.A(G113), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT5), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n331), .B1(new_n240), .B2(new_n332), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n330), .A2(new_n333), .B1(new_n245), .B2(new_n246), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n323), .A2(new_n329), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n324), .A2(new_n325), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT4), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G101), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n326), .A2(KEYINPUT4), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n313), .B1(new_n324), .B2(new_n325), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n338), .B(new_n248), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(G110), .B(G122), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n335), .A2(new_n341), .A3(new_n343), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(KEYINPUT6), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT6), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n342), .A2(new_n348), .A3(new_n344), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n195), .A2(new_n196), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n189), .ZN(new_n351));
  INV_X1    g165(.A(new_n224), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n189), .A2(new_n191), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n351), .A2(new_n352), .B1(new_n353), .B2(new_n222), .ZN(new_n354));
  INV_X1    g168(.A(G125), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n199), .A2(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G953), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G224), .ZN(new_n360));
  XOR2_X1   g174(.A(new_n358), .B(new_n360), .Z(new_n361));
  NAND3_X1  g175(.A1(new_n347), .A2(new_n349), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n347), .A2(KEYINPUT83), .A3(new_n349), .A4(new_n361), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(KEYINPUT84), .A2(KEYINPUT7), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n356), .A2(new_n357), .A3(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n360), .A2(KEYINPUT7), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n314), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n322), .B1(new_n371), .B2(new_n324), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n373), .A2(new_n334), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n334), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n343), .B(KEYINPUT8), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n370), .A2(new_n346), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n284), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n307), .B1(new_n366), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n307), .ZN(new_n382));
  AOI211_X1 g196(.A(new_n382), .B(new_n379), .C1(new_n364), .C2(new_n365), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n306), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G469), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n309), .A2(new_n312), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n386), .B1(new_n317), .B2(new_n318), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n326), .B(KEYINPUT4), .C1(new_n387), .C2(new_n313), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n388), .A2(new_n200), .A3(new_n219), .A4(new_n338), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n323), .A2(KEYINPUT10), .A3(new_n329), .A4(new_n225), .ZN(new_n390));
  INV_X1    g204(.A(new_n217), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n223), .B1(new_n353), .B2(new_n224), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n372), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n389), .A2(new_n390), .A3(new_n391), .A4(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G110), .B(G140), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n359), .A2(G227), .ZN(new_n398));
  XNOR2_X1  g212(.A(new_n397), .B(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  OR3_X1    g215(.A1(new_n372), .A2(KEYINPUT81), .A3(new_n225), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT81), .B1(new_n372), .B2(new_n225), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n393), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n217), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT12), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(KEYINPUT12), .A3(new_n217), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n401), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n389), .A2(new_n390), .A3(new_n395), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n217), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n400), .B1(new_n411), .B2(new_n396), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n385), .B(new_n284), .C1(new_n409), .C2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n385), .A2(new_n284), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT82), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n401), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n396), .A2(KEYINPUT82), .A3(new_n400), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n411), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n410), .A2(new_n217), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n420), .B1(new_n408), .B2(new_n407), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n421), .B2(new_n400), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n413), .B(new_n415), .C1(new_n422), .C2(new_n385), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT9), .B(G234), .ZN(new_n424));
  OAI21_X1  g238(.A(G221), .B1(new_n424), .B2(G902), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT15), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G478), .ZN(new_n428));
  OR2_X1    g242(.A1(KEYINPUT88), .A2(G122), .ZN(new_n429));
  NAND2_X1  g243(.A1(KEYINPUT88), .A2(G122), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n237), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n237), .A2(G122), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NOR3_X1   g247(.A1(new_n431), .A2(KEYINPUT89), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT89), .ZN(new_n435));
  INV_X1    g249(.A(new_n430), .ZN(new_n436));
  NOR2_X1   g250(.A1(KEYINPUT88), .A2(G122), .ZN(new_n437));
  OAI21_X1  g251(.A(G116), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n435), .B1(new_n438), .B2(new_n432), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n308), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT90), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT89), .B1(new_n431), .B2(new_n433), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n438), .A2(new_n435), .A3(new_n432), .ZN(new_n443));
  AOI21_X1  g257(.A(G107), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT90), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G128), .B(G143), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(G134), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n432), .A2(KEYINPUT14), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n449), .A2(new_n438), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n448), .B1(G107), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n441), .A2(new_n446), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(KEYINPUT13), .B1(new_n221), .B2(G143), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n454), .A2(new_n207), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(new_n447), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n434), .A2(new_n439), .A3(new_n308), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(new_n444), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G217), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n424), .A2(new_n460), .A3(G953), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n453), .A2(new_n458), .A3(new_n461), .ZN(new_n464));
  AOI21_X1  g278(.A(G902), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT91), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n428), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n465), .A2(new_n466), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n453), .A2(new_n458), .A3(new_n461), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n461), .B1(new_n453), .B2(new_n458), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n284), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT91), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n467), .B1(new_n473), .B2(new_n428), .ZN(new_n474));
  INV_X1    g288(.A(G475), .ZN(new_n475));
  XNOR2_X1  g289(.A(G125), .B(G140), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(new_n188), .ZN(new_n477));
  INV_X1    g291(.A(G237), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n359), .A3(G214), .ZN(new_n479));
  NAND2_X1  g293(.A1(KEYINPUT85), .A2(G143), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(KEYINPUT85), .A2(G143), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OR2_X1    g297(.A1(KEYINPUT85), .A2(G143), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(G214), .A3(new_n251), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT18), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(new_n215), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n484), .A2(new_n480), .B1(new_n251), .B2(G214), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n479), .A2(new_n482), .ZN(new_n490));
  OAI21_X1  g304(.A(G131), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI221_X1 g305(.A(new_n477), .B1(new_n486), .B2(new_n488), .C1(new_n491), .C2(new_n487), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n483), .A2(new_n215), .A3(new_n485), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT17), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT86), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT86), .A4(new_n495), .ZN(new_n497));
  INV_X1    g311(.A(G140), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G125), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n355), .A2(G140), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(KEYINPUT16), .ZN(new_n501));
  OR3_X1    g315(.A1(new_n355), .A2(KEYINPUT16), .A3(G140), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n502), .A3(G146), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(G146), .B1(new_n501), .B2(new_n502), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n486), .A2(KEYINPUT17), .A3(G131), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n497), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n492), .B1(new_n496), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(G113), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(new_n311), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n511), .B(new_n492), .C1(new_n496), .C2(new_n508), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n475), .B1(new_n515), .B2(new_n284), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT19), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n476), .B(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n503), .B1(new_n518), .B2(G146), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n492), .B1(new_n494), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n512), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT87), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(G475), .A2(G902), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n514), .A2(new_n521), .A3(KEYINPUT87), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT20), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT20), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n522), .A2(new_n529), .A3(new_n525), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n516), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(G234), .A2(G237), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n532), .A2(G952), .A3(new_n359), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n532), .A2(G902), .A3(G953), .ZN(new_n534));
  XNOR2_X1  g348(.A(KEYINPUT21), .B(G898), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n474), .A2(new_n531), .A3(new_n537), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n384), .A2(new_n426), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n460), .B1(G234), .B2(new_n284), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n221), .A2(G119), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n235), .A2(G128), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT24), .B(G110), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT73), .B1(new_n235), .B2(G128), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT23), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT23), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n542), .A2(KEYINPUT73), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n550), .A3(new_n543), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n551), .A2(KEYINPUT74), .A3(G110), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT74), .B1(new_n551), .B2(G110), .ZN(new_n553));
  OAI221_X1 g367(.A(new_n546), .B1(new_n505), .B2(new_n504), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n544), .A2(new_n545), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n551), .B2(G110), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n476), .A2(new_n188), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n503), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n359), .A2(G221), .A3(G234), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT75), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT22), .B(G137), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n554), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n554), .B2(new_n558), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n284), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT76), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(KEYINPUT25), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n565), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n563), .ZN(new_n571));
  INV_X1    g385(.A(new_n568), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n571), .A2(new_n284), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n541), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n540), .A2(G902), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT77), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n570), .A2(KEYINPUT77), .A3(new_n563), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n305), .A2(new_n539), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  AND3_X1   g397(.A1(new_n423), .A2(new_n581), .A3(new_n425), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n274), .A2(new_n284), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT92), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(G472), .ZN(new_n587));
  AOI21_X1  g401(.A(G902), .B1(new_n265), .B2(new_n273), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT92), .B1(new_n588), .B2(new_n299), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  AOI211_X1 g404(.A(KEYINPUT69), .B(new_n278), .C1(new_n265), .C2(new_n273), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n276), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n584), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n537), .B(new_n306), .C1(new_n381), .C2(new_n383), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n528), .A2(new_n530), .ZN(new_n595));
  INV_X1    g409(.A(new_n516), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OR3_X1    g411(.A1(new_n469), .A2(new_n470), .A3(KEYINPUT33), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT33), .B1(new_n469), .B2(new_n470), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n598), .A2(G478), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G478), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(new_n284), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n465), .B2(new_n601), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n597), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n594), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n593), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G104), .ZN(new_n609));
  XNOR2_X1  g423(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  INV_X1    g425(.A(KEYINPUT94), .ZN(new_n612));
  INV_X1    g426(.A(new_n528), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n527), .A2(KEYINPUT20), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n474), .ZN(new_n616));
  INV_X1    g430(.A(new_n614), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(KEYINPUT94), .A3(new_n528), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n615), .A2(new_n616), .A3(new_n596), .A4(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n594), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n593), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G107), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G9));
  AND2_X1   g437(.A1(new_n590), .A2(new_n592), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n384), .A2(new_n426), .ZN(new_n625));
  INV_X1    g439(.A(new_n574), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n554), .A2(new_n558), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n562), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n576), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n626), .A2(KEYINPUT95), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT95), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n634), .B1(new_n574), .B2(new_n631), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(new_n538), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n624), .A2(new_n625), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  NAND4_X1  g454(.A1(new_n633), .A2(new_n635), .A3(new_n425), .A4(new_n423), .ZN(new_n641));
  INV_X1    g455(.A(new_n304), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n642), .B1(new_n592), .B2(new_n281), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n641), .B1(new_n643), .B2(new_n303), .ZN(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n533), .B1(new_n534), .B2(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n619), .A2(new_n384), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  NAND2_X1  g463(.A1(new_n366), .A2(new_n380), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n382), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n366), .A2(new_n307), .A3(new_n380), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n653), .B(KEYINPUT38), .Z(new_n654));
  INV_X1    g468(.A(new_n306), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n626), .A2(new_n632), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n474), .A2(new_n531), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR4_X1   g472(.A1(new_n654), .A2(new_n655), .A3(new_n656), .A4(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n260), .A2(new_n255), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n286), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n284), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n261), .B1(new_n249), .B2(new_n257), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n643), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n646), .B(KEYINPUT39), .Z(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n426), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT40), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n659), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G143), .ZN(G45));
  INV_X1    g485(.A(new_n646), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n597), .A2(new_n605), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT96), .B1(new_n384), .B2(new_n673), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n531), .A2(new_n604), .A3(new_n646), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT96), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n653), .A2(new_n675), .A3(new_n676), .A4(new_n306), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n644), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  OAI21_X1  g494(.A(new_n284), .B1(new_n409), .B2(new_n412), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G469), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n425), .A3(new_n413), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n305), .A2(new_n607), .A3(new_n581), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NAND4_X1  g501(.A1(new_n620), .A2(new_n305), .A3(new_n581), .A4(new_n684), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  INV_X1    g503(.A(KEYINPUT97), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(new_n384), .B2(new_n683), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n653), .A2(KEYINPUT97), .A3(new_n306), .A4(new_n684), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n305), .A3(new_n637), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  XNOR2_X1  g509(.A(new_n657), .B(KEYINPUT99), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n287), .A2(new_n261), .B1(new_n272), .B2(KEYINPUT31), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n265), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n275), .ZN(new_n699));
  AOI22_X1  g513(.A1(KEYINPUT98), .A2(new_n699), .B1(new_n585), .B2(G472), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT98), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n698), .A2(new_n701), .A3(new_n275), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n384), .A2(new_n536), .A3(new_n683), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n696), .A2(new_n581), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NAND2_X1  g520(.A1(new_n585), .A2(G472), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n699), .A2(KEYINPUT98), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n656), .A4(new_n702), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(KEYINPUT100), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT100), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n700), .A2(new_n711), .A3(new_n656), .A4(new_n702), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n693), .A3(new_n675), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  NAND3_X1  g529(.A1(new_n651), .A2(new_n306), .A3(new_n652), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n716), .A2(new_n673), .A3(new_n426), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n717), .A2(KEYINPUT42), .ZN(new_n718));
  INV_X1    g532(.A(new_n581), .ZN(new_n719));
  OR3_X1    g533(.A1(new_n279), .A2(KEYINPUT101), .A3(KEYINPUT32), .ZN(new_n720));
  OAI21_X1  g534(.A(KEYINPUT101), .B1(new_n279), .B2(KEYINPUT32), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n720), .A2(new_n304), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n719), .B1(new_n722), .B2(new_n303), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n716), .A2(new_n426), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n305), .A2(new_n724), .A3(new_n581), .A4(new_n675), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT42), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n718), .A2(new_n723), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n215), .ZN(G33));
  NOR2_X1   g542(.A1(new_n619), .A2(new_n646), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n305), .A3(new_n581), .A4(new_n724), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G134), .ZN(G36));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n422), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT102), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n385), .B1(new_n422), .B2(new_n732), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n414), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n413), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n425), .A3(new_n666), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n624), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n597), .A2(new_n604), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT43), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n744), .A3(new_n656), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n716), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n741), .B(new_n748), .C1(new_n746), .C2(new_n745), .ZN(new_n749));
  XOR2_X1   g563(.A(KEYINPUT103), .B(G137), .Z(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G39));
  NAND2_X1  g565(.A1(new_n739), .A2(new_n425), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n753), .A2(KEYINPUT104), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(KEYINPUT104), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n739), .B(new_n425), .C1(KEYINPUT104), .C2(new_n753), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n305), .A2(new_n581), .A3(new_n673), .A4(new_n716), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G140), .ZN(G42));
  INV_X1    g574(.A(new_n716), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n684), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n581), .A2(new_n533), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n665), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n597), .A3(new_n605), .ZN(new_n765));
  INV_X1    g579(.A(G952), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n744), .A2(new_n533), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n703), .A2(new_n581), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI211_X1 g583(.A(new_n766), .B(G953), .C1(new_n769), .C2(new_n693), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n767), .A2(new_n762), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(KEYINPUT112), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n772), .A2(new_n723), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT48), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n765), .B(new_n770), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n684), .A2(new_n655), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT110), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(new_n654), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT111), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n769), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n780), .A2(KEYINPUT111), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT50), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n597), .A2(new_n605), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n772), .A2(new_n713), .B1(new_n764), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n682), .A2(new_n413), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n425), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n756), .B2(new_n757), .ZN(new_n790));
  INV_X1    g604(.A(new_n769), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n716), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n785), .B(new_n787), .C1(new_n790), .C2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n777), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n785), .A2(KEYINPUT51), .A3(new_n787), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n790), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n790), .A2(new_n798), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n800), .A3(new_n792), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(new_n801), .A3(KEYINPUT114), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n796), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT114), .B1(new_n797), .B2(new_n801), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n384), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT105), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n597), .A2(new_n474), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n806), .A2(new_n807), .A3(new_n537), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n616), .A2(new_n531), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT105), .B1(new_n594), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n809), .A2(new_n593), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n638), .A3(new_n608), .A4(new_n582), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n713), .A2(new_n717), .ZN(new_n814));
  INV_X1    g628(.A(new_n641), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n516), .A2(new_n646), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n474), .A2(new_n615), .A3(new_n618), .A4(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n305), .A2(new_n815), .A3(new_n761), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n814), .A2(new_n730), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n813), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n718), .A2(new_n723), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n725), .A2(new_n726), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n694), .A2(new_n705), .A3(new_n688), .A4(new_n685), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n820), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT106), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n644), .B1(new_n678), .B2(new_n647), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n426), .A2(new_n656), .A3(new_n646), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n665), .A2(new_n696), .A3(new_n806), .A4(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n714), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT107), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n828), .A2(new_n714), .A3(KEYINPUT107), .A4(new_n830), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT52), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n831), .A2(KEYINPUT52), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n827), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n833), .A2(new_n834), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n727), .A2(new_n824), .A3(new_n813), .A4(new_n819), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n833), .A2(KEYINPUT52), .A3(new_n834), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n840), .B1(new_n839), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT54), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n825), .A2(KEYINPUT109), .A3(new_n823), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT109), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n727), .B2(new_n824), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n813), .A2(new_n819), .A3(new_n839), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n853), .A2(new_n835), .A3(new_n836), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n846), .A2(new_n839), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n854), .B1(new_n855), .B2(KEYINPUT108), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT108), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n846), .A2(new_n858), .A3(new_n839), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n848), .A2(new_n860), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n805), .A2(new_n861), .B1(G952), .B2(G953), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n788), .A2(KEYINPUT49), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n581), .A2(new_n306), .A3(new_n425), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n743), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n654), .A2(new_n643), .A3(new_n866), .A4(new_n664), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n867), .ZN(G75));
  NOR2_X1   g682(.A1(new_n359), .A2(G952), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT115), .Z(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n837), .A2(new_n849), .A3(new_n851), .A4(new_n852), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n835), .A2(new_n826), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT53), .B1(new_n873), .B2(new_n845), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n872), .B1(new_n874), .B2(new_n858), .ZN(new_n875));
  INV_X1    g689(.A(new_n859), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n284), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT56), .B1(new_n878), .B2(G210), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n347), .A2(new_n349), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n361), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT55), .Z(new_n882));
  OR2_X1    g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n882), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n871), .B1(new_n883), .B2(new_n884), .ZN(G51));
  NAND2_X1  g699(.A1(new_n734), .A2(new_n735), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n877), .A2(new_n284), .A3(new_n886), .ZN(new_n887));
  XNOR2_X1  g701(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(new_n414), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT54), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n857), .B1(new_n856), .B2(new_n859), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n409), .A2(new_n412), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT117), .Z(new_n894));
  AOI21_X1  g708(.A(new_n887), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT118), .B1(new_n895), .B2(new_n869), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT118), .ZN(new_n897));
  INV_X1    g711(.A(new_n869), .ZN(new_n898));
  INV_X1    g712(.A(new_n894), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n855), .A2(KEYINPUT108), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n859), .A3(new_n872), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n860), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n903), .B2(new_n889), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n897), .B(new_n898), .C1(new_n904), .C2(new_n887), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n896), .A2(new_n905), .ZN(G54));
  NAND3_X1  g720(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT119), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n524), .A2(new_n526), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n907), .B2(new_n909), .ZN(new_n911));
  INV_X1    g725(.A(new_n909), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n898), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(G60));
  XNOR2_X1  g729(.A(new_n602), .B(KEYINPUT59), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n848), .B2(new_n860), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n598), .A2(new_n599), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n870), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n916), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n903), .A2(new_n921), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(KEYINPUT120), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(KEYINPUT120), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(G63));
  INV_X1    g739(.A(KEYINPUT61), .ZN(new_n926));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT60), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n901), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n870), .B1(new_n930), .B2(new_n630), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n578), .A2(new_n579), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n901), .B2(new_n929), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n926), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT121), .ZN(new_n935));
  INV_X1    g749(.A(new_n931), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT122), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n926), .B1(new_n933), .B2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n936), .B(new_n938), .C1(new_n937), .C2(new_n933), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT121), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n940), .B(new_n926), .C1(new_n931), .C2(new_n933), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n935), .A2(new_n939), .A3(new_n941), .ZN(G66));
  INV_X1    g756(.A(G224), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n535), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n824), .A2(new_n813), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n944), .B1(new_n945), .B2(G953), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n880), .B1(G898), .B2(new_n359), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT123), .Z(new_n948));
  XNOR2_X1  g762(.A(new_n946), .B(new_n948), .ZN(G69));
  NOR3_X1   g763(.A1(new_n716), .A2(new_n426), .A3(new_n667), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n810), .A2(new_n606), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n950), .A2(new_n305), .A3(new_n581), .A4(new_n951), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n749), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n670), .A2(new_n714), .A3(new_n828), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n953), .A2(new_n759), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n359), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n229), .A2(new_n233), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(new_n518), .Z(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n741), .A2(new_n806), .A3(new_n696), .A4(new_n723), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n962), .A2(new_n714), .A3(new_n828), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n749), .A2(new_n730), .ZN(new_n964));
  AND2_X1   g778(.A1(new_n759), .A2(new_n823), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n359), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n960), .B1(G900), .B2(G953), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n359), .B1(G227), .B2(G900), .ZN(new_n968));
  AOI22_X1  g782(.A1(new_n966), .A2(new_n967), .B1(KEYINPUT124), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n961), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n968), .A2(KEYINPUT124), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n970), .B(new_n971), .Z(G72));
  XNOR2_X1  g786(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n299), .A2(new_n284), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n297), .A2(new_n272), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n847), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT127), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n945), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n979), .A2(KEYINPUT126), .A3(new_n975), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT126), .B1(new_n979), .B2(new_n975), .ZN(new_n981));
  OAI211_X1 g795(.A(new_n249), .B(new_n660), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n945), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n975), .B1(new_n957), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n869), .B1(new_n984), .B2(new_n663), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n978), .A2(new_n982), .A3(new_n985), .ZN(G57));
endmodule


