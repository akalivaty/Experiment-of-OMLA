//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT88), .B(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT66), .A2(G953), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT66), .A2(G953), .ZN(new_n192));
  OAI211_X1 g006(.A(G214), .B(new_n190), .C1(new_n191), .C2(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT86), .B(G143), .Z(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G953), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT86), .A2(G143), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n196), .A2(G214), .A3(new_n190), .A4(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n198), .A3(G131), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT87), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT87), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n195), .A2(new_n198), .A3(new_n201), .A4(G131), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n195), .A2(new_n198), .ZN(new_n204));
  INV_X1    g018(.A(G131), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(G125), .B(G140), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT73), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  OR3_X1    g025(.A1(new_n209), .A2(new_n211), .A3(G140), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT16), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n211), .A2(KEYINPUT16), .A3(G140), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n214), .A2(G146), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT19), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n208), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n213), .B2(new_n218), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n207), .B(new_n217), .C1(G146), .C2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n204), .B1(new_n222), .B2(new_n205), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n208), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n213), .B2(new_n224), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n223), .B(new_n226), .C1(new_n222), .C2(new_n199), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n189), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT17), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n203), .A2(new_n229), .A3(new_n206), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n200), .A2(KEYINPUT17), .A3(new_n202), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT89), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT16), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(new_n210), .B2(new_n212), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n224), .B1(new_n234), .B2(new_n215), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n217), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT89), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n200), .A2(new_n238), .A3(KEYINPUT17), .A4(new_n202), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n230), .A2(new_n232), .A3(new_n237), .A4(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n189), .A3(new_n227), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT90), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n240), .A2(KEYINPUT90), .A3(new_n189), .A4(new_n227), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n228), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(G475), .A2(G902), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT20), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT91), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(KEYINPUT91), .B(KEYINPUT20), .C1(new_n245), .C2(new_n247), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n243), .A2(new_n244), .ZN(new_n252));
  INV_X1    g066(.A(new_n228), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT20), .B1(new_n247), .B2(KEYINPUT92), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n254), .B(new_n255), .C1(KEYINPUT92), .C2(new_n247), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n250), .A2(new_n251), .A3(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n189), .B1(new_n240), .B2(new_n227), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n243), .B2(new_n244), .ZN(new_n259));
  OAI21_X1  g073(.A(G475), .B1(new_n259), .B2(G902), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n257), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT96), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT94), .B(G952), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(G953), .ZN(new_n264));
  NAND2_X1  g078(.A1(G234), .A2(G237), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  XOR2_X1   g081(.A(KEYINPUT21), .B(G898), .Z(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(KEYINPUT95), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n196), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(G902), .A3(new_n265), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n267), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  XNOR2_X1  g090(.A(G128), .B(G143), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n276), .B1(new_n277), .B2(KEYINPUT13), .ZN(new_n278));
  INV_X1    g092(.A(G143), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G128), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n278), .B1(KEYINPUT13), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(G116), .B(G122), .ZN(new_n282));
  INV_X1    g096(.A(G107), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n282), .B(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n277), .A2(new_n276), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n281), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n277), .B(new_n276), .ZN(new_n287));
  INV_X1    g101(.A(G116), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n288), .A2(KEYINPUT14), .A3(G122), .ZN(new_n289));
  INV_X1    g103(.A(new_n282), .ZN(new_n290));
  OAI211_X1 g104(.A(G107), .B(new_n289), .C1(new_n290), .C2(KEYINPUT14), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n282), .A2(new_n283), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n293), .B(KEYINPUT93), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n286), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  XOR2_X1   g109(.A(KEYINPUT9), .B(G234), .Z(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G217), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n297), .A2(new_n298), .A3(G953), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n295), .B(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G902), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G478), .ZN(new_n304));
  OR2_X1    g118(.A1(new_n304), .A2(KEYINPUT15), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n303), .B(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n261), .A2(new_n262), .A3(new_n275), .A4(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n257), .A2(new_n275), .A3(new_n260), .A4(new_n306), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT96), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G472), .ZN(new_n311));
  XOR2_X1   g125(.A(G116), .B(G119), .Z(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT2), .B(G113), .ZN(new_n313));
  XOR2_X1   g127(.A(new_n312), .B(new_n313), .Z(new_n314));
  INV_X1    g128(.A(KEYINPUT11), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n315), .B1(new_n276), .B2(G137), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n276), .A2(G137), .ZN(new_n317));
  INV_X1    g131(.A(G137), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT11), .A3(G134), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G131), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT64), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n316), .A2(new_n319), .A3(new_n205), .A4(new_n317), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n320), .A2(KEYINPUT64), .A3(G131), .ZN(new_n325));
  XNOR2_X1  g139(.A(G143), .B(G146), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT0), .ZN(new_n327));
  INV_X1    g141(.A(G128), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT0), .B(G128), .Z(new_n330));
  OAI21_X1  g144(.A(new_n329), .B1(new_n326), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n324), .A2(new_n325), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT1), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n326), .A2(new_n333), .A3(G128), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n279), .A2(G146), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT1), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n334), .B(new_n337), .C1(G128), .C2(new_n326), .ZN(new_n338));
  INV_X1    g152(.A(new_n317), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n276), .A2(G137), .ZN(new_n340));
  OAI21_X1  g154(.A(G131), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n323), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n314), .B1(new_n332), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n343), .B(KEYINPUT70), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n332), .A2(new_n342), .A3(new_n314), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(KEYINPUT28), .ZN(new_n347));
  INV_X1    g161(.A(new_n345), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n348), .A2(KEYINPUT28), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n196), .A2(G210), .A3(new_n190), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(G101), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(KEYINPUT29), .ZN(new_n356));
  AOI21_X1  g170(.A(G902), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n332), .A2(new_n342), .A3(KEYINPUT30), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT65), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n332), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n324), .A2(new_n331), .A3(KEYINPUT65), .A4(new_n325), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n342), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT30), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n358), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n314), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n345), .ZN(new_n367));
  INV_X1    g181(.A(new_n355), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT29), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n348), .B1(new_n362), .B2(new_n365), .ZN(new_n370));
  XOR2_X1   g184(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n371));
  OAI21_X1  g185(.A(new_n349), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n369), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n311), .B1(new_n357), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT32), .ZN(new_n375));
  AOI211_X1 g189(.A(new_n368), .B(new_n348), .C1(new_n364), .C2(new_n365), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT31), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n376), .A2(KEYINPUT67), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT67), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n366), .A2(new_n355), .A3(new_n345), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(KEYINPUT31), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n372), .A2(new_n368), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n366), .A2(new_n377), .A3(new_n355), .A4(new_n345), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n378), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(G472), .A2(G902), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n375), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT69), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT67), .B1(new_n376), .B2(new_n377), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n380), .A2(new_n379), .A3(KEYINPUT31), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n390), .A2(new_n382), .A3(new_n391), .A4(new_n383), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(KEYINPUT32), .A3(new_n386), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT32), .B1(new_n392), .B2(new_n386), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT69), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n374), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  OR2_X1    g211(.A1(KEYINPUT24), .A2(G110), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT24), .A2(G110), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT71), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT71), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n402), .A3(new_n399), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G119), .B(G128), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT23), .ZN(new_n406));
  INV_X1    g220(.A(G119), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n407), .B2(G128), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n328), .A2(KEYINPUT23), .A3(G119), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n408), .B(new_n409), .C1(G119), .C2(new_n328), .ZN(new_n410));
  OAI22_X1  g224(.A1(new_n404), .A2(new_n405), .B1(G110), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n217), .A3(new_n225), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT74), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(G110), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n401), .A2(new_n405), .A3(new_n403), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT72), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n236), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n411), .A2(new_n217), .A3(KEYINPUT74), .A4(new_n225), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n414), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT75), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT75), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n414), .A2(new_n418), .A3(new_n422), .A4(new_n419), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n196), .A2(G221), .A3(G234), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT22), .B(G137), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n421), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n420), .A2(KEYINPUT75), .A3(new_n426), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n302), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n298), .B1(G234), .B2(new_n302), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT25), .ZN(new_n434));
  AOI21_X1  g248(.A(G902), .B1(new_n428), .B2(new_n429), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT76), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n433), .A2(G902), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n397), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n324), .A2(new_n325), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT80), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(KEYINPUT12), .ZN(new_n447));
  INV_X1    g261(.A(G104), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT3), .B1(new_n448), .B2(G107), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT3), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n283), .A3(G104), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n449), .B(new_n451), .C1(G104), .C2(new_n283), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n452), .A2(G101), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n283), .A2(G104), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n448), .A2(G107), .ZN(new_n455));
  OAI21_X1  g269(.A(G101), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n338), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n338), .B1(new_n453), .B2(new_n456), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n445), .B(new_n447), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n459), .A2(new_n460), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(new_n444), .ZN(new_n463));
  XOR2_X1   g277(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n464));
  OAI21_X1  g278(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n457), .A2(KEYINPUT79), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT79), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n453), .A2(new_n467), .A3(new_n456), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n466), .A2(KEYINPUT10), .A3(new_n338), .A4(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT78), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n470), .A2(KEYINPUT10), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(KEYINPUT10), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n471), .B(new_n472), .C1(new_n457), .C2(new_n458), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n452), .A2(G101), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n453), .A2(KEYINPUT4), .A3(new_n474), .ZN(new_n475));
  OR2_X1    g289(.A1(new_n474), .A2(KEYINPUT4), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n331), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n469), .A2(new_n473), .A3(new_n444), .A4(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  XOR2_X1   g293(.A(G110), .B(G140), .Z(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(KEYINPUT77), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n196), .A2(G227), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n465), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n469), .A2(new_n473), .A3(new_n477), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n445), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(new_n487), .B2(new_n478), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n443), .B(new_n302), .C1(new_n485), .C2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n484), .B1(new_n465), .B2(new_n479), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(new_n478), .A3(new_n483), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(G469), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(G469), .A2(G902), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G221), .B1(new_n297), .B2(G902), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(G214), .B1(G237), .B2(G902), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT5), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(new_n407), .A3(G116), .ZN(new_n501));
  OAI211_X1 g315(.A(G113), .B(new_n501), .C1(new_n312), .C2(new_n500), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n312), .A2(new_n313), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n466), .A2(new_n468), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n365), .A2(new_n475), .A3(new_n476), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XOR2_X1   g321(.A(G110), .B(G122), .Z(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  XOR2_X1   g324(.A(new_n504), .B(new_n457), .Z(new_n511));
  XOR2_X1   g325(.A(new_n508), .B(KEYINPUT8), .Z(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n331), .A2(new_n211), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(G125), .B2(new_n338), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT83), .B(G224), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n517), .A2(G953), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n518), .B(KEYINPUT84), .Z(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT7), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n515), .A2(KEYINPUT82), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT82), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n514), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n523), .A2(KEYINPUT7), .A3(new_n519), .A4(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n510), .A2(new_n513), .A3(new_n522), .A4(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT81), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT6), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n507), .A2(new_n508), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n530), .B1(new_n507), .B2(new_n508), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n532), .A2(new_n533), .A3(new_n509), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n523), .A2(new_n525), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(new_n519), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n302), .B(new_n527), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT85), .ZN(new_n539));
  OAI21_X1  g353(.A(G210), .B1(G237), .B2(G902), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n540), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n537), .A2(KEYINPUT85), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n499), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n310), .A2(new_n442), .A3(new_n497), .A4(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(G101), .ZN(G3));
  NAND2_X1  g360(.A1(new_n301), .A2(KEYINPUT33), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT33), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n300), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(G478), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n304), .A2(new_n302), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n301), .A2(new_n304), .A3(new_n302), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT97), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n257), .B2(new_n260), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n537), .A2(new_n540), .ZN(new_n557));
  INV_X1    g371(.A(new_n533), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n558), .A2(new_n510), .A3(new_n531), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n535), .B(new_n520), .ZN(new_n560));
  AOI21_X1  g374(.A(G902), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n542), .A3(new_n527), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n557), .A2(new_n562), .A3(new_n498), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(new_n274), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n556), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT98), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n556), .A2(KEYINPUT98), .A3(new_n564), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n385), .A2(new_n387), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n311), .B1(new_n392), .B2(new_n302), .ZN(new_n571));
  OR3_X1    g385(.A1(new_n570), .A2(new_n571), .A3(new_n496), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n441), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT99), .B(KEYINPUT100), .Z(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT34), .B(G104), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n574), .B(new_n577), .ZN(G6));
  INV_X1    g392(.A(KEYINPUT20), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n254), .A2(new_n579), .A3(new_n246), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT101), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT101), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n254), .A2(new_n582), .A3(new_n579), .A4(new_n246), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n581), .A2(new_n250), .A3(new_n251), .A4(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n306), .ZN(new_n585));
  AND4_X1   g399(.A1(new_n260), .A2(new_n564), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n573), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT35), .B(G107), .Z(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(G9));
  INV_X1    g403(.A(new_n572), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n427), .A2(KEYINPUT36), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n420), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n439), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT102), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n438), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n310), .A2(new_n544), .A3(new_n590), .A4(new_n595), .ZN(new_n596));
  XOR2_X1   g410(.A(KEYINPUT37), .B(G110), .Z(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G12));
  INV_X1    g412(.A(new_n374), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n392), .A2(KEYINPUT32), .A3(new_n386), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n600), .A2(new_n395), .A3(KEYINPUT69), .ZN(new_n601));
  INV_X1    g415(.A(new_n396), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G900), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n267), .B1(new_n273), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AND4_X1   g420(.A1(new_n260), .A2(new_n584), .A3(new_n585), .A4(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n595), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n608), .A2(new_n563), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n603), .A2(new_n607), .A3(new_n497), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G128), .ZN(G30));
  XNOR2_X1  g425(.A(new_n605), .B(KEYINPUT39), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n497), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n541), .A2(new_n543), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(KEYINPUT38), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n498), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n394), .A2(new_n396), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n302), .B1(new_n346), .B2(new_n355), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n368), .B1(new_n366), .B2(new_n345), .ZN(new_n622));
  OAI21_X1  g436(.A(G472), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n257), .A2(new_n260), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n585), .ZN(new_n627));
  NOR4_X1   g441(.A1(new_n619), .A2(new_n625), .A3(new_n595), .A4(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT103), .B(G143), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G45));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n554), .B(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n626), .A2(new_n632), .A3(new_n606), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n634), .A2(new_n603), .A3(new_n497), .A4(new_n609), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G146), .ZN(G48));
  OAI21_X1  g450(.A(new_n302), .B1(new_n485), .B2(new_n488), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(G469), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(KEYINPUT104), .A3(new_n489), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n637), .A2(new_n640), .A3(G469), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n495), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n397), .A2(new_n441), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n569), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(KEYINPUT105), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT41), .B(G113), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G15));
  INV_X1    g462(.A(new_n441), .ZN(new_n649));
  INV_X1    g463(.A(new_n495), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n639), .B2(new_n641), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n603), .A2(new_n586), .A3(new_n649), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G116), .ZN(G18));
  NOR3_X1   g467(.A1(new_n643), .A2(new_n608), .A3(new_n563), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n308), .A2(KEYINPUT96), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n308), .A2(KEYINPUT96), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n654), .B(new_n603), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT106), .B(G119), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G21));
  INV_X1    g473(.A(new_n563), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n626), .A2(new_n585), .A3(new_n651), .A4(new_n660), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n350), .A2(new_n368), .B1(KEYINPUT31), .B2(new_n380), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n387), .B1(new_n662), .B2(new_n383), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n571), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n649), .A2(new_n664), .ZN(new_n665));
  OR3_X1    g479(.A1(new_n661), .A2(new_n665), .A3(new_n274), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G122), .ZN(G24));
  NOR2_X1   g481(.A1(new_n643), .A2(new_n563), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n664), .A2(new_n595), .ZN(new_n669));
  AND4_X1   g483(.A1(KEYINPUT107), .A2(new_n626), .A3(new_n632), .A4(new_n606), .ZN(new_n670));
  AOI21_X1  g484(.A(KEYINPUT107), .B1(new_n556), .B2(new_n606), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n668), .B(new_n669), .C1(new_n670), .C2(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G125), .ZN(G27));
  NOR2_X1   g487(.A1(new_n670), .A2(new_n671), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT108), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n492), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n492), .A2(new_n675), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n676), .A2(new_n489), .A3(new_n493), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n495), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n541), .A2(new_n498), .A3(new_n543), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n388), .A2(new_n393), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n649), .B1(new_n683), .B2(new_n374), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n682), .A2(KEYINPUT42), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n397), .A2(new_n681), .A3(new_n441), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n633), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n556), .A2(KEYINPUT107), .A3(new_n606), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n687), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI211_X1 g509(.A(KEYINPUT109), .B(KEYINPUT42), .C1(new_n688), .C2(new_n692), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n686), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G131), .ZN(G33));
  NOR2_X1   g512(.A1(new_n679), .A2(new_n680), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n603), .A2(new_n649), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n607), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n276), .ZN(G36));
  INV_X1    g517(.A(new_n680), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n257), .A2(new_n260), .A3(new_n632), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT43), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n570), .A2(new_n571), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n257), .A2(new_n632), .A3(new_n708), .A4(new_n260), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n706), .A2(new_n707), .A3(new_n595), .A4(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n704), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT110), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n714), .B(new_n704), .C1(new_n710), .C2(new_n711), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n490), .A2(new_n491), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n717), .B(G469), .C1(new_n723), .C2(G902), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n721), .A2(G469), .A3(new_n722), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(KEYINPUT46), .A3(new_n493), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n724), .A2(new_n489), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n495), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n612), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n710), .A2(new_n711), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n716), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G137), .ZN(G39));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n728), .B(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n603), .A2(new_n649), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n734), .A2(new_n634), .A3(new_n704), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G140), .ZN(G42));
  AND2_X1   g551(.A1(new_n706), .A2(new_n709), .ZN(new_n738));
  INV_X1    g552(.A(new_n665), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(new_n267), .A3(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n617), .B(KEYINPUT38), .Z(new_n741));
  NOR2_X1   g555(.A1(new_n643), .A2(new_n498), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n741), .B1(new_n743), .B2(KEYINPUT114), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n743), .A2(KEYINPUT114), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n740), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n740), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n642), .B(KEYINPUT113), .Z(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n495), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n751), .B(new_n704), .C1(new_n734), .C2(new_n753), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n643), .A2(new_n680), .A3(new_n266), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n625), .A2(new_n649), .A3(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n756), .A2(new_n626), .A3(new_n632), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n738), .A2(new_n755), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(KEYINPUT116), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n757), .B1(new_n759), .B2(new_n669), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n750), .A2(new_n754), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n556), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n264), .B1(new_n756), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n759), .A2(new_n685), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n766), .A2(KEYINPUT48), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(KEYINPUT48), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n763), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n761), .A2(new_n762), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n751), .A2(new_n668), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n694), .B1(new_n674), .B2(new_n700), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT109), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n693), .A2(new_n687), .A3(new_n694), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n702), .B1(new_n777), .B2(new_n686), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n682), .A2(new_n669), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n661), .A2(new_n665), .A3(new_n274), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(new_n569), .B2(new_n644), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n626), .A2(new_n585), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n626), .B2(new_n555), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n275), .A3(new_n544), .A4(new_n573), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n781), .A2(new_n652), .A3(new_n657), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n585), .A2(new_n605), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n704), .A2(new_n260), .A3(new_n584), .A4(new_n786), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n787), .A2(KEYINPUT111), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n397), .A2(new_n496), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n608), .B1(new_n787), .B2(KEYINPUT111), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n545), .A2(new_n596), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n785), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n626), .A2(new_n608), .A3(new_n585), .A4(new_n660), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n679), .A2(new_n605), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n624), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n672), .A2(new_n610), .A3(new_n635), .A4(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n778), .A2(new_n779), .A3(new_n794), .A4(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n798), .B(KEYINPUT52), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n556), .A2(KEYINPUT98), .A3(new_n564), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT98), .B1(new_n556), .B2(new_n564), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n603), .A2(new_n649), .A3(new_n651), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n666), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n657), .A2(new_n652), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n545), .A2(new_n596), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n812), .A3(new_n791), .A4(new_n784), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n804), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(KEYINPUT53), .A3(new_n779), .A4(new_n778), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n803), .A2(new_n815), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(KEYINPUT54), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n803), .A2(new_n815), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n801), .A2(KEYINPUT112), .A3(new_n802), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(KEYINPUT54), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n772), .A2(new_n773), .A3(new_n817), .A4(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(G952), .B2(G953), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n642), .B(KEYINPUT49), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n741), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n649), .A2(new_n495), .A3(new_n498), .ZN(new_n826));
  OR4_X1    g640(.A1(new_n624), .A2(new_n825), .A3(new_n705), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n823), .A2(new_n827), .ZN(G75));
  XNOR2_X1  g642(.A(new_n559), .B(new_n536), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT55), .Z(new_n830));
  INV_X1    g644(.A(G210), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n831), .B(new_n302), .C1(new_n803), .C2(new_n815), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n832), .B2(KEYINPUT56), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n196), .A2(G952), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n816), .A2(G210), .A3(G902), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n837));
  INV_X1    g651(.A(new_n830), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n833), .A2(new_n835), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n833), .A2(KEYINPUT117), .A3(new_n835), .A4(new_n839), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(G51));
  XNOR2_X1  g658(.A(new_n816), .B(KEYINPUT54), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n493), .B(KEYINPUT57), .Z(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n485), .A2(new_n488), .ZN(new_n848));
  XOR2_X1   g662(.A(new_n848), .B(KEYINPUT118), .Z(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n302), .B1(new_n803), .B2(new_n815), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(G469), .A3(new_n723), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n834), .B1(new_n850), .B2(new_n852), .ZN(G54));
  NAND3_X1  g667(.A1(new_n851), .A2(KEYINPUT58), .A3(G475), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(new_n245), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n245), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n855), .A2(new_n856), .A3(new_n834), .ZN(G60));
  XNOR2_X1  g671(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(new_n551), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n547), .B2(new_n549), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n845), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n547), .A2(new_n549), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n817), .B2(new_n821), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n861), .B(new_n835), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(G63));
  NAND2_X1  g679(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n866));
  OR2_X1    g680(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n867));
  XNOR2_X1  g681(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n298), .A2(new_n302), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n868), .B(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n803), .B2(new_n815), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n872), .A2(new_n592), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n835), .B1(new_n872), .B2(new_n430), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n866), .B(new_n867), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n873), .A2(new_n874), .A3(KEYINPUT121), .A4(KEYINPUT61), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(G66));
  NAND3_X1  g692(.A1(new_n811), .A2(new_n812), .A3(new_n784), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n196), .ZN(new_n880));
  OAI21_X1  g694(.A(G953), .B1(new_n270), .B2(new_n517), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n534), .B1(G898), .B2(new_n196), .ZN(new_n883));
  XOR2_X1   g697(.A(KEYINPUT122), .B(KEYINPUT123), .Z(new_n884));
  XNOR2_X1  g698(.A(new_n883), .B(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n882), .B(new_n885), .ZN(G69));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n196), .B1(G227), .B2(G900), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n731), .A2(new_n736), .ZN(new_n889));
  INV_X1    g703(.A(new_n614), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n783), .A2(new_n442), .A3(new_n890), .A4(new_n704), .ZN(new_n891));
  INV_X1    g705(.A(new_n628), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n672), .A2(new_n610), .A3(new_n635), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n892), .A2(KEYINPUT62), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT62), .B1(new_n892), .B2(new_n893), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n889), .B(new_n891), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n364), .B(new_n220), .Z(new_n897));
  NOR2_X1   g711(.A1(new_n897), .A2(new_n271), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n702), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n627), .A2(new_n563), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n729), .A2(new_n902), .A3(new_n685), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n697), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n731), .A2(new_n736), .A3(new_n893), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n196), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n196), .A2(G900), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n906), .A2(KEYINPUT125), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n900), .B1(new_n913), .B2(new_n897), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n887), .B(new_n888), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n906), .A2(KEYINPUT125), .A3(new_n908), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT125), .B1(new_n906), .B2(new_n908), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n897), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n899), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT126), .B1(new_n920), .B2(KEYINPUT124), .ZN(new_n921));
  INV_X1    g735(.A(new_n888), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n920), .B2(KEYINPUT126), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n916), .B1(new_n921), .B2(new_n923), .ZN(G72));
  NOR2_X1   g738(.A1(new_n367), .A2(new_n355), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n904), .A2(new_n905), .A3(new_n879), .ZN(new_n926));
  NAND2_X1  g740(.A1(G472), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT63), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n925), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n896), .B2(new_n879), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n931), .A2(KEYINPUT127), .A3(new_n622), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT127), .B1(new_n931), .B2(new_n622), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n835), .B(new_n930), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n819), .A2(new_n820), .ZN(new_n935));
  NOR4_X1   g749(.A1(new_n935), .A2(new_n622), .A3(new_n929), .A4(new_n925), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n936), .ZN(G57));
endmodule


