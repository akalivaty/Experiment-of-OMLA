//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n543, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n588,
    new_n589, new_n592, new_n594, new_n595, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1094,
    new_n1095, new_n1096;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G236), .A3(G238), .A4(G235), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  XNOR2_X1  g029(.A(G325), .B(KEYINPUT66), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n465));
  OAI22_X1  g040(.A1(new_n460), .A2(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  OR2_X1    g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n468), .A2(new_n469), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n481), .B1(G136), .B2(new_n470), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n471), .A2(KEYINPUT70), .A3(G138), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n483), .B1(new_n460), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n478), .A2(G126), .A3(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(KEYINPUT70), .A2(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(KEYINPUT4), .C1(new_n459), .C2(new_n458), .ZN(new_n489));
  OR2_X1    g064(.A1(G102), .A2(G2105), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT69), .A2(G114), .ZN(new_n491));
  OAI21_X1  g066(.A(G2105), .B1(KEYINPUT69), .B2(G114), .ZN(new_n492));
  OAI211_X1 g067(.A(G2104), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n485), .A2(new_n486), .A3(new_n489), .A4(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OR2_X1    g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n507), .A2(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n503), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND3_X1  g092(.A1(new_n500), .A2(G63), .A3(G651), .ZN(new_n518));
  XOR2_X1   g093(.A(new_n518), .B(KEYINPUT71), .Z(new_n519));
  AOI21_X1  g094(.A(new_n497), .B1(new_n504), .B2(new_n505), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G51), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  INV_X1    g098(.A(G89), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n521), .B(new_n523), .C1(new_n524), .C2(new_n513), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n519), .A2(new_n525), .ZN(G168));
  AOI22_X1  g101(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n527), .A2(new_n502), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT72), .B(G52), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n507), .A2(new_n529), .B1(new_n513), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n528), .A2(new_n531), .ZN(G301));
  INV_X1    g107(.A(G301), .ZN(G171));
  AOI22_X1  g108(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT73), .ZN(new_n535));
  OR3_X1    g110(.A1(new_n534), .A2(new_n535), .A3(new_n502), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n534), .B2(new_n502), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n504), .A2(new_n505), .B1(new_n498), .B2(new_n499), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n538), .A2(G81), .B1(new_n520), .B2(G43), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT74), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(new_n520), .A2(G53), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT9), .ZN(new_n549));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  XOR2_X1   g125(.A(KEYINPUT75), .B(G65), .Z(new_n551));
  NOR2_X1   g126(.A1(new_n510), .A2(new_n509), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n553), .A2(G651), .B1(G91), .B2(new_n538), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n549), .A2(new_n554), .ZN(G299));
  INV_X1    g130(.A(G168), .ZN(G286));
  INV_X1    g131(.A(G74), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n498), .A2(new_n557), .A3(new_n499), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n520), .A2(G49), .B1(new_n558), .B2(G651), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n538), .B2(G87), .ZN(new_n561));
  INV_X1    g136(.A(G87), .ZN(new_n562));
  NOR3_X1   g137(.A1(new_n513), .A2(KEYINPUT76), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n559), .B1(new_n561), .B2(new_n563), .ZN(G288));
  OAI211_X1 g139(.A(G48), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n565));
  INV_X1    g140(.A(G86), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n513), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(G61), .B1(new_n510), .B2(new_n509), .ZN(new_n568));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n502), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(G305));
  XOR2_X1   g147(.A(KEYINPUT77), .B(G47), .Z(new_n573));
  AOI22_X1  g148(.A1(new_n538), .A2(G85), .B1(new_n520), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n502), .B2(new_n575), .ZN(G290));
  NAND2_X1  g151(.A1(G301), .A2(G868), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n538), .A2(G92), .ZN(new_n578));
  XOR2_X1   g153(.A(new_n578), .B(KEYINPUT10), .Z(new_n579));
  NAND2_X1  g154(.A1(G79), .A2(G543), .ZN(new_n580));
  XOR2_X1   g155(.A(KEYINPUT78), .B(G66), .Z(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n552), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(G54), .B2(new_n520), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n577), .B1(new_n585), .B2(G868), .ZN(G284));
  OAI21_X1  g161(.A(new_n577), .B1(new_n585), .B2(G868), .ZN(G321));
  INV_X1    g162(.A(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(G299), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n589), .B1(new_n588), .B2(G168), .ZN(G297));
  OAI21_X1  g165(.A(new_n589), .B1(new_n588), .B2(G168), .ZN(G280));
  INV_X1    g166(.A(G559), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n585), .B1(new_n592), .B2(G860), .ZN(G148));
  NAND2_X1  g168(.A1(new_n540), .A2(new_n588), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n584), .A2(G559), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n588), .ZN(G323));
  XNOR2_X1  g171(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g172(.A1(new_n478), .A2(new_n472), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT12), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT13), .ZN(new_n600));
  INV_X1    g175(.A(G2100), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n470), .A2(G135), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n471), .A2(G111), .ZN(new_n605));
  OAI21_X1  g180(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n606));
  INV_X1    g181(.A(G123), .ZN(new_n607));
  OAI221_X1 g182(.A(new_n604), .B1(new_n605), .B2(new_n606), .C1(new_n479), .C2(new_n607), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(G2096), .Z(new_n609));
  NAND3_X1  g184(.A1(new_n602), .A2(new_n603), .A3(new_n609), .ZN(G156));
  INV_X1    g185(.A(KEYINPUT14), .ZN(new_n611));
  XNOR2_X1  g186(.A(G2427), .B(G2438), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2430), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT15), .B(G2435), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n614), .B2(new_n613), .ZN(new_n616));
  XNOR2_X1  g191(.A(G2451), .B(G2454), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT16), .ZN(new_n618));
  XNOR2_X1  g193(.A(G1341), .B(G1348), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n616), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2443), .B(G2446), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  AND3_X1   g199(.A1(new_n623), .A2(G14), .A3(new_n624), .ZN(G401));
  XNOR2_X1  g200(.A(G2067), .B(G2678), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT79), .Z(new_n627));
  XNOR2_X1  g202(.A(G2072), .B(G2078), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT80), .Z(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2084), .B(G2090), .Z(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n628), .B(KEYINPUT17), .Z(new_n633));
  OAI211_X1 g208(.A(new_n630), .B(new_n632), .C1(new_n627), .C2(new_n633), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n631), .A2(new_n626), .A3(new_n628), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT18), .Z(new_n636));
  NAND3_X1  g211(.A1(new_n627), .A2(new_n633), .A3(new_n631), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n634), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2096), .B(G2100), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(G227));
  XOR2_X1   g215(.A(G1971), .B(G1976), .Z(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT19), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1956), .B(G2474), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1961), .B(G1966), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NOR3_X1   g221(.A1(new_n642), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n642), .A2(new_n645), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT20), .Z(new_n649));
  AOI211_X1 g224(.A(new_n647), .B(new_n649), .C1(new_n642), .C2(new_n646), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT81), .ZN(new_n651));
  XOR2_X1   g226(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1991), .B(G1996), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT82), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1981), .B(G1986), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G229));
  INV_X1    g234(.A(G16), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n660), .A2(G23), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(G288), .B2(G16), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT33), .B(G1976), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(G166), .A2(new_n660), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n660), .B2(G22), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n666), .A2(G1971), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n666), .A2(G1971), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n662), .A2(new_n663), .ZN(new_n670));
  NOR2_X1   g245(.A1(G6), .A2(G16), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n571), .B2(G16), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT32), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G1981), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n669), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT34), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  OR2_X1    g253(.A1(G25), .A2(G29), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n470), .A2(G131), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n471), .A2(G107), .ZN(new_n681));
  OAI21_X1  g256(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n682));
  INV_X1    g257(.A(G119), .ZN(new_n683));
  OAI221_X1 g258(.A(new_n680), .B1(new_n681), .B2(new_n682), .C1(new_n683), .C2(new_n479), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT83), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n679), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT35), .B(G1991), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  MUX2_X1   g268(.A(G24), .B(G290), .S(G16), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(G1986), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n677), .A2(new_n678), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT36), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT31), .B(G11), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT88), .B(G28), .Z(new_n700));
  AOI21_X1  g275(.A(G29), .B1(new_n700), .B2(KEYINPUT30), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(KEYINPUT30), .B2(new_n700), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n699), .B(new_n702), .C1(new_n608), .C2(new_n689), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n660), .A2(G21), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G168), .B2(new_n660), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT87), .B(G1966), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n703), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n660), .A2(G5), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G171), .B2(new_n660), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT89), .Z(new_n711));
  INV_X1    g286(.A(G1961), .ZN(new_n712));
  OAI221_X1 g287(.A(new_n708), .B1(new_n705), .B2(new_n707), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT90), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n711), .A2(new_n712), .ZN(new_n715));
  NOR2_X1   g290(.A1(G16), .A2(G19), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n541), .B2(G16), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n715), .B1(G1341), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n470), .A2(G140), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n471), .A2(G116), .ZN(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n721));
  INV_X1    g296(.A(G128), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n719), .B1(new_n720), .B2(new_n721), .C1(new_n722), .C2(new_n479), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n689), .A2(G26), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT28), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G2067), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n585), .A2(new_n660), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G4), .B2(new_n660), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT84), .B(G1348), .Z(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n729), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n731), .A2(new_n733), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n660), .A2(G20), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT92), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT23), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G299), .B2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1956), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n689), .A2(G27), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G164), .B2(new_n689), .ZN(new_n743));
  INV_X1    g318(.A(G2078), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n689), .A2(G32), .ZN(new_n746));
  INV_X1    g321(.A(new_n479), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G129), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n470), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT26), .Z(new_n751));
  AND3_X1   g326(.A1(new_n748), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n746), .B1(new_n752), .B2(new_n689), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n741), .A2(new_n745), .A3(new_n755), .ZN(new_n756));
  NOR4_X1   g331(.A1(new_n718), .A2(new_n735), .A3(new_n736), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n717), .A2(G1341), .ZN(new_n758));
  NOR2_X1   g333(.A1(G29), .A2(G35), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G162), .B2(G29), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G2090), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT24), .ZN(new_n764));
  INV_X1    g339(.A(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(G29), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n764), .B2(new_n765), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G160), .B2(new_n689), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT86), .Z(new_n769));
  INV_X1    g344(.A(G2084), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n689), .A2(G33), .ZN(new_n772));
  NAND2_X1  g347(.A1(G115), .A2(G2104), .ZN(new_n773));
  INV_X1    g348(.A(G127), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n773), .B1(new_n460), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n775), .A2(G2105), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT25), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n470), .A2(G139), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT85), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n772), .B1(new_n781), .B2(new_n689), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(G2072), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n761), .A2(new_n762), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(G2072), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n771), .A2(new_n783), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  AOI211_X1 g361(.A(new_n763), .B(new_n786), .C1(new_n770), .C2(new_n769), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n698), .A2(new_n714), .A3(new_n757), .A4(new_n787), .ZN(G150));
  INV_X1    g363(.A(G150), .ZN(G311));
  AOI22_X1  g364(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(new_n502), .ZN(new_n791));
  INV_X1    g366(.A(G55), .ZN(new_n792));
  INV_X1    g367(.A(G93), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n507), .A2(new_n792), .B1(new_n513), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT93), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G860), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT95), .B(KEYINPUT37), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n797), .A2(new_n540), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n541), .A2(new_n795), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT38), .Z(new_n804));
  NOR2_X1   g379(.A1(new_n584), .A2(new_n592), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(KEYINPUT39), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT94), .Z(new_n809));
  INV_X1    g384(.A(G860), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n807), .B2(KEYINPUT39), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n800), .B1(new_n809), .B2(new_n811), .ZN(G145));
  XNOR2_X1  g387(.A(new_n752), .B(new_n723), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G164), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n814), .A2(KEYINPUT96), .A3(new_n781), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n781), .B(KEYINPUT96), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n688), .B(new_n599), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n819));
  INV_X1    g394(.A(G118), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(G2105), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n470), .A2(G142), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT97), .Z(new_n823));
  AOI211_X1 g398(.A(new_n821), .B(new_n823), .C1(G130), .C2(new_n747), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n818), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT98), .Z(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n817), .B2(new_n825), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n608), .B(new_n474), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(G162), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G37), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n825), .B1(new_n817), .B2(KEYINPUT99), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(KEYINPUT99), .B2(new_n817), .ZN(new_n834));
  INV_X1    g409(.A(new_n830), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n827), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n831), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g413(.A1(new_n797), .A2(new_n588), .ZN(new_n839));
  XNOR2_X1  g414(.A(G303), .B(KEYINPUT100), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G305), .ZN(new_n841));
  XNOR2_X1  g416(.A(G288), .B(G290), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n842), .A2(new_n843), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n841), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT42), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT102), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n584), .B(G299), .Z(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT41), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n803), .B(new_n595), .ZN(new_n853));
  MUX2_X1   g428(.A(new_n851), .B(new_n852), .S(new_n853), .Z(new_n854));
  AOI21_X1  g429(.A(new_n849), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n854), .A2(new_n850), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n855), .B(new_n856), .Z(new_n857));
  OAI21_X1  g432(.A(new_n839), .B1(new_n857), .B2(new_n588), .ZN(G295));
  OAI21_X1  g433(.A(new_n839), .B1(new_n857), .B2(new_n588), .ZN(G331));
  XNOR2_X1  g434(.A(G168), .B(G171), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n803), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT104), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n803), .A2(new_n860), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n863), .A2(new_n851), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n848), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n861), .A2(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n852), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n869), .A2(new_n832), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT104), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n861), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n863), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n852), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n864), .A2(new_n861), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n848), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n870), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n865), .A2(new_n868), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n848), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n870), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n879), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n880), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n870), .A2(KEYINPUT105), .A3(new_n883), .A4(new_n879), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n884), .B2(new_n885), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT43), .B1(new_n878), .B2(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n870), .A2(new_n891), .A3(new_n877), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n888), .B(new_n890), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n887), .B1(new_n894), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g470(.A(G1384), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n494), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT45), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(KEYINPUT107), .B(G40), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n467), .A2(new_n473), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT108), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n723), .B(new_n728), .ZN(new_n905));
  INV_X1    g480(.A(G1996), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n906), .B2(new_n752), .ZN(new_n907));
  INV_X1    g482(.A(new_n902), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(G1996), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n903), .A2(new_n907), .B1(new_n752), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n910), .A2(new_n687), .A3(new_n686), .A4(new_n691), .ZN(new_n911));
  OR2_X1    g486(.A1(new_n723), .A2(G2067), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n904), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n909), .B(KEYINPUT46), .Z(new_n914));
  AND2_X1   g489(.A1(new_n905), .A2(new_n752), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n904), .B2(new_n915), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n916), .B(KEYINPUT47), .Z(new_n917));
  XNOR2_X1  g492(.A(new_n688), .B(new_n691), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n918), .A2(KEYINPUT109), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(KEYINPUT109), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n919), .A2(new_n903), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n910), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n908), .A2(G1986), .A3(G290), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n924), .B(KEYINPUT48), .Z(new_n925));
  AOI211_X1 g500(.A(new_n913), .B(new_n917), .C1(new_n923), .C2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(G290), .B(G1986), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n922), .B1(new_n902), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n896), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT45), .B1(new_n494), .B2(new_n896), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n930), .A2(new_n931), .A3(new_n901), .ZN(new_n932));
  OAI21_X1  g507(.A(KEYINPUT118), .B1(new_n932), .B2(new_n707), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n897), .A2(KEYINPUT50), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT50), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n494), .A2(new_n935), .A3(new_n896), .ZN(new_n936));
  INV_X1    g511(.A(new_n901), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n770), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n896), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n899), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT118), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(new_n706), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n933), .A2(new_n940), .A3(new_n944), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n945), .A2(G8), .A3(G168), .ZN(new_n946));
  OAI21_X1  g521(.A(G1981), .B1(new_n567), .B2(new_n570), .ZN(new_n947));
  INV_X1    g522(.A(G61), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(new_n498), .B2(new_n499), .ZN(new_n949));
  INV_X1    g524(.A(new_n569), .ZN(new_n950));
  OAI21_X1  g525(.A(G651), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1981), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n506), .A2(new_n500), .A3(G86), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n565), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n947), .A2(KEYINPUT49), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT114), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n947), .A2(new_n954), .A3(KEYINPUT114), .A4(KEYINPUT49), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(G8), .B1(new_n897), .B2(new_n901), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT49), .B1(new_n947), .B2(new_n954), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n960), .ZN(new_n964));
  OAI211_X1 g539(.A(G1976), .B(new_n559), .C1(new_n561), .C2(new_n563), .ZN(new_n965));
  INV_X1    g540(.A(G1976), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT52), .B1(G288), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n965), .B(G8), .C1(new_n897), .C2(new_n901), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n969), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT113), .B1(new_n969), .B2(KEYINPUT52), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n963), .B(new_n968), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n946), .A2(KEYINPUT63), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n932), .B2(G1971), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT111), .B1(new_n938), .B2(G2090), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n901), .B1(new_n897), .B2(KEYINPUT50), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n979));
  INV_X1    g554(.A(G2090), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n936), .ZN(new_n981));
  INV_X1    g556(.A(G1971), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n942), .A2(KEYINPUT110), .A3(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n976), .A2(new_n977), .A3(new_n981), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G303), .A2(G8), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n985), .B(KEYINPUT55), .Z(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(G8), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT112), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n984), .A2(new_n989), .A3(G8), .A4(new_n986), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n984), .A2(G8), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n974), .B(new_n991), .C1(new_n986), .C2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G8), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n938), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n978), .A2(KEYINPUT117), .A3(new_n936), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n980), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n942), .A2(new_n982), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n994), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(new_n986), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(new_n972), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n991), .A2(KEYINPUT119), .A3(new_n1002), .A4(new_n946), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT63), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n973), .B1(new_n986), .B2(new_n1000), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n988), .B2(new_n990), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT119), .B1(new_n1007), .B2(new_n946), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n993), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n991), .A2(new_n972), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G288), .A2(G1976), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT116), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n963), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n954), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n960), .B(KEYINPUT115), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1010), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1009), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT56), .B(G2072), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  OAI22_X1  g594(.A1(new_n939), .A2(G1956), .B1(new_n942), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G299), .A2(KEYINPUT121), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(G299), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1956), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n932), .A2(new_n1018), .B1(new_n938), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n897), .A2(new_n901), .ZN(new_n1030));
  AOI22_X1  g605(.A1(new_n938), .A2(new_n733), .B1(new_n728), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n585), .A3(new_n1032), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT122), .B(KEYINPUT58), .Z(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(G1341), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n942), .A2(G1996), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(KEYINPUT123), .A3(new_n541), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(KEYINPUT59), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n584), .B1(new_n1031), .B2(KEYINPUT60), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(KEYINPUT60), .B2(new_n1031), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1031), .A2(KEYINPUT60), .A3(new_n584), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT61), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1026), .A2(new_n1029), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1026), .B(new_n1033), .C1(new_n1042), .C2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n933), .A2(new_n940), .A3(G168), .A4(new_n944), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G8), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(KEYINPUT51), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n945), .A2(G286), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1051), .A2(G8), .A3(new_n1048), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1050), .B1(new_n1052), .B2(KEYINPUT51), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n942), .B2(G2078), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n938), .A2(new_n712), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n932), .A2(KEYINPUT53), .A3(new_n744), .ZN(new_n1059));
  AOI21_X1  g634(.A(G301), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(KEYINPUT54), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n473), .A2(KEYINPUT53), .A3(G40), .A4(new_n744), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT124), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n466), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n471), .B1(new_n466), .B2(new_n1063), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1062), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1066), .A2(new_n899), .A3(new_n941), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1056), .A2(new_n1067), .A3(new_n1057), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1061), .B1(G171), .B2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1059), .A2(new_n1056), .A3(G301), .A4(new_n1057), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT125), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1068), .A2(G171), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT54), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1069), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1047), .A2(new_n1054), .A3(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1054), .A2(KEYINPUT62), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1060), .B1(new_n1053), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1078), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1017), .A2(KEYINPUT120), .B1(new_n1082), .B2(new_n1007), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1009), .A2(new_n1084), .A3(new_n1016), .ZN(new_n1085));
  AOI211_X1 g660(.A(KEYINPUT126), .B(new_n929), .C1(new_n1083), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT126), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1017), .A2(KEYINPUT120), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1082), .A2(new_n1007), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1087), .B1(new_n1090), .B2(new_n928), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n926), .B1(new_n1086), .B2(new_n1091), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g667(.A1(new_n880), .A2(new_n886), .ZN(new_n1094));
  INV_X1    g668(.A(G319), .ZN(new_n1095));
  NOR3_X1   g669(.A1(G401), .A2(new_n1095), .A3(G227), .ZN(new_n1096));
  AND4_X1   g670(.A1(new_n658), .A2(new_n837), .A3(new_n1094), .A4(new_n1096), .ZN(G308));
  NAND4_X1  g671(.A1(new_n658), .A2(new_n837), .A3(new_n1094), .A4(new_n1096), .ZN(G225));
endmodule


