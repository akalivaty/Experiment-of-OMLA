//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018;
  INV_X1    g000(.A(G155gat), .ZN(new_n202));
  INV_X1    g001(.A(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G148gat), .ZN(new_n208));
  INV_X1    g007(.A(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G141gat), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(new_n205), .A2(KEYINPUT2), .ZN(new_n212));
  OAI211_X1 g011(.A(KEYINPUT74), .B(new_n206), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n206), .A2(KEYINPUT74), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT74), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n204), .A2(new_n215), .A3(new_n205), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n208), .A2(new_n210), .B1(KEYINPUT2), .B2(new_n205), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT68), .ZN(new_n219));
  INV_X1    g018(.A(G113gat), .ZN(new_n220));
  INV_X1    g019(.A(G120gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G113gat), .B2(G120gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n219), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G127gat), .B(G134gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n226), .B(new_n219), .C1(new_n222), .C2(new_n224), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n213), .A2(new_n218), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n218), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n228), .A2(new_n229), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n213), .A2(new_n218), .A3(KEYINPUT3), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n232), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G225gat), .A2(G233gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT39), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n233), .A2(new_n236), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(new_n230), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n244), .B1(new_n246), .B2(new_n241), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G1gat), .B(G29gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT0), .ZN(new_n250));
  XNOR2_X1  g049(.A(G57gat), .B(G85gat), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n250), .B(new_n251), .Z(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT78), .B(KEYINPUT39), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n240), .A2(new_n242), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n248), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT40), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n248), .A2(KEYINPUT40), .A3(new_n252), .A4(new_n254), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT5), .B1(new_n246), .B2(new_n241), .ZN(new_n259));
  INV_X1    g058(.A(new_n233), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n231), .B1(new_n260), .B2(new_n237), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n230), .A2(KEYINPUT4), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n239), .A2(new_n261), .A3(new_n241), .A4(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n232), .A2(KEYINPUT5), .A3(new_n241), .A4(new_n239), .ZN(new_n265));
  INV_X1    g064(.A(new_n252), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n257), .A2(new_n258), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G8gat), .B(G36gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(G64gat), .B(G92gat), .ZN(new_n270));
  XOR2_X1   g069(.A(new_n269), .B(new_n270), .Z(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT26), .ZN(new_n275));
  NAND2_X1  g074(.A1(G169gat), .A2(G176gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n273), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(KEYINPUT27), .B(G183gat), .ZN(new_n279));
  INV_X1    g078(.A(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  XOR2_X1   g080(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n282));
  OAI211_X1 g081(.A(new_n277), .B(new_n278), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n281), .A2(new_n282), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT25), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n288));
  INV_X1    g087(.A(G183gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n289), .B2(new_n280), .ZN(new_n290));
  NAND3_X1  g089(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT64), .B(G176gat), .ZN(new_n293));
  INV_X1    g092(.A(G169gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT23), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n296));
  OAI22_X1  g095(.A1(new_n293), .A2(new_n295), .B1(new_n296), .B2(new_n273), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n287), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n291), .B(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n290), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT25), .B1(new_n295), .B2(G176gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n273), .B1(KEYINPUT23), .B2(new_n276), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n298), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G226gat), .A2(G233gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n286), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT69), .B(G211gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT70), .B(G218gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT22), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g117(.A(G197gat), .B(G204gat), .Z(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n313), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT22), .B1(new_n314), .B2(new_n315), .ZN(new_n322));
  NOR3_X1   g121(.A1(new_n322), .A2(new_n312), .A3(new_n319), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n306), .A2(KEYINPUT66), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT66), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n298), .A2(new_n305), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n285), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(new_n308), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n309), .B(new_n324), .C1(new_n328), .C2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n328), .A2(new_n308), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n286), .A2(new_n306), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n308), .A2(KEYINPUT29), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n324), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n272), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(KEYINPUT73), .B(new_n272), .C1(new_n334), .C2(new_n339), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n335), .A2(new_n338), .ZN(new_n345));
  INV_X1    g144(.A(new_n324), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(new_n333), .A3(new_n271), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT30), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n347), .A2(new_n333), .A3(new_n350), .A4(new_n271), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n268), .B1(new_n344), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT38), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT37), .ZN(new_n355));
  AOI221_X4 g154(.A(new_n346), .B1(new_n336), .B2(new_n337), .C1(new_n328), .C2(new_n308), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n309), .B1(new_n328), .B2(new_n332), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n346), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(KEYINPUT79), .A3(new_n346), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n333), .A3(new_n355), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n272), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n354), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n355), .B1(new_n347), .B2(new_n333), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT80), .B1(new_n366), .B2(new_n271), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n363), .A2(KEYINPUT38), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT37), .B1(new_n334), .B2(new_n339), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n369), .A2(new_n370), .A3(new_n272), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n365), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n264), .A2(new_n265), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT6), .B1(new_n374), .B2(new_n252), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n267), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n264), .A2(KEYINPUT6), .A3(new_n265), .A4(new_n266), .ZN(new_n377));
  AND3_X1   g176(.A1(new_n376), .A2(new_n377), .A3(new_n348), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n353), .B1(new_n373), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G22gat), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT29), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n321), .B2(new_n323), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT75), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT3), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n318), .A2(new_n313), .A3(new_n320), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n312), .B1(new_n322), .B2(new_n319), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT75), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n233), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n235), .A2(new_n329), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n324), .ZN(new_n391));
  INV_X1    g190(.A(G228gat), .ZN(new_n392));
  INV_X1    g191(.A(G233gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT76), .B1(new_n389), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n388), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n234), .B1(new_n387), .B2(KEYINPUT75), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n260), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT76), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n394), .A4(new_n391), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n318), .A2(new_n320), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n310), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n329), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n403), .A2(new_n310), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n234), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n260), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n394), .B1(new_n408), .B2(new_n391), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n380), .B1(new_n402), .B2(new_n410), .ZN(new_n411));
  AOI211_X1 g210(.A(G22gat), .B(new_n409), .C1(new_n396), .C2(new_n401), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT77), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT31), .B(G50gat), .ZN(new_n415));
  XOR2_X1   g214(.A(new_n414), .B(new_n415), .Z(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NOR4_X1   g216(.A1(new_n411), .A2(new_n412), .A3(new_n413), .A4(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n411), .A2(new_n412), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n416), .B1(new_n419), .B2(KEYINPUT77), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n413), .B1(new_n411), .B2(new_n412), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n327), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n326), .B1(new_n298), .B2(new_n305), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n286), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n236), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n328), .A2(new_n237), .ZN(new_n427));
  INV_X1    g226(.A(G227gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n393), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT32), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n328), .A2(new_n237), .ZN(new_n433));
  AOI211_X1 g232(.A(new_n236), .B(new_n285), .C1(new_n325), .C2(new_n327), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT34), .B1(new_n435), .B2(new_n429), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n426), .A2(new_n427), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT34), .ZN(new_n438));
  INV_X1    g237(.A(new_n429), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT33), .B1(new_n435), .B2(new_n429), .ZN(new_n441));
  XNOR2_X1  g240(.A(G15gat), .B(G43gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n436), .B(new_n440), .C1(new_n441), .C2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n444), .B1(new_n430), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n438), .B1(new_n437), .B2(new_n439), .ZN(new_n448));
  AOI211_X1 g247(.A(KEYINPUT34), .B(new_n429), .C1(new_n426), .C2(new_n427), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n432), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n445), .A2(new_n450), .A3(new_n432), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(KEYINPUT36), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT36), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n445), .A2(new_n450), .A3(new_n432), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(new_n451), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n379), .A2(new_n422), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n402), .A2(new_n410), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(G22gat), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n402), .A2(new_n380), .A3(new_n410), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(KEYINPUT77), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n421), .A3(new_n417), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n419), .A2(KEYINPUT77), .A3(new_n416), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n352), .A2(new_n344), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n376), .A2(new_n377), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n456), .A2(new_n451), .ZN(new_n471));
  AND4_X1   g270(.A1(KEYINPUT81), .A2(new_n352), .A3(new_n344), .A4(new_n468), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n471), .A2(new_n472), .A3(new_n463), .A4(new_n464), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT35), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT35), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n422), .A2(new_n475), .A3(new_n471), .A4(new_n472), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n458), .A2(new_n470), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT82), .B(G29gat), .ZN(new_n478));
  INV_X1    g277(.A(G36gat), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT83), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G29gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(new_n479), .A3(KEYINPUT14), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT14), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(G29gat), .B2(G36gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT83), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT82), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(G29gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n487), .B(G36gat), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT15), .ZN(new_n492));
  INV_X1    g291(.A(G50gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(G43gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n492), .B1(new_n494), .B2(KEYINPUT84), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n480), .A2(new_n486), .A3(new_n491), .A4(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G43gat), .B(G50gat), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n488), .A2(G29gat), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n479), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n485), .B1(new_n502), .B2(new_n487), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n503), .A2(new_n497), .A3(new_n495), .A4(new_n480), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n480), .A2(new_n491), .A3(new_n486), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n492), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n499), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT16), .ZN(new_n509));
  AOI21_X1  g308(.A(G1gat), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n380), .A2(G15gat), .ZN(new_n511));
  INV_X1    g310(.A(G15gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(G22gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G8gat), .ZN(new_n516));
  INV_X1    g315(.A(G8gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n508), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n510), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n510), .B1(new_n516), .B2(new_n518), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n507), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n498), .A2(new_n496), .B1(new_n505), .B2(new_n492), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n519), .A2(new_n520), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n524), .A3(new_n504), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT13), .Z(new_n529));
  NAND3_X1  g328(.A1(new_n507), .A2(new_n521), .A3(KEYINPUT87), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n525), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n507), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n523), .A2(KEYINPUT17), .A3(new_n504), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n532), .B1(new_n536), .B2(new_n521), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n528), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT18), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n531), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n507), .A2(new_n533), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT17), .B1(new_n523), .B2(new_n504), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n521), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n543), .A2(KEYINPUT18), .A3(new_n528), .A4(new_n525), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n544), .A2(KEYINPUT86), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(KEYINPUT86), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n540), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G197gat), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT11), .B(G169gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n551), .B(KEYINPUT12), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n540), .B(new_n554), .C1(new_n545), .C2(new_n546), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n477), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(KEYINPUT41), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT92), .ZN(new_n562));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n560), .A2(KEYINPUT41), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT8), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n568), .B1(G85gat), .B2(G92gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AND2_X1   g371(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n573));
  NOR2_X1   g372(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT93), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT7), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(new_n571), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n575), .A2(KEYINPUT94), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT94), .B1(new_n575), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n570), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G99gat), .B(G106gat), .Z(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n585));
  NAND2_X1  g384(.A1(KEYINPUT93), .A2(KEYINPUT7), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n571), .B1(new_n578), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n574), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n575), .A2(KEYINPUT94), .A3(new_n579), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n583), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n592), .A3(new_n570), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n584), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n566), .B1(new_n594), .B2(new_n507), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n594), .B1(new_n541), .B2(new_n542), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT95), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n592), .B1(new_n591), .B2(new_n570), .ZN(new_n598));
  AOI211_X1 g397(.A(new_n583), .B(new_n569), .C1(new_n589), .C2(new_n590), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n600), .B1(new_n534), .B2(new_n535), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n595), .B1(new_n597), .B2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G190gat), .B(G218gat), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI211_X1 g406(.A(new_n605), .B(new_n595), .C1(new_n597), .C2(new_n603), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n565), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT20), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n612), .B(KEYINPUT89), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n611), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G71gat), .B(G78gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT88), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  XNOR2_X1  g420(.A(G57gat), .B(G64gat), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n620), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n619), .B(new_n618), .C1(new_n622), .C2(new_n623), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n627), .A2(KEYINPUT21), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n627), .B(KEYINPUT91), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n524), .B1(new_n631), .B2(KEYINPUT21), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n630), .A2(new_n632), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n617), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n635), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n637), .A2(new_n633), .A3(new_n616), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n595), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n596), .A2(KEYINPUT95), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n601), .A2(new_n602), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n605), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n604), .A2(new_n606), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n564), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n609), .A2(new_n639), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT96), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT96), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n609), .A2(new_n646), .A3(new_n649), .A4(new_n639), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT97), .B1(new_n598), .B2(new_n599), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT97), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n584), .A2(new_n652), .A3(new_n593), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n653), .A3(new_n627), .ZN(new_n654));
  INV_X1    g453(.A(new_n627), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n600), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT10), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n631), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(G230gat), .A2(G233gat), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT10), .B1(new_n654), .B2(new_n656), .ZN(new_n664));
  INV_X1    g463(.A(new_n661), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT98), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n662), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n657), .A2(new_n663), .ZN(new_n668));
  XOR2_X1   g467(.A(G120gat), .B(G148gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT99), .ZN(new_n670));
  XNOR2_X1  g469(.A(G176gat), .B(G204gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n670), .B(new_n671), .Z(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n664), .A2(new_n665), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n663), .B(KEYINPUT100), .Z(new_n677));
  OAI21_X1  g476(.A(new_n668), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n672), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT101), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT101), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n675), .A2(new_n682), .A3(new_n679), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n648), .A2(new_n650), .A3(new_n681), .A4(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n675), .A2(new_n682), .A3(new_n679), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n682), .B1(new_n675), .B2(new_n679), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n689), .A2(KEYINPUT102), .A3(new_n648), .A4(new_n650), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n558), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n468), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n376), .A2(KEYINPUT103), .A3(new_n377), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g499(.A1(new_n693), .A2(new_n467), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT16), .B(G8gat), .Z(new_n702));
  AOI21_X1  g501(.A(KEYINPUT42), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  OAI21_X1  g503(.A(G8gat), .B1(new_n693), .B2(new_n467), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(new_n706), .B2(KEYINPUT42), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT104), .ZN(G1325gat));
  NAND2_X1  g507(.A1(new_n454), .A2(new_n457), .ZN(new_n709));
  OAI21_X1  g508(.A(G15gat), .B1(new_n693), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n471), .A2(new_n512), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n710), .B1(new_n693), .B2(new_n711), .ZN(G1326gat));
  NOR3_X1   g511(.A1(new_n477), .A2(new_n422), .A3(new_n557), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n692), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT43), .B(G22gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  NAND2_X1  g515(.A1(new_n681), .A2(new_n683), .ZN(new_n717));
  INV_X1    g516(.A(new_n646), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n564), .B1(new_n644), .B2(new_n645), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n717), .A2(new_n639), .A3(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n558), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(new_n478), .A3(new_n698), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n474), .A2(new_n476), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n379), .A2(new_n422), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(new_n470), .A3(new_n709), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n720), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT106), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n731), .B(KEYINPUT44), .C1(new_n477), .C2(new_n720), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n470), .A2(KEYINPUT107), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT107), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n465), .A2(new_n469), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n458), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n725), .ZN(new_n737));
  INV_X1    g536(.A(new_n720), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n737), .A2(new_n729), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n730), .A2(new_n732), .A3(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n556), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n553), .A2(KEYINPUT105), .A3(new_n555), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n745), .A2(new_n639), .A3(new_n717), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(new_n698), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n724), .B1(new_n748), .B2(new_n478), .ZN(G1328gat));
  NAND3_X1  g548(.A1(new_n722), .A2(new_n479), .A3(new_n466), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT108), .B(KEYINPUT46), .Z(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n747), .A2(new_n466), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n753), .B2(new_n479), .ZN(G1329gat));
  INV_X1    g553(.A(new_n709), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n755), .A3(new_n746), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G43gat), .ZN(new_n757));
  INV_X1    g556(.A(G43gat), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n722), .A2(new_n758), .A3(new_n471), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT47), .B1(new_n760), .B2(KEYINPUT109), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n762), .B(new_n763), .C1(new_n757), .C2(new_n759), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n761), .A2(new_n764), .ZN(G1330gat));
  AOI21_X1  g564(.A(new_n493), .B1(new_n747), .B2(new_n465), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT48), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n713), .A2(new_n493), .A3(new_n721), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  OR3_X1    g568(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n766), .B2(new_n769), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(G1331gat));
  NAND4_X1  g571(.A1(new_n745), .A2(new_n648), .A3(new_n650), .A4(new_n717), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n736), .B2(new_n725), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n698), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT110), .B(G57gat), .Z(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(G1332gat));
  AOI21_X1  g576(.A(new_n467), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT111), .ZN(new_n780));
  NOR2_X1   g579(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(G1333gat));
  INV_X1    g581(.A(G71gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n774), .A2(new_n783), .A3(new_n471), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n774), .A2(new_n755), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n785), .B2(new_n783), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g586(.A1(new_n774), .A2(new_n465), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g588(.A1(new_n744), .A2(new_n639), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n737), .A2(new_n738), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n737), .A2(KEYINPUT51), .A3(new_n738), .A4(new_n790), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n689), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(G85gat), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n796), .A3(new_n698), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n790), .A2(new_n717), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n740), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n800), .A2(new_n698), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n797), .B1(new_n801), .B2(new_n796), .ZN(G1336gat));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n466), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G92gat), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n467), .A2(G92gat), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT52), .B1(new_n795), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n793), .A2(KEYINPUT112), .A3(new_n794), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n791), .A2(new_n809), .A3(new_n792), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n689), .A2(G92gat), .A3(new_n467), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n803), .A2(G92gat), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n807), .B1(new_n813), .B2(new_n814), .ZN(G1337gat));
  AOI21_X1  g614(.A(G99gat), .B1(new_n795), .B2(new_n471), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n755), .A2(G99gat), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n800), .B2(new_n817), .ZN(G1338gat));
  NAND2_X1  g617(.A1(new_n793), .A2(new_n794), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n422), .A2(G106gat), .A3(new_n689), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT53), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n740), .A2(new_n465), .A3(new_n799), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(G106gat), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n822), .A2(new_n823), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n821), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n822), .A2(new_n828), .A3(G106gat), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n822), .B2(G106gat), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n808), .A2(new_n810), .A3(new_n820), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n827), .B1(new_n832), .B2(new_n833), .ZN(G1339gat));
  NOR2_X1   g633(.A1(new_n684), .A2(new_n744), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n836), .B1(new_n676), .B2(new_n677), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n667), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n677), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n836), .B(new_n839), .C1(new_n664), .C2(new_n665), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n672), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(KEYINPUT55), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n675), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n841), .B1(new_n667), .B2(new_n837), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(KEYINPUT55), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT115), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n838), .A2(new_n842), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n850), .A2(new_n851), .A3(new_n675), .A4(new_n843), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n847), .A2(new_n744), .A3(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n527), .A2(new_n530), .ZN(new_n854));
  OAI22_X1  g653(.A1(new_n854), .A2(new_n529), .B1(new_n537), .B2(new_n528), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n551), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n555), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n687), .B2(new_n688), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT116), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n717), .A2(new_n860), .A3(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n720), .B1(new_n853), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n847), .A2(new_n852), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n856), .B(new_n555), .C1(new_n718), .C2(new_n719), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n639), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n835), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n698), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n471), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n465), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n872), .A2(new_n467), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(G113gat), .B1(new_n875), .B2(new_n744), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n870), .A2(new_n465), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n871), .A2(new_n466), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n471), .A3(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(new_n220), .A3(new_n557), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n876), .A2(new_n880), .ZN(G1340gat));
  AOI21_X1  g680(.A(G120gat), .B1(new_n875), .B2(new_n717), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n879), .A2(new_n221), .A3(new_n689), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(G1341gat));
  INV_X1    g683(.A(G127gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n875), .A2(new_n885), .A3(new_n639), .ZN(new_n886));
  OAI21_X1  g685(.A(G127gat), .B1(new_n879), .B2(new_n869), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1342gat));
  INV_X1    g687(.A(G134gat), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n720), .A2(new_n466), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n872), .A2(new_n889), .A3(new_n874), .A4(new_n890), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT56), .ZN(new_n892));
  OAI21_X1  g691(.A(G134gat), .B1(new_n879), .B2(new_n720), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(KEYINPUT56), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(KEYINPUT117), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n892), .B(new_n893), .C1(new_n895), .C2(new_n896), .ZN(G1343gat));
  NAND2_X1  g696(.A1(new_n709), .A2(new_n878), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT118), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n898), .A2(KEYINPUT118), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n835), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n847), .A2(new_n744), .A3(new_n852), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n859), .A3(new_n861), .ZN(new_n905));
  AOI22_X1  g704(.A1(new_n905), .A2(new_n720), .B1(new_n864), .B2(new_n866), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n906), .B2(new_n639), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT57), .B1(new_n907), .B2(new_n465), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n422), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n867), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n849), .B1(new_n845), .B2(new_n913), .ZN(new_n914));
  AOI211_X1 g713(.A(KEYINPUT119), .B(new_n841), .C1(new_n667), .C2(new_n837), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n556), .A2(new_n675), .A3(new_n843), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n858), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(new_n720), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n869), .B1(new_n912), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n911), .B1(new_n920), .B2(new_n903), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n902), .B1(new_n908), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(G141gat), .B1(new_n922), .B2(new_n557), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT122), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n755), .A2(new_n422), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT120), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n907), .A2(new_n467), .A3(new_n698), .A4(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n557), .A2(G141gat), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n924), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n927), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(KEYINPUT122), .A3(new_n928), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n923), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT58), .ZN(new_n934));
  AOI21_X1  g733(.A(KEYINPUT121), .B1(new_n931), .B2(new_n928), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n927), .A2(new_n936), .A3(new_n929), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n935), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G141gat), .B1(new_n922), .B2(new_n745), .ZN(new_n939));
  AOI22_X1  g738(.A1(new_n933), .A2(new_n934), .B1(new_n938), .B2(new_n939), .ZN(G1344gat));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n941));
  AOI211_X1 g740(.A(new_n941), .B(G148gat), .C1(new_n931), .C2(new_n717), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n922), .B2(new_n689), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n944), .B1(new_n870), .B2(new_n911), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n686), .A2(new_n557), .A3(new_n690), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n865), .A2(new_n844), .A3(new_n846), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n947), .B1(new_n918), .B2(new_n720), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n946), .B1(new_n948), .B2(new_n639), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT125), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n946), .B(new_n951), .C1(new_n948), .C2(new_n639), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n950), .A2(new_n465), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n909), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n907), .A2(KEYINPUT124), .A3(new_n910), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n945), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  OR3_X1    g755(.A1(new_n900), .A2(KEYINPUT123), .A3(new_n901), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT123), .B1(new_n900), .B2(new_n901), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n689), .A2(new_n941), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n943), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n942), .B1(new_n961), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g761(.A(G155gat), .B1(new_n922), .B2(new_n869), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n931), .A2(new_n202), .A3(new_n639), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1346gat));
  OAI21_X1  g764(.A(G162gat), .B1(new_n922), .B2(new_n720), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n907), .A2(new_n698), .A3(new_n926), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n890), .A2(new_n203), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(G1347gat));
  NAND2_X1  g768(.A1(new_n871), .A2(new_n466), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n970), .A2(new_n873), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n877), .A2(new_n971), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n972), .A2(new_n294), .A3(new_n557), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n870), .A2(new_n698), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n873), .A2(new_n465), .A3(new_n467), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n976), .A2(KEYINPUT126), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(KEYINPUT126), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n977), .A2(new_n744), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n973), .B1(new_n979), .B2(new_n294), .ZN(G1348gat));
  AND4_X1   g779(.A1(new_n293), .A2(new_n877), .A3(new_n717), .A4(new_n971), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n977), .A2(new_n717), .A3(new_n978), .ZN(new_n982));
  INV_X1    g781(.A(G176gat), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(G1349gat));
  OAI21_X1  g783(.A(G183gat), .B1(new_n972), .B2(new_n869), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n974), .A2(new_n279), .A3(new_n639), .A4(new_n975), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g786(.A(new_n987), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g787(.A(G190gat), .B1(new_n972), .B2(new_n720), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(KEYINPUT127), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT127), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n991), .B(G190gat), .C1(new_n972), .C2(new_n720), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n990), .A2(KEYINPUT61), .A3(new_n992), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT61), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n989), .A2(KEYINPUT127), .A3(new_n994), .ZN(new_n995));
  NAND4_X1  g794(.A1(new_n977), .A2(new_n280), .A3(new_n738), .A4(new_n978), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(G1351gat));
  NOR3_X1   g796(.A1(new_n755), .A2(new_n467), .A3(new_n422), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n974), .A2(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(new_n999), .ZN(new_n1000));
  AOI21_X1  g799(.A(G197gat), .B1(new_n1000), .B2(new_n744), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n755), .A2(new_n970), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n956), .A2(new_n1002), .ZN(new_n1003));
  AND2_X1   g802(.A1(new_n556), .A2(G197gat), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(G1352gat));
  NAND2_X1  g804(.A1(new_n1003), .A2(new_n717), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(G204gat), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n689), .A2(G204gat), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n974), .A2(new_n998), .A3(new_n1008), .ZN(new_n1009));
  XOR2_X1   g808(.A(new_n1009), .B(KEYINPUT62), .Z(new_n1010));
  NAND2_X1  g809(.A1(new_n1007), .A2(new_n1010), .ZN(G1353gat));
  OR3_X1    g810(.A1(new_n999), .A2(new_n314), .A3(new_n869), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n956), .A2(new_n639), .A3(new_n1002), .ZN(new_n1013));
  AND3_X1   g812(.A1(new_n1013), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1014));
  AOI21_X1  g813(.A(KEYINPUT63), .B1(new_n1013), .B2(G211gat), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(G1354gat));
  AOI21_X1  g815(.A(G218gat), .B1(new_n1000), .B2(new_n738), .ZN(new_n1017));
  AND2_X1   g816(.A1(new_n738), .A2(new_n315), .ZN(new_n1018));
  AOI21_X1  g817(.A(new_n1017), .B1(new_n1003), .B2(new_n1018), .ZN(G1355gat));
endmodule


