//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1254, new_n1255,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G107), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI22_X1  g0019(.A1(new_n202), .A2(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  XOR2_X1   g0023(.A(KEYINPUT64), .B(G238), .Z(new_n224));
  OAI211_X1 g0024(.A(new_n221), .B(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  OAI21_X1  g0027(.A(new_n213), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n216), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NOR2_X1   g0045(.A1(G20), .A2(G33), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  OR2_X1    g0047(.A1(new_n247), .A2(KEYINPUT73), .ZN(new_n248));
  XOR2_X1   g0048(.A(KEYINPUT8), .B(G58), .Z(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(KEYINPUT73), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n210), .A2(G33), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT15), .B(G87), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n251), .B1(new_n210), .B2(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n209), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(KEYINPUT67), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT67), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G1), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n259), .A2(new_n261), .A3(G13), .A4(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n255), .A2(new_n257), .B1(new_n252), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(new_n259), .A2(new_n261), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(KEYINPUT70), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT70), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n259), .A2(new_n261), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(new_n210), .ZN(new_n269));
  INV_X1    g0069(.A(new_n257), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n266), .A2(new_n269), .A3(new_n262), .A4(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G77), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n264), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G169), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT66), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT66), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G33), .A3(G41), .ZN(new_n280));
  INV_X1    g0080(.A(new_n209), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  INV_X1    g0083(.A(G45), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(new_n259), .A3(new_n261), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G244), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n283), .B2(new_n284), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n282), .A2(G274), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT72), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n288), .A2(KEYINPUT72), .A3(new_n290), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT3), .B(G33), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(G232), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(G1698), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n297), .B1(new_n218), .B2(new_n295), .C1(new_n298), .C2(new_n224), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n281), .A2(new_n277), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n293), .A2(new_n294), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n275), .B1(new_n276), .B2(new_n303), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n303), .A2(G179), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(G200), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n275), .B(new_n307), .C1(new_n308), .C2(new_n303), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n287), .A2(G226), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n311), .A2(new_n290), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n295), .A2(G222), .A3(new_n296), .ZN(new_n313));
  INV_X1    g0113(.A(G223), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n313), .B1(new_n252), .B2(new_n295), .C1(new_n298), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n301), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT68), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT68), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n312), .A2(new_n319), .A3(new_n316), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G179), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n272), .A2(G50), .ZN(new_n324));
  NOR2_X1   g0124(.A1(KEYINPUT8), .A2(G58), .ZN(new_n325));
  INV_X1    g0125(.A(G58), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(KEYINPUT69), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT69), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G58), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n325), .B1(new_n330), .B2(KEYINPUT8), .ZN(new_n331));
  INV_X1    g0131(.A(new_n253), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n246), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n257), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n263), .A2(new_n202), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n324), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n318), .A2(new_n276), .A3(new_n320), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n323), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT71), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT71), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n310), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n318), .A2(new_n320), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT9), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n346), .A2(G200), .B1(new_n347), .B2(new_n338), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n321), .A2(G190), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n324), .A2(KEYINPUT9), .A3(new_n336), .A4(new_n337), .ZN(new_n351));
  XOR2_X1   g0151(.A(new_n351), .B(KEYINPUT74), .Z(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT10), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n352), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT10), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n354), .A2(new_n348), .A3(new_n355), .A4(new_n349), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT18), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT69), .B(G58), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n206), .B1(new_n359), .B2(new_n223), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(G20), .B1(G159), .B2(new_n246), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT7), .ZN(new_n362));
  NOR2_X1   g0162(.A1(KEYINPUT3), .A2(G33), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT79), .B(G33), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n363), .B1(new_n364), .B2(KEYINPUT3), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n362), .B1(new_n365), .B2(new_n210), .ZN(new_n366));
  AND2_X1   g0166(.A1(KEYINPUT79), .A2(G33), .ZN(new_n367));
  NOR2_X1   g0167(.A1(KEYINPUT79), .A2(G33), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT3), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n363), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n369), .A2(new_n362), .A3(new_n210), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(G68), .ZN(new_n372));
  OAI211_X1 g0172(.A(KEYINPUT16), .B(new_n361), .C1(new_n366), .C2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT16), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n201), .B1(new_n330), .B2(G68), .ZN(new_n375));
  INV_X1    g0175(.A(G159), .ZN(new_n376));
  OAI22_X1  g0176(.A1(new_n375), .A2(new_n210), .B1(new_n376), .B2(new_n247), .ZN(new_n377));
  NAND2_X1  g0177(.A1(KEYINPUT3), .A2(G33), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n378), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n364), .B2(KEYINPUT3), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n210), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n362), .B1(new_n381), .B2(new_n363), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n223), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n374), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n373), .A2(new_n384), .A3(new_n257), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n271), .A2(new_n331), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n263), .B2(new_n331), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G87), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n217), .A2(G1698), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(G223), .B2(G1698), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n389), .B1(new_n365), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n301), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n282), .A2(new_n286), .A3(G232), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n394), .A2(new_n290), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G169), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(new_n395), .A3(G179), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n358), .B1(new_n388), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n388), .A2(new_n399), .A3(new_n358), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n396), .A2(G200), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n393), .A2(new_n395), .A3(G190), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n405), .A2(KEYINPUT17), .A3(new_n385), .A4(new_n387), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n385), .A2(new_n403), .A3(new_n387), .A4(new_n404), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT17), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n401), .A2(new_n402), .A3(new_n406), .A4(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n345), .A2(new_n357), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n272), .A2(G68), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n263), .A2(new_n223), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n414), .B(KEYINPUT12), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n223), .A2(G20), .ZN(new_n416));
  OAI221_X1 g0216(.A(new_n416), .B1(new_n253), .B2(new_n252), .C1(new_n247), .C2(new_n202), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n257), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT11), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT11), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(new_n420), .A3(new_n257), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n413), .A2(new_n415), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n282), .A2(new_n286), .A3(G238), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n290), .ZN(new_n426));
  AND2_X1   g0226(.A1(KEYINPUT3), .A2(G33), .ZN(new_n427));
  OAI211_X1 g0227(.A(G232), .B(G1698), .C1(new_n427), .C2(new_n363), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT75), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT75), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n295), .A2(new_n430), .A3(G232), .A4(G1698), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G97), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n295), .A2(G226), .A3(new_n296), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n429), .A2(new_n431), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n426), .B1(new_n434), .B2(new_n301), .ZN(new_n435));
  XNOR2_X1  g0235(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n435), .B(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT14), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n439), .A3(G169), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n434), .A2(new_n301), .ZN(new_n441));
  INV_X1    g0241(.A(new_n426), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n437), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT13), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n443), .B(G179), .C1(new_n444), .C2(new_n435), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n439), .B1(new_n438), .B2(G169), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n424), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n443), .B(G190), .C1(new_n444), .C2(new_n435), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n423), .ZN(new_n450));
  AOI211_X1 g0250(.A(new_n436), .B(new_n426), .C1(new_n301), .C2(new_n434), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n437), .B1(new_n441), .B2(new_n442), .ZN(new_n452));
  OAI21_X1  g0252(.A(G200), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT77), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT77), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(G200), .C1(new_n451), .C2(new_n452), .ZN(new_n456));
  AOI211_X1 g0256(.A(KEYINPUT78), .B(new_n450), .C1(new_n454), .C2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT78), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(new_n456), .ZN(new_n459));
  INV_X1    g0259(.A(new_n450), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n448), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n412), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n369), .A2(new_n370), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(G244), .A3(G1698), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(G238), .A3(new_n296), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n364), .A2(G116), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n301), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n259), .A2(new_n261), .A3(G45), .ZN(new_n470));
  OR2_X1    g0270(.A1(new_n470), .A2(G274), .ZN(new_n471));
  INV_X1    g0271(.A(G250), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n471), .A2(new_n282), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G200), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n464), .A2(new_n210), .A3(G68), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT87), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT87), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n464), .A2(new_n480), .A3(new_n210), .A4(G68), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(G97), .A3(new_n332), .ZN(new_n483));
  NOR3_X1   g0283(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n484), .B1(new_n210), .B2(new_n432), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(new_n482), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n479), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n487), .A2(new_n257), .B1(new_n263), .B2(new_n254), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n474), .B1(new_n468), .B2(new_n301), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G190), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n259), .A2(new_n261), .A3(G33), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n262), .A2(new_n270), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G87), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n477), .A2(new_n488), .A3(new_n490), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n487), .A2(new_n257), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n263), .A2(new_n254), .ZN(new_n497));
  OR2_X1    g0297(.A1(new_n492), .A2(new_n254), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n476), .A2(new_n276), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n489), .A2(new_n322), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n295), .A2(KEYINPUT4), .A3(G244), .A4(new_n296), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n505), .B(new_n506), .C1(new_n472), .C2(new_n298), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n464), .A2(G244), .A3(new_n296), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n507), .B1(new_n510), .B2(KEYINPUT83), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT83), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n508), .A2(new_n512), .A3(new_n509), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n300), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  XOR2_X1   g0314(.A(KEYINPUT5), .B(G41), .Z(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(new_n470), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n209), .B1(KEYINPUT66), .B2(new_n277), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n516), .B1(new_n280), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(G257), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(G274), .A3(new_n282), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n276), .B1(new_n514), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n520), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n518), .B2(G257), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n508), .A2(new_n512), .A3(new_n509), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n512), .B1(new_n508), .B2(new_n509), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n525), .A2(new_n526), .A3(new_n507), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n322), .B(new_n524), .C1(new_n527), .C2(new_n300), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT6), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n529), .A2(KEYINPUT80), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n529), .A2(KEYINPUT80), .ZN(new_n531));
  INV_X1    g0331(.A(G97), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(new_n218), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n530), .A2(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  XNOR2_X1  g0335(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(G97), .A3(new_n218), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G20), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT81), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n246), .A2(G77), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n210), .B1(new_n535), .B2(new_n537), .ZN(new_n543));
  INV_X1    g0343(.A(new_n541), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT81), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n380), .A2(new_n382), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G107), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n257), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n492), .A2(G97), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(G97), .B2(new_n263), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT82), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT82), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n550), .B(new_n553), .C1(G97), .C2(new_n263), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n522), .A2(new_n528), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(G190), .B(new_n524), .C1(new_n527), .C2(new_n300), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT85), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n511), .A2(new_n513), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n301), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT85), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(G190), .A4(new_n524), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n556), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n521), .B1(new_n561), .B2(new_n301), .ZN(new_n566));
  INV_X1    g0366(.A(G200), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT84), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n524), .B1(new_n527), .B2(new_n300), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT84), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(G200), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n558), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT89), .ZN(new_n574));
  OAI211_X1 g0374(.A(G270), .B(new_n282), .C1(new_n515), .C2(new_n470), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n520), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT88), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n219), .A2(new_n296), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n577), .B1(new_n365), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n295), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G303), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n464), .A2(G257), .A3(new_n296), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n464), .A2(KEYINPUT88), .A3(new_n578), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n580), .A2(new_n582), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n576), .B1(new_n585), .B2(new_n301), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n262), .A2(new_n270), .A3(new_n491), .A4(G116), .ZN(new_n587));
  INV_X1    g0387(.A(G116), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n256), .A2(new_n209), .B1(G20), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n506), .B(new_n210), .C1(G33), .C2(new_n532), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n589), .A2(KEYINPUT20), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT20), .B1(new_n589), .B2(new_n590), .ZN(new_n592));
  OAI221_X1 g0392(.A(new_n587), .B1(G116), .B2(new_n262), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n586), .A2(G179), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(G169), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n586), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n574), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n593), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n600), .A2(new_n276), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n585), .A2(new_n301), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(KEYINPUT21), .C1(new_n602), .C2(new_n576), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(KEYINPUT89), .A3(new_n594), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n586), .A2(G190), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n605), .B(new_n600), .C1(new_n567), .C2(new_n586), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n597), .B1(new_n586), .B2(new_n596), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n599), .A2(new_n604), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(G264), .B(new_n282), .C1(new_n515), .C2(new_n470), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n464), .A2(G250), .A3(new_n296), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n464), .A2(G257), .A3(G1698), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n364), .A2(G294), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n610), .B1(new_n614), .B2(new_n301), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n520), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n276), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n610), .B(new_n523), .C1(new_n614), .C2(new_n301), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n322), .ZN(new_n619));
  NAND2_X1  g0419(.A1(KEYINPUT22), .A2(G87), .ZN(new_n620));
  NOR3_X1   g0420(.A1(new_n365), .A2(G20), .A3(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n210), .B(G87), .C1(new_n427), .C2(new_n363), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT22), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n364), .A2(new_n210), .A3(G116), .ZN(new_n625));
  OAI22_X1  g0425(.A1(new_n210), .A2(G107), .B1(KEYINPUT90), .B2(KEYINPUT23), .ZN(new_n626));
  XNOR2_X1  g0426(.A(KEYINPUT90), .B(KEYINPUT23), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(G20), .A3(new_n218), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n624), .A2(new_n625), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT91), .B1(new_n621), .B2(new_n629), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n625), .A2(new_n628), .A3(new_n626), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n464), .A2(KEYINPUT22), .A3(new_n210), .A4(G87), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT91), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .A4(new_n624), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n630), .A2(KEYINPUT24), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n257), .B1(new_n630), .B2(KEYINPUT24), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n262), .A2(G107), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n638), .B(KEYINPUT25), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n218), .B2(new_n492), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n617), .B(new_n619), .C1(new_n637), .C2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n636), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n630), .A2(new_n634), .A3(KEYINPUT24), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n615), .A2(new_n308), .A3(new_n520), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n618), .B2(G200), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n608), .A2(new_n648), .ZN(new_n649));
  AND4_X1   g0449(.A1(new_n463), .A2(new_n504), .A3(new_n573), .A4(new_n649), .ZN(G372));
  NAND2_X1  g0450(.A1(new_n406), .A2(new_n409), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n305), .B(new_n304), .C1(new_n457), .C2(new_n461), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n448), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n401), .A2(new_n402), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n357), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n342), .A2(new_n344), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n595), .A2(new_n598), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n641), .A2(new_n659), .A3(new_n607), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n573), .A2(new_n504), .A3(new_n647), .A4(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n502), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n503), .A2(new_n557), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(KEYINPUT26), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n503), .B2(new_n557), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n662), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n463), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n658), .A2(new_n669), .ZN(G369));
  INV_X1    g0470(.A(G13), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G20), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n265), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n600), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT92), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n680), .B1(new_n608), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n681), .B2(new_n608), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n659), .A2(new_n607), .A3(new_n680), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n641), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n678), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n641), .B(new_n647), .C1(new_n644), .C2(new_n679), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(KEYINPUT93), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(KEYINPUT93), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n687), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n641), .A2(new_n678), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n599), .A2(new_n604), .A3(new_n607), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n679), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n699), .B1(new_n695), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n698), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n214), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n484), .A2(new_n588), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(G1), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n710), .B1(new_n207), .B2(new_n707), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT28), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n489), .A2(new_n615), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT94), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n586), .A2(G179), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT94), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n489), .A2(new_n615), .A3(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n714), .A2(new_n566), .A3(new_n715), .A4(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n586), .A2(G179), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n569), .A2(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n489), .A2(new_n615), .A3(new_n716), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n716), .B1(new_n489), .B2(new_n615), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n722), .A2(new_n725), .A3(KEYINPUT30), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n586), .A2(new_n489), .A3(G179), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n727), .A2(new_n569), .A3(new_n616), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n720), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(KEYINPUT31), .B1(new_n729), .B2(new_n678), .ZN(new_n732));
  OAI21_X1  g0532(.A(KEYINPUT95), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n729), .A2(new_n678), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT31), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT95), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n736), .A2(new_n737), .A3(new_n730), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n649), .A2(new_n573), .A3(new_n504), .A4(new_n679), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n733), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI211_X1 g0542(.A(KEYINPUT29), .B(new_n678), .C1(new_n661), .C2(new_n667), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n569), .A2(new_n276), .B1(new_n549), .B2(new_n555), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n744), .A2(new_n502), .A3(new_n495), .A4(new_n528), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT96), .B1(new_n745), .B2(new_n665), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT97), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n666), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT96), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n663), .A2(new_n749), .A3(KEYINPUT26), .ZN(new_n750));
  OAI211_X1 g0550(.A(KEYINPUT97), .B(new_n665), .C1(new_n503), .C2(new_n557), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n746), .A2(new_n748), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n641), .A2(new_n599), .A3(new_n604), .A4(new_n607), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n573), .A2(new_n504), .A3(new_n647), .A4(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n752), .A2(new_n502), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n679), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n743), .B1(new_n756), .B2(KEYINPUT29), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n742), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n712), .B1(new_n759), .B2(G1), .ZN(G364));
  AOI21_X1  g0560(.A(new_n258), .B1(new_n672), .B2(G45), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n706), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G330), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n685), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT98), .Z(new_n766));
  AOI211_X1 g0566(.A(new_n763), .B(new_n766), .C1(G330), .C2(new_n686), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n209), .B1(G20), .B2(new_n276), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n210), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n308), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(G283), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n210), .A2(new_n322), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G190), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G322), .ZN(new_n778));
  INV_X1    g0578(.A(G294), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n308), .A2(G179), .A3(G200), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n210), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n777), .A2(new_n778), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n775), .A2(new_n567), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n773), .B(new_n782), .C1(G326), .C2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n774), .A2(new_n308), .A3(G200), .ZN(new_n785));
  XOR2_X1   g0585(.A(KEYINPUT33), .B(G317), .Z(new_n786));
  INV_X1    g0586(.A(G329), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G190), .A2(G200), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n770), .A2(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n785), .A2(new_n786), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n774), .A2(new_n788), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n295), .B(new_n790), .C1(G311), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G303), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n795));
  OR2_X1    g0595(.A1(new_n795), .A2(KEYINPUT100), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(KEYINPUT100), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n784), .B(new_n793), .C1(new_n794), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n789), .A2(new_n376), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT99), .B(KEYINPUT32), .Z(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n801), .B1(new_n493), .B2(new_n795), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n800), .B2(new_n801), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n295), .B1(new_n785), .B2(new_n223), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G77), .B2(new_n792), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n771), .A2(new_n218), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G50), .B2(new_n783), .ZN(new_n807));
  INV_X1    g0607(.A(new_n781), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G97), .A2(new_n808), .B1(new_n776), .B2(new_n330), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n803), .A2(new_n805), .A3(new_n807), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n769), .B1(new_n799), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n464), .A2(new_n705), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(new_n284), .B2(new_n208), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(new_n284), .B2(new_n241), .ZN(new_n815));
  INV_X1    g0615(.A(G355), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n295), .A2(new_n214), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(G116), .B2(new_n214), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G13), .A2(G33), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(G20), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n768), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n763), .B1(new_n819), .B2(new_n824), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n811), .B(new_n825), .C1(new_n685), .C2(new_n822), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n767), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  NOR2_X1   g0628(.A1(new_n768), .A2(new_n820), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n762), .B(new_n706), .C1(new_n252), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n785), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n831), .A2(G150), .B1(new_n792), .B2(G159), .ZN(new_n832));
  INV_X1    g0632(.A(new_n783), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  INV_X1    g0634(.A(G143), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n832), .B1(new_n833), .B2(new_n834), .C1(new_n835), .C2(new_n777), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT34), .ZN(new_n837));
  INV_X1    g0637(.A(G132), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n464), .B1(new_n838), .B2(new_n789), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n781), .A2(new_n359), .B1(new_n771), .B2(new_n223), .ZN(new_n840));
  INV_X1    g0640(.A(new_n798), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n839), .B(new_n840), .C1(new_n841), .C2(G50), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n833), .A2(new_n794), .B1(new_n771), .B2(new_n493), .ZN(new_n843));
  INV_X1    g0643(.A(new_n789), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n295), .B1(new_n844), .B2(G311), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n588), .B2(new_n791), .C1(new_n772), .C2(new_n785), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n843), .B(new_n846), .C1(G107), .C2(new_n841), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G97), .A2(new_n808), .B1(new_n776), .B2(G294), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT101), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n837), .A2(new_n842), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n309), .B1(new_n275), .B2(new_n679), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n306), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n306), .B2(new_n678), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n830), .B1(new_n769), .B2(new_n850), .C1(new_n854), .C2(new_n821), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n668), .A2(new_n679), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(new_n854), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n763), .B1(new_n858), .B2(new_n742), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(new_n742), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n855), .B1(new_n860), .B2(new_n861), .ZN(G384));
  NOR2_X1   g0662(.A1(new_n265), .A2(new_n672), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT106), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n423), .A2(new_n679), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n462), .A2(new_n865), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n448), .B1(new_n423), .B2(new_n679), .C1(new_n457), .C2(new_n461), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n853), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n739), .A2(new_n736), .A3(new_n730), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n388), .A2(new_n399), .ZN(new_n871));
  INV_X1    g0671(.A(new_n676), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n388), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n873), .A3(new_n407), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n373), .A2(new_n257), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT7), .B1(new_n464), .B2(G20), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(G68), .A3(new_n371), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT16), .B1(new_n879), .B2(new_n361), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n387), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n399), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n872), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n882), .A2(new_n883), .A3(new_n407), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n875), .A2(new_n876), .B1(new_n884), .B2(KEYINPUT37), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n407), .B(KEYINPUT17), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n388), .A2(new_n399), .A3(new_n358), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n887), .A2(new_n400), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n883), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n870), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n871), .A2(new_n873), .A3(new_n407), .A4(new_n876), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n893), .B(KEYINPUT38), .C1(new_n411), .C2(new_n883), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n868), .A2(new_n869), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n864), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(new_n864), .A3(new_n897), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n873), .ZN(new_n902));
  INV_X1    g0702(.A(new_n876), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n874), .A2(new_n903), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n410), .A2(new_n902), .B1(new_n904), .B2(new_n892), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT104), .B1(new_n905), .B2(KEYINPUT38), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT104), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n904), .A2(new_n892), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n873), .B1(new_n886), .B2(new_n888), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n907), .B(new_n870), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n906), .A2(new_n910), .A3(new_n894), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n911), .A2(new_n868), .A3(KEYINPUT40), .A4(new_n869), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n901), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n463), .A2(new_n869), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n764), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n890), .A2(new_n894), .A3(KEYINPUT39), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n448), .A2(new_n678), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n866), .A2(new_n867), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n668), .A2(new_n679), .A3(new_n854), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n306), .A2(new_n678), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT102), .Z(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n895), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n654), .A2(new_n676), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n924), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n463), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT105), .B1(new_n757), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT105), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT29), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n755), .B2(new_n679), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n936), .B(new_n463), .C1(new_n938), .C2(new_n743), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n657), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n933), .B(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n863), .B1(new_n916), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n916), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n538), .A2(KEYINPUT35), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n944), .A2(G116), .A3(new_n211), .A4(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT36), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n208), .B(G77), .C1(new_n223), .C2(new_n359), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(G50), .B2(new_n223), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(new_n671), .A3(new_n268), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n943), .A2(new_n947), .A3(new_n950), .ZN(G367));
  NAND2_X1  g0751(.A1(new_n556), .A2(new_n678), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n573), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n558), .A2(new_n678), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n695), .A2(new_n702), .A3(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n956), .A2(KEYINPUT42), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n573), .A2(new_n688), .A3(new_n952), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n678), .B1(new_n958), .B2(new_n557), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(new_n956), .B2(KEYINPUT42), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n488), .A2(new_n494), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n678), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n504), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n962), .A2(new_n502), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n957), .A2(new_n960), .B1(KEYINPUT43), .B2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n967), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n955), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n698), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n970), .B(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n706), .B(KEYINPUT41), .Z(new_n974));
  INV_X1    g0774(.A(KEYINPUT44), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT107), .ZN(new_n976));
  INV_X1    g0776(.A(new_n694), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n702), .B1(new_n977), .B2(new_n692), .ZN(new_n978));
  INV_X1    g0778(.A(new_n699), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n976), .B1(new_n980), .B2(new_n971), .ZN(new_n981));
  AOI211_X1 g0781(.A(KEYINPUT107), .B(new_n955), .C1(new_n978), .C2(new_n979), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n975), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT107), .B1(new_n703), .B2(new_n955), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n980), .A2(new_n976), .A3(new_n971), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(KEYINPUT44), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT45), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n980), .B2(new_n971), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n703), .A2(KEYINPUT45), .A3(new_n955), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n983), .A2(new_n986), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n697), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n695), .B(new_n702), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(new_n687), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n994), .A2(new_n758), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n983), .A2(new_n986), .A3(new_n698), .A4(new_n990), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n992), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n974), .B1(new_n997), .B2(new_n759), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n973), .B1(new_n998), .B2(new_n762), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n823), .B1(new_n214), .B2(new_n254), .C1(new_n813), .C2(new_n237), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n1000), .A2(new_n763), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n785), .A2(new_n376), .B1(new_n791), .B2(new_n202), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n581), .B(new_n1002), .C1(G137), .C2(new_n844), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n795), .A2(new_n359), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n781), .A2(new_n223), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G150), .B2(new_n776), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n771), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n783), .A2(G143), .B1(new_n1007), .B2(G77), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n588), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n841), .A2(G116), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1010), .B1(new_n1011), .B2(KEYINPUT46), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n785), .A2(new_n779), .B1(new_n791), .B2(new_n772), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G317), .B2(new_n844), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1007), .A2(G97), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G107), .A2(new_n808), .B1(new_n776), .B2(G303), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n464), .B1(new_n783), .B2(G311), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1009), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT47), .Z(new_n1020));
  INV_X1    g0820(.A(new_n822), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1001), .B1(new_n769), .B2(new_n1020), .C1(new_n965), .C2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n999), .A2(new_n1022), .ZN(G387));
  NOR2_X1   g0823(.A1(new_n995), .A2(new_n707), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n994), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1024), .B1(new_n759), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n696), .A2(new_n822), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n709), .A2(new_n817), .B1(G107), .B2(new_n214), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n234), .A2(new_n284), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n249), .A2(new_n202), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT50), .Z(new_n1031));
  AOI211_X1 g0831(.A(G45), .B(new_n708), .C1(G68), .C2(G77), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n813), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1028), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n763), .B1(new_n1034), .B2(new_n824), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n795), .A2(new_n252), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n781), .A2(new_n254), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(G50), .C2(new_n776), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n331), .A2(new_n831), .ZN(new_n1039));
  INV_X1    g0839(.A(G150), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n791), .A2(new_n223), .B1(new_n789), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1041), .A2(new_n365), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n783), .A2(G159), .B1(new_n1007), .B2(G97), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1038), .A2(new_n1039), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n464), .B1(G326), .B2(new_n844), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n781), .A2(new_n772), .B1(new_n795), .B2(new_n779), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n831), .A2(G311), .B1(new_n792), .B2(G303), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n776), .A2(G317), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(new_n778), .C2(new_n833), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1046), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n1050), .B2(new_n1049), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1045), .B1(new_n588), .B2(new_n771), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1044), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1035), .B1(new_n1056), .B2(new_n768), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1025), .A2(new_n762), .B1(new_n1027), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1026), .A2(new_n1058), .ZN(G393));
  NAND3_X1  g0859(.A1(new_n992), .A2(new_n762), .A3(new_n996), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n823), .B1(new_n532), .B2(new_n214), .C1(new_n813), .C2(new_n244), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT108), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n763), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n792), .A2(new_n249), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n202), .B2(new_n785), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT109), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n464), .B1(new_n835), .B2(new_n789), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G150), .A2(new_n783), .B1(new_n776), .B2(G159), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT51), .Z(new_n1072));
  OAI22_X1  g0872(.A1(new_n781), .A2(new_n252), .B1(new_n771), .B2(new_n493), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n795), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(G68), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1070), .A2(new_n1072), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT110), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G311), .A2(new_n776), .B1(new_n783), .B2(G317), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT52), .Z(new_n1080));
  OAI22_X1  g0880(.A1(new_n791), .A2(new_n779), .B1(new_n789), .B2(new_n778), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n295), .B(new_n1081), .C1(G303), .C2(new_n831), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n795), .A2(new_n772), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n806), .B(new_n1083), .C1(G116), .C2(new_n808), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1080), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1078), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1065), .B1(new_n1087), .B2(new_n768), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n955), .B2(new_n1021), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n997), .A2(new_n706), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n995), .B1(new_n992), .B2(new_n996), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1060), .B(new_n1089), .C1(new_n1090), .C2(new_n1091), .ZN(G390));
  NOR2_X1   g0892(.A1(new_n929), .A2(new_n923), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n755), .A2(new_n679), .A3(new_n854), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n925), .B1(new_n1094), .B2(new_n928), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n911), .A2(new_n922), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1093), .A2(new_n921), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n853), .A2(new_n764), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n869), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1099), .A2(new_n925), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n925), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n740), .A2(new_n1102), .A3(new_n1098), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n1095), .B2(new_n1096), .C1(new_n1093), .C2(new_n921), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n920), .A2(new_n820), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n829), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n763), .B1(new_n331), .B2(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n785), .A2(new_n218), .B1(new_n791), .B2(new_n532), .ZN(new_n1110));
  AOI211_X1 g0910(.A(new_n295), .B(new_n1110), .C1(G294), .C2(new_n844), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n841), .A2(G87), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n808), .A2(G77), .B1(new_n1007), .B2(G68), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G116), .A2(new_n776), .B1(new_n783), .B2(G283), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(KEYINPUT54), .B(G143), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n785), .A2(new_n834), .B1(new_n791), .B2(new_n1116), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT114), .Z(new_n1118));
  NOR2_X1   g0918(.A1(new_n795), .A2(new_n1040), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT53), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n581), .B1(new_n1007), .B2(G50), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1118), .B(new_n1120), .C1(KEYINPUT115), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(KEYINPUT115), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G159), .A2(new_n808), .B1(new_n776), .B2(G132), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n783), .A2(G128), .B1(G125), .B2(new_n844), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1123), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1115), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1109), .B1(new_n1127), .B2(new_n768), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1106), .A2(new_n762), .B1(new_n1107), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n926), .A2(new_n928), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1102), .B1(new_n740), .B2(new_n1098), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n1100), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1099), .A2(new_n925), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1103), .A2(new_n928), .A3(new_n1094), .A4(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n935), .A2(new_n939), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n463), .A2(G330), .A3(new_n869), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT111), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n658), .A4(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT112), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n940), .A2(new_n1135), .A3(KEYINPUT112), .A4(new_n1138), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(new_n1105), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT113), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1141), .A2(KEYINPUT113), .A3(new_n1105), .A4(new_n1142), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1139), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n707), .B1(new_n1106), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1129), .B1(new_n1145), .B2(new_n1149), .ZN(G378));
  NAND2_X1  g0950(.A1(new_n357), .A2(new_n340), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n338), .A2(new_n872), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n357), .A2(new_n340), .A3(new_n1152), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1156), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1152), .B1(new_n357), .B2(new_n340), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n341), .B(new_n1153), .C1(new_n353), .C2(new_n356), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1157), .A2(new_n1161), .A3(KEYINPUT118), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT118), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT119), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n912), .A2(G330), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1164), .A2(new_n901), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n896), .A2(new_n864), .A3(new_n897), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1166), .B1(new_n1168), .B2(new_n898), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1156), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1159), .A2(new_n1160), .A3(new_n1158), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT119), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT118), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1157), .A2(new_n1161), .A3(KEYINPUT118), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1169), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1167), .B1(new_n1173), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n933), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1167), .B(new_n932), .C1(new_n1173), .C2(new_n1178), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n940), .A2(new_n1138), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1135), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1182), .B1(new_n1105), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1180), .A2(new_n1181), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1180), .A2(new_n1184), .A3(KEYINPUT57), .A4(new_n1181), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n706), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1180), .A2(new_n762), .A3(new_n1181), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n763), .B1(G50), .B2(new_n1108), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n831), .A2(G97), .B1(new_n844), .B2(G283), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n254), .B2(new_n791), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n777), .A2(new_n218), .B1(new_n833), .B2(new_n588), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n771), .A2(new_n359), .ZN(new_n1195));
  NOR4_X1   g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1005), .A4(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n365), .A2(new_n283), .ZN(new_n1197));
  OAI21_X1  g0997(.A(KEYINPUT116), .B1(new_n1197), .B2(new_n1036), .ZN(new_n1198));
  OR3_X1    g0998(.A1(new_n1197), .A2(KEYINPUT116), .A3(new_n1036), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1196), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT58), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1197), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n795), .A2(new_n1116), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT117), .Z(new_n1204));
  OAI22_X1  g1004(.A1(new_n785), .A2(new_n838), .B1(new_n791), .B2(new_n834), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G125), .B2(new_n783), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(G150), .A2(new_n808), .B1(new_n776), .B2(G128), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1204), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(KEYINPUT59), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1007), .A2(G159), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n844), .C2(G124), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1201), .B(new_n1202), .C1(new_n1209), .C2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1191), .B1(new_n1214), .B2(new_n768), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1164), .B2(new_n821), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1190), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1189), .A2(new_n1218), .ZN(G375));
  NOR2_X1   g1019(.A1(new_n1182), .A2(new_n1135), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n974), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1221), .A2(new_n1222), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n925), .A2(new_n820), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n763), .B1(G68), .B2(new_n1108), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n831), .A2(G116), .B1(new_n792), .B2(G107), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1226), .B1(new_n779), .B2(new_n833), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT120), .Z(new_n1228));
  OAI221_X1 g1028(.A(new_n581), .B1(new_n789), .B2(new_n794), .C1(new_n252), .C2(new_n771), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1037), .B(new_n1229), .C1(G283), .C2(new_n776), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(new_n532), .C2(new_n798), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT121), .Z(new_n1232));
  NAND2_X1  g1032(.A1(new_n776), .A2(G137), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1233), .B1(new_n785), .B2(new_n1116), .C1(new_n833), .C2(new_n838), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n791), .A2(new_n1040), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n365), .B(new_n1235), .C1(G128), .C2(new_n844), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1195), .B1(G50), .B2(new_n808), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1236), .B(new_n1237), .C1(new_n376), .C2(new_n798), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1234), .B1(new_n1239), .B2(KEYINPUT122), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(KEYINPUT122), .B2(new_n1239), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1232), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1225), .B1(new_n1242), .B2(new_n768), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1135), .A2(new_n762), .B1(new_n1224), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1223), .A2(new_n1244), .ZN(G381));
  INV_X1    g1045(.A(G390), .ZN(new_n1246));
  INV_X1    g1046(.A(G384), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1026), .A2(new_n827), .A3(new_n1058), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1249), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1250), .A2(G387), .A3(G381), .ZN(new_n1251));
  INV_X1    g1051(.A(G378), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1251), .A2(new_n1252), .A3(new_n1218), .A4(new_n1189), .ZN(G407));
  NAND2_X1  g1053(.A1(new_n677), .A2(G213), .ZN(new_n1254));
  OR3_X1    g1054(.A1(G375), .A2(G378), .A3(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(G407), .A2(G213), .A3(new_n1255), .ZN(G409));
  NAND3_X1  g1056(.A1(new_n999), .A2(new_n1022), .A3(G390), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G390), .B1(new_n999), .B2(new_n1022), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n827), .B1(new_n1026), .B2(new_n1058), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1258), .A2(new_n1259), .B1(new_n1249), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1259), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1249), .A2(new_n1260), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1257), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT61), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT123), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1185), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1217), .A2(new_n1267), .B1(new_n1268), .B2(new_n1222), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1190), .A2(KEYINPUT123), .A3(new_n1216), .ZN(new_n1270));
  AOI21_X1  g1070(.A(G378), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1189), .A2(G378), .A3(new_n1218), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1254), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1139), .A2(KEYINPUT60), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1220), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n940), .A2(new_n1138), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(KEYINPUT60), .A3(new_n1183), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n706), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1244), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1247), .ZN(new_n1280));
  OAI211_X1 g1080(.A(G384), .B(new_n1244), .C1(new_n1275), .C2(new_n1278), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n677), .A2(G213), .A3(G2897), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1283), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1280), .A2(new_n1281), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT62), .B1(new_n1273), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1282), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1254), .B(new_n1289), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1266), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(KEYINPUT124), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1189), .A2(G378), .A3(new_n1218), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1217), .A2(new_n1267), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1268), .A2(new_n1222), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1295), .A2(new_n1270), .A3(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1294), .B1(new_n1297), .B2(G378), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT124), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1254), .A4(new_n1289), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT62), .B1(new_n1293), .B2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1265), .B1(new_n1292), .B2(new_n1301), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1273), .A2(KEYINPUT125), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT125), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1298), .B2(new_n1254), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1287), .A2(KEYINPUT126), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT126), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1284), .B2(new_n1286), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(new_n1303), .A2(new_n1305), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT63), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1293), .A2(new_n1310), .A3(new_n1300), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1298), .A2(KEYINPUT63), .A3(new_n1254), .A4(new_n1289), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1265), .A2(KEYINPUT61), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1309), .A2(new_n1311), .A3(new_n1312), .A4(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1302), .A2(new_n1314), .ZN(G405));
  NAND2_X1  g1115(.A1(G375), .A2(new_n1252), .ZN(new_n1316));
  AOI22_X1  g1116(.A1(new_n1316), .A2(new_n1294), .B1(KEYINPUT127), .B2(new_n1282), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(KEYINPUT127), .B2(new_n1282), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT127), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1316), .A2(new_n1289), .A3(new_n1319), .A4(new_n1294), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1265), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(new_n1321), .B(new_n1322), .ZN(G402));
endmodule


