//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:19 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT29), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT72), .A2(G953), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT72), .A2(G953), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G237), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(G210), .A3(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT27), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G101), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n194), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT11), .B1(new_n197), .B2(G137), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n199));
  INV_X1    g013(.A(G137), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n197), .A2(G137), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n203), .B1(new_n202), .B2(new_n204), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT0), .A2(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(G143), .B(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT0), .A3(G128), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n209), .A3(new_n211), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT1), .B1(new_n210), .B2(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT65), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n225), .B(KEYINPUT1), .C1(new_n210), .C2(G146), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(G128), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n222), .B1(new_n227), .B2(new_n212), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT64), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n200), .B2(G134), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n200), .A2(G134), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n197), .A2(KEYINPUT64), .A3(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G131), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n199), .B1(G134), .B2(new_n200), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n197), .A2(KEYINPUT11), .A3(G137), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n203), .B(new_n204), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  OAI22_X1  g052(.A1(new_n207), .A2(new_n218), .B1(new_n228), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT68), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G119), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n243), .A3(G116), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT69), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G116), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n246), .A2(new_n248), .A3(G119), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT2), .ZN(new_n251));
  INV_X1    g065(.A(G113), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT67), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(KEYINPUT2), .B2(G113), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT2), .A2(G113), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n250), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n244), .A2(new_n249), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n253), .A2(new_n255), .B1(KEYINPUT2), .B2(G113), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT70), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AND4_X1   g076(.A1(KEYINPUT70), .A2(new_n261), .A3(new_n244), .A4(new_n249), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n239), .A2(new_n264), .ZN(new_n265));
  OR2_X1    g079(.A1(new_n265), .A2(KEYINPUT28), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n228), .B2(new_n238), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n234), .A2(new_n237), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n226), .A2(G128), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n225), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n212), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n221), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n269), .A2(new_n273), .A3(KEYINPUT66), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n217), .B(new_n215), .C1(new_n205), .C2(new_n206), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n268), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n265), .B1(new_n264), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT73), .B(KEYINPUT28), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n196), .B(new_n266), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT30), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n204), .B1(new_n235), .B2(new_n236), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G131), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n237), .ZN(new_n284));
  INV_X1    g098(.A(new_n218), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n273), .A2(new_n269), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT71), .B1(new_n286), .B2(KEYINPUT30), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n269), .A2(new_n273), .ZN(new_n288));
  AND4_X1   g102(.A1(KEYINPUT71), .A2(new_n288), .A3(KEYINPUT30), .A4(new_n275), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n281), .B(new_n264), .C1(new_n287), .C2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n250), .B2(new_n258), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n261), .A2(KEYINPUT70), .A3(new_n244), .A4(new_n249), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n288), .A2(new_n294), .A3(new_n275), .A4(new_n259), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n188), .B(new_n279), .C1(new_n296), .C2(new_n196), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n239), .A2(new_n264), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT74), .A3(new_n295), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT74), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n239), .A2(new_n264), .A3(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(KEYINPUT28), .A3(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n302), .A2(KEYINPUT29), .A3(new_n196), .A4(new_n266), .ZN(new_n303));
  INV_X1    g117(.A(G902), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n187), .B1(new_n297), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n266), .B1(new_n277), .B2(new_n278), .ZN(new_n307));
  INV_X1    g121(.A(new_n196), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n265), .ZN(new_n310));
  AND3_X1   g124(.A1(new_n290), .A2(KEYINPUT31), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT31), .B1(new_n290), .B2(new_n310), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n309), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G472), .A2(G902), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT32), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT32), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n317), .A3(new_n314), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n306), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G217), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n320), .B1(G234), .B2(new_n304), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT22), .B(G137), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G125), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G140), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n327), .A2(new_n329), .A3(new_n330), .A4(KEYINPUT16), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT16), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT16), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(new_n326), .A3(G125), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT76), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n331), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G146), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n327), .A2(new_n329), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n208), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n219), .B1(new_n241), .B2(new_n243), .ZN(new_n342));
  NOR2_X1   g156(.A1(G119), .A2(G128), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT75), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(KEYINPUT24), .B(G110), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT75), .ZN(new_n346));
  INV_X1    g160(.A(new_n343), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT68), .B(G119), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n346), .B(new_n347), .C1(new_n348), .C2(new_n219), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n344), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n350), .A2(KEYINPUT77), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n344), .A2(new_n352), .A3(new_n345), .A4(new_n349), .ZN(new_n353));
  INV_X1    g167(.A(G110), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT23), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n348), .B2(G128), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n347), .B1(new_n348), .B2(new_n219), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n354), .B(new_n356), .C1(new_n357), .C2(new_n355), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n341), .B1(new_n351), .B2(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n208), .B(new_n331), .C1(new_n332), .C2(new_n335), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n337), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n356), .B1(new_n357), .B2(new_n355), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G110), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n344), .A2(new_n349), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n362), .B(new_n364), .C1(new_n345), .C2(new_n365), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n360), .A2(KEYINPUT78), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT78), .B1(new_n360), .B2(new_n366), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n325), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n360), .A2(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n324), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT25), .B1(new_n372), .B2(new_n304), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n374));
  AOI211_X1 g188(.A(new_n374), .B(G902), .C1(new_n369), .C2(new_n371), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n321), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n371), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT78), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n360), .A2(new_n366), .A3(KEYINPUT78), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n377), .B1(new_n381), .B2(new_n325), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n372), .A2(KEYINPUT79), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n321), .A2(G902), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n376), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n319), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT91), .ZN(new_n391));
  OR2_X1    g205(.A1(KEYINPUT72), .A2(G953), .ZN(new_n392));
  NAND2_X1  g206(.A1(KEYINPUT72), .A2(G953), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n392), .A2(G214), .A3(new_n192), .A4(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n210), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n191), .A2(G143), .A3(G214), .A4(new_n192), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G131), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT17), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(new_n396), .A3(new_n203), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n361), .ZN(new_n402));
  OAI211_X1 g216(.A(KEYINPUT76), .B(new_n334), .C1(new_n338), .C2(new_n333), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n208), .B1(new_n403), .B2(new_n331), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n203), .B1(new_n395), .B2(new_n396), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(KEYINPUT17), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n401), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n338), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT85), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n410), .A2(G146), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n340), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT86), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n395), .A2(new_n396), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(KEYINPUT18), .A2(G131), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n415), .A2(new_n416), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G113), .B(G122), .ZN(new_n420));
  INV_X1    g234(.A(G104), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n422), .B(KEYINPUT87), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n408), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n422), .B1(new_n408), .B2(new_n419), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n424), .B1(new_n425), .B2(KEYINPUT88), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT88), .ZN(new_n427));
  AOI211_X1 g241(.A(new_n427), .B(new_n422), .C1(new_n408), .C2(new_n419), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n304), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G475), .ZN(new_n430));
  NOR2_X1   g244(.A1(G475), .A2(G902), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n408), .A2(new_n419), .A3(new_n423), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT19), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n410), .B2(new_n411), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n339), .A2(KEYINPUT19), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n208), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n400), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n436), .B(new_n337), .C1(new_n437), .C2(new_n406), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n422), .B1(new_n419), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n431), .B1(new_n432), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT20), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n442), .B(new_n431), .C1(new_n432), .C2(new_n439), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n430), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(G478), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(KEYINPUT15), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n246), .A2(new_n248), .A3(KEYINPUT14), .A4(G122), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G107), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n246), .A2(new_n248), .A3(G122), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n245), .A2(G122), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT14), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n450), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n219), .A2(G143), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n219), .A2(G143), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n197), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n210), .A2(G128), .ZN(new_n461));
  OAI21_X1  g275(.A(G134), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G107), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n451), .A2(new_n464), .A3(new_n452), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT90), .B1(new_n456), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n460), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n453), .A2(G107), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n469), .B2(new_n465), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT13), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n471), .B1(new_n219), .B2(G143), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n210), .A2(KEYINPUT13), .A3(G128), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n459), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G134), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT89), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT89), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n474), .A2(new_n477), .A3(G134), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(G107), .B(new_n449), .C1(new_n453), .C2(KEYINPUT14), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n481), .A2(new_n482), .A3(new_n465), .A4(new_n463), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n467), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT9), .B(G234), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n485), .A2(new_n320), .A3(G953), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n467), .A2(new_n480), .A3(new_n483), .A4(new_n486), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n448), .B1(new_n490), .B2(new_n304), .ZN(new_n491));
  AOI211_X1 g305(.A(G902), .B(new_n447), .C1(new_n488), .C2(new_n489), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n445), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g309(.A(G221), .B1(new_n485), .B2(G902), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G469), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n191), .A2(G227), .ZN(new_n499));
  XOR2_X1   g313(.A(G110), .B(G140), .Z(new_n500));
  XOR2_X1   g314(.A(new_n499), .B(new_n500), .Z(new_n501));
  NAND2_X1  g315(.A1(new_n421), .A2(G107), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n421), .A2(G107), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT80), .ZN(new_n504));
  AOI21_X1  g318(.A(KEYINPUT3), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n504), .A2(new_n464), .A3(KEYINPUT3), .A4(G104), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n502), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT4), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(G101), .ZN(new_n510));
  INV_X1    g324(.A(G101), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n502), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n505), .B2(new_n507), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT4), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT3), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n464), .A2(G104), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n516), .B1(new_n517), .B2(KEYINPUT80), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n506), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n511), .B1(new_n519), .B2(new_n502), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n510), .B(new_n285), .C1(new_n515), .C2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n511), .B1(new_n517), .B2(new_n502), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n219), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n221), .B1(new_n524), .B2(new_n216), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n514), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT10), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n522), .B1(new_n519), .B2(new_n513), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n273), .A2(KEYINPUT10), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n521), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT81), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n521), .A2(KEYINPUT81), .A3(new_n528), .A4(new_n530), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n284), .A3(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n521), .A2(new_n207), .A3(new_n528), .A4(new_n530), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n501), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n536), .A2(new_n501), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n526), .B1(new_n273), .B2(new_n529), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n284), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT12), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT82), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n539), .A2(KEYINPUT12), .A3(new_n284), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n512), .B1(new_n518), .B2(new_n506), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n272), .B(new_n221), .C1(new_n546), .C2(new_n522), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n541), .B(new_n207), .C1(new_n547), .C2(new_n526), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT12), .B1(new_n539), .B2(new_n284), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT82), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n538), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n498), .B(new_n304), .C1(new_n537), .C2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n501), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n536), .B1(new_n548), .B2(new_n549), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n535), .A2(new_n538), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(G469), .B1(new_n555), .B2(G902), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n497), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n495), .A2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT84), .ZN(new_n559));
  XNOR2_X1  g373(.A(G110), .B(G122), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n560), .B(KEYINPUT8), .Z(new_n561));
  INV_X1    g375(.A(KEYINPUT5), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n348), .A2(new_n562), .A3(G116), .ZN(new_n563));
  OAI211_X1 g377(.A(G113), .B(new_n563), .C1(new_n250), .C2(new_n562), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n262), .B2(new_n263), .ZN(new_n565));
  INV_X1    g379(.A(new_n529), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n529), .B(new_n564), .C1(new_n262), .C2(new_n263), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n561), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n272), .A2(new_n328), .A3(new_n221), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n218), .A2(G125), .ZN(new_n571));
  INV_X1    g385(.A(G224), .ZN(new_n572));
  OR2_X1    g386(.A1(new_n572), .A2(G953), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n573), .A2(KEYINPUT7), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n570), .B(new_n571), .C1(KEYINPUT83), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(KEYINPUT83), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n576), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n570), .A2(new_n571), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n559), .B1(new_n569), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n561), .ZN(new_n582));
  INV_X1    g396(.A(new_n568), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n529), .B1(new_n294), .B2(new_n564), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n579), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n576), .B2(new_n575), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(KEYINPUT84), .A3(new_n587), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n292), .A2(new_n293), .B1(new_n258), .B2(new_n250), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n510), .B1(new_n515), .B2(new_n520), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n568), .B(new_n560), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n581), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n568), .B1(new_n589), .B2(new_n590), .ZN(new_n593));
  INV_X1    g407(.A(new_n560), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n595), .A2(KEYINPUT6), .A3(new_n591), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT6), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n593), .A2(new_n597), .A3(new_n594), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n570), .A2(new_n571), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n599), .B(new_n573), .Z(new_n600));
  NAND3_X1  g414(.A1(new_n596), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n592), .A2(new_n601), .A3(new_n304), .ZN(new_n602));
  OAI21_X1  g416(.A(G210), .B1(G237), .B2(G902), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n592), .A2(new_n601), .A3(new_n304), .A4(new_n603), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G952), .ZN(new_n608));
  AOI211_X1 g422(.A(G953), .B(new_n608), .C1(G234), .C2(G237), .ZN(new_n609));
  AOI211_X1 g423(.A(new_n304), .B(new_n191), .C1(G234), .C2(G237), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT21), .B(G898), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(G214), .B1(G237), .B2(G902), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n607), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n391), .B1(new_n558), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n614), .ZN(new_n617));
  AOI211_X1 g431(.A(new_n612), .B(new_n617), .C1(new_n605), .C2(new_n606), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n618), .A2(KEYINPUT91), .A3(new_n557), .A4(new_n495), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n390), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G101), .ZN(G3));
  INV_X1    g435(.A(new_n557), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n389), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n290), .A2(new_n310), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT31), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n290), .A2(new_n310), .A3(KEYINPUT31), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n626), .A2(new_n627), .B1(new_n308), .B2(new_n307), .ZN(new_n628));
  OAI21_X1  g442(.A(G472), .B1(new_n628), .B2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n315), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n615), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT92), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(KEYINPUT92), .A2(KEYINPUT33), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n481), .A2(new_n465), .A3(new_n463), .ZN(new_n637));
  AOI22_X1  g451(.A1(new_n637), .A2(KEYINPUT90), .B1(new_n470), .B2(new_n479), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n486), .B1(new_n638), .B2(new_n483), .ZN(new_n639));
  INV_X1    g453(.A(new_n489), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n635), .B(new_n636), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n488), .A2(new_n633), .A3(new_n634), .A4(new_n489), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n446), .A2(G902), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n490), .A2(new_n304), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n446), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n445), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n632), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT93), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT34), .B(G104), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  AOI22_X1  g467(.A1(G475), .A2(new_n429), .B1(new_n441), .B2(new_n443), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n494), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n632), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT35), .B(G107), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  INV_X1    g472(.A(KEYINPUT36), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n381), .A2(new_n659), .A3(new_n324), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n379), .B(new_n380), .C1(KEYINPUT36), .C2(new_n325), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n660), .A2(new_n387), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n374), .B1(new_n382), .B2(G902), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n372), .A2(KEYINPUT25), .A3(new_n304), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n662), .B1(new_n665), .B2(new_n321), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n630), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n616), .A2(new_n619), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT37), .B(G110), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT94), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n668), .B(new_n670), .ZN(G12));
  INV_X1    g485(.A(new_n662), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n376), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n557), .ZN(new_n674));
  INV_X1    g488(.A(new_n655), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n617), .B1(new_n605), .B2(new_n606), .ZN(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n610), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g492(.A1(new_n678), .A2(KEYINPUT95), .ZN(new_n679));
  INV_X1    g493(.A(new_n609), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(KEYINPUT95), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n675), .A2(new_n676), .A3(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n674), .A2(new_n319), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n219), .ZN(G30));
  AOI211_X1 g500(.A(new_n617), .B(new_n493), .C1(new_n430), .C2(new_n444), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n666), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT97), .Z(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT98), .B(KEYINPUT39), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n682), .B(new_n690), .Z(new_n691));
  NAND2_X1  g505(.A1(new_n557), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n692), .B(KEYINPUT40), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n607), .B(KEYINPUT38), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n316), .A2(new_n318), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n296), .A2(new_n308), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n299), .A2(new_n301), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n304), .B1(new_n698), .B2(new_n196), .ZN(new_n699));
  OAI21_X1  g513(.A(G472), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT96), .ZN(new_n702));
  OR3_X1    g516(.A1(new_n689), .A2(new_n695), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  NAND2_X1  g518(.A1(new_n607), .A2(new_n614), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n430), .A2(new_n444), .B1(new_n645), .B2(new_n647), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n683), .ZN(new_n707));
  OAI21_X1  g521(.A(KEYINPUT99), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n643), .A2(new_n644), .B1(new_n446), .B2(new_n646), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n654), .A2(new_n709), .A3(new_n682), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT99), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n676), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n674), .A2(new_n319), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(new_n208), .ZN(G48));
  NAND2_X1  g530(.A1(new_n297), .A2(new_n305), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G472), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n313), .A2(new_n317), .A3(new_n314), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n317), .B1(new_n313), .B2(new_n314), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n321), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n663), .B2(new_n664), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n384), .A2(new_n387), .A3(new_n385), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n721), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n538), .A2(new_n545), .A3(new_n550), .ZN(new_n727));
  INV_X1    g541(.A(new_n536), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n207), .B1(new_n531), .B2(new_n532), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n728), .B1(new_n729), .B2(new_n534), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n727), .B1(new_n730), .B2(new_n501), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n304), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(G469), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n496), .A3(new_n552), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT100), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n734), .A2(new_n735), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n726), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n618), .A3(new_n706), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND3_X1  g556(.A1(new_n739), .A2(new_n618), .A3(new_n675), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  NOR2_X1   g558(.A1(new_n705), .A2(new_n734), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n445), .A2(new_n612), .A3(new_n494), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n721), .A3(new_n673), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G119), .ZN(G21));
  NAND4_X1  g562(.A1(new_n676), .A2(new_n613), .A3(new_n494), .A4(new_n445), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n737), .A2(new_n749), .A3(new_n738), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n302), .A2(new_n266), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n308), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n752), .B1(new_n311), .B2(new_n312), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n753), .A2(KEYINPUT101), .A3(new_n314), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT101), .B1(new_n753), .B2(new_n314), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n629), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n389), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n750), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G122), .ZN(G24));
  NOR2_X1   g573(.A1(new_n756), .A2(new_n666), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(KEYINPUT102), .A3(new_n710), .A4(new_n745), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT102), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT101), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n196), .B1(new_n302), .B2(new_n266), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n626), .B2(new_n627), .ZN(new_n765));
  INV_X1    g579(.A(new_n314), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n753), .A2(KEYINPUT101), .A3(new_n314), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n673), .A2(new_n769), .A3(new_n629), .A4(new_n710), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n733), .A2(new_n552), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n676), .A3(new_n496), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n762), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n761), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G125), .ZN(G27));
  INV_X1    g590(.A(KEYINPUT104), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT103), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n552), .A2(new_n778), .A3(new_n556), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n778), .B1(new_n552), .B2(new_n556), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n605), .A2(new_n614), .A3(new_n606), .A4(new_n496), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n777), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n782), .A2(new_n779), .A3(new_n780), .A4(KEYINPUT104), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n390), .B(new_n710), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  XOR2_X1   g600(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT106), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n306), .B1(new_n696), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n316), .A2(KEYINPUT106), .A3(new_n318), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n389), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n710), .A2(KEYINPUT42), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n552), .A2(new_n556), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT103), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n552), .A2(new_n778), .A3(new_n556), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT104), .B1(new_n797), .B2(new_n782), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n781), .A2(new_n783), .A3(new_n777), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n793), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g614(.A1(new_n786), .A2(new_n788), .B1(new_n792), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(new_n203), .ZN(G33));
  NAND2_X1  g616(.A1(new_n798), .A2(new_n799), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n655), .A2(new_n682), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n390), .A3(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  NAND3_X1  g620(.A1(new_n605), .A2(new_n614), .A3(new_n606), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n445), .A2(new_n709), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT43), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n673), .A2(new_n630), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n807), .B1(new_n812), .B2(KEYINPUT44), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n555), .A2(KEYINPUT45), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n555), .A2(KEYINPUT45), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(G469), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(G469), .A2(G902), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT46), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(KEYINPUT46), .A3(new_n817), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n820), .A2(new_n552), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT107), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n822), .A2(new_n823), .A3(new_n496), .A4(new_n691), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(new_n496), .A3(new_n691), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT107), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT44), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n827), .B1(new_n810), .B2(new_n811), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n813), .A2(new_n824), .A3(new_n826), .A4(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G137), .ZN(G39));
  AND2_X1   g644(.A1(new_n822), .A2(new_n496), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n831), .A2(KEYINPUT47), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(KEYINPUT47), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n725), .A2(new_n707), .A3(new_n807), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n319), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G140), .ZN(G42));
  NAND2_X1  g651(.A1(new_n771), .A2(KEYINPUT49), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n614), .A3(new_n496), .A4(new_n808), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT49), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n840), .B2(new_n772), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n694), .A2(new_n389), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n702), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n783), .A2(new_n609), .A3(new_n772), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n389), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n702), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n846), .A2(KEYINPUT113), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(KEYINPUT113), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n654), .A3(new_n709), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n757), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n850), .A2(new_n680), .A3(new_n810), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n694), .A2(new_n614), .A3(new_n734), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT50), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n851), .A2(KEYINPUT50), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n810), .A2(new_n844), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n760), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT51), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n497), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n832), .A2(new_n833), .A3(new_n863), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n850), .A2(new_n810), .A3(new_n680), .A4(new_n807), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n849), .A2(new_n857), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT115), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n847), .A2(new_n706), .A3(new_n848), .ZN(new_n869));
  AOI211_X1 g683(.A(new_n608), .B(G953), .C1(new_n851), .C2(new_n745), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n792), .A2(new_n858), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(KEYINPUT48), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT116), .Z(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(KEYINPUT48), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT117), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n871), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n868), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT112), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n857), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n855), .A2(KEYINPUT112), .A3(new_n856), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n849), .A2(new_n880), .A3(new_n859), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n882), .A2(new_n883), .B1(new_n864), .B2(new_n865), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT51), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n685), .B1(new_n761), .B2(new_n774), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n687), .A2(new_n795), .A3(new_n607), .A4(new_n796), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n376), .A2(new_n672), .A3(new_n496), .A4(new_n683), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n714), .A2(new_n713), .B1(new_n890), .B2(new_n701), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n887), .A2(KEYINPUT52), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT52), .B1(new_n887), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT109), .ZN(new_n896));
  INV_X1    g710(.A(new_n770), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n803), .A2(new_n897), .ZN(new_n898));
  NOR4_X1   g712(.A1(new_n807), .A2(new_n494), .A3(new_n445), .A4(new_n682), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n714), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n805), .A2(new_n898), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n801), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n649), .A2(new_n655), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT108), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n706), .A2(KEYINPUT108), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n623), .A3(new_n631), .ZN(new_n907));
  INV_X1    g721(.A(new_n749), .ZN(new_n908));
  INV_X1    g722(.A(new_n738), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n909), .A3(new_n736), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n907), .B(new_n747), .C1(new_n850), .C2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n737), .A2(new_n738), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(new_n390), .A3(new_n618), .A4(new_n903), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n620), .A2(new_n668), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n896), .B1(new_n902), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n673), .A2(new_n746), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n773), .A2(new_n918), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n750), .A2(new_n757), .B1(new_n919), .B2(new_n721), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n619), .B(new_n616), .C1(new_n390), .C2(new_n667), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n920), .A2(new_n913), .A3(new_n907), .A4(new_n921), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n922), .A2(new_n801), .A3(new_n901), .A4(KEYINPUT109), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n895), .B1(new_n917), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT53), .ZN(new_n925));
  AOI22_X1  g739(.A1(new_n803), .A2(new_n897), .B1(new_n714), .B2(new_n899), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n726), .B1(new_n799), .B2(new_n798), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n787), .B1(new_n927), .B2(new_n710), .ZN(new_n928));
  INV_X1    g742(.A(new_n793), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n929), .B1(new_n784), .B2(new_n785), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n789), .B1(new_n719), .B2(new_n720), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n931), .A2(new_n791), .A3(new_n718), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n725), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n805), .B(new_n926), .C1(new_n928), .C2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT109), .B1(new_n935), .B2(new_n922), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n902), .A2(new_n916), .A3(new_n896), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT110), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n939), .B1(new_n892), .B2(new_n893), .ZN(new_n940));
  INV_X1    g754(.A(new_n685), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n775), .A2(new_n891), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT52), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n887), .A2(KEYINPUT52), .A3(new_n891), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n944), .A2(KEYINPUT110), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT53), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n938), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n925), .A2(KEYINPUT54), .A3(new_n949), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n935), .A2(new_n948), .A3(new_n922), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n892), .A2(new_n893), .A3(new_n939), .ZN(new_n952));
  AOI21_X1  g766(.A(KEYINPUT110), .B1(new_n944), .B2(new_n945), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT54), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n894), .B1(new_n936), .B2(new_n937), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n954), .B(new_n955), .C1(new_n956), .C2(KEYINPUT53), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n950), .A2(new_n957), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n878), .A2(new_n886), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(G952), .A2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n843), .B1(new_n959), .B2(new_n960), .ZN(G75));
  AOI22_X1  g775(.A1(new_n924), .A2(new_n948), .B1(new_n947), .B2(new_n951), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n304), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(G210), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT56), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n596), .A2(new_n598), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT118), .Z(new_n967));
  XNOR2_X1  g781(.A(new_n600), .B(KEYINPUT55), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n964), .A2(new_n965), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n964), .B2(new_n965), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n191), .A2(G952), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(G51));
  NOR3_X1   g787(.A1(new_n962), .A2(new_n304), .A3(new_n816), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT119), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n954), .B1(new_n956), .B2(KEYINPUT53), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT54), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n957), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n817), .B(KEYINPUT57), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n731), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n972), .B1(new_n975), .B2(new_n981), .ZN(G54));
  NAND3_X1  g796(.A1(new_n963), .A2(KEYINPUT58), .A3(G475), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n432), .A2(new_n439), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n985), .A2(new_n986), .A3(new_n972), .ZN(G60));
  NAND2_X1  g801(.A1(G478), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT59), .Z(new_n989));
  AOI21_X1  g803(.A(new_n989), .B1(new_n641), .B2(new_n642), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n924), .A2(new_n948), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n955), .B1(new_n991), .B2(new_n954), .ZN(new_n992));
  INV_X1    g806(.A(new_n957), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n990), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n972), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n989), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n643), .B1(new_n958), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(KEYINPUT120), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n972), .B1(new_n978), .B2(new_n990), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT120), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n989), .B1(new_n950), .B2(new_n957), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n1000), .B(new_n1001), .C1(new_n643), .C2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n999), .A2(new_n1003), .ZN(G63));
  NAND2_X1  g818(.A1(G217), .A2(G902), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT60), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n962), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1007), .A2(new_n660), .A3(new_n661), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n386), .B(KEYINPUT121), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1009), .B1(new_n962), .B2(new_n1006), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1008), .A2(new_n995), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT61), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1008), .A2(KEYINPUT61), .A3(new_n995), .A4(new_n1010), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(G66));
  OAI21_X1  g829(.A(G953), .B1(new_n611), .B2(new_n572), .ZN(new_n1016));
  INV_X1    g830(.A(new_n191), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1016), .B1(new_n916), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n967), .B1(G898), .B2(new_n191), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT122), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1018), .B(new_n1020), .ZN(G69));
  AOI21_X1  g835(.A(new_n191), .B1(G227), .B2(G900), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n836), .A2(new_n805), .A3(new_n829), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n687), .A2(new_n607), .ZN(new_n1024));
  AND4_X1   g838(.A1(new_n792), .A2(new_n826), .A3(new_n824), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n801), .ZN(new_n1027));
  INV_X1    g841(.A(new_n715), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n887), .A2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n1026), .A2(new_n191), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n281), .B1(new_n287), .B2(new_n289), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n434), .A2(new_n435), .ZN(new_n1032));
  XOR2_X1   g846(.A(new_n1031), .B(new_n1032), .Z(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(G900), .B2(new_n1017), .ZN(new_n1034));
  AND2_X1   g848(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1033), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n692), .A2(new_n807), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n390), .A2(new_n906), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n829), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1039), .A2(KEYINPUT123), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT123), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n829), .A2(new_n1041), .A3(new_n1038), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n703), .A2(new_n1029), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1044), .A2(KEYINPUT62), .ZN(new_n1045));
  INV_X1    g859(.A(KEYINPUT62), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n703), .A2(new_n1029), .A3(new_n1046), .ZN(new_n1047));
  NAND4_X1  g861(.A1(new_n1043), .A2(new_n836), .A3(new_n1045), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1036), .B1(new_n1048), .B2(new_n191), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1022), .B1(new_n1035), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1048), .A2(new_n191), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1051), .A2(new_n1033), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1052), .A2(KEYINPUT124), .ZN(new_n1053));
  INV_X1    g867(.A(KEYINPUT124), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g870(.A(new_n1022), .B(KEYINPUT125), .Z(new_n1057));
  AOI21_X1  g871(.A(new_n1057), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1058));
  AOI21_X1  g872(.A(KEYINPUT126), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g873(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1060));
  AOI211_X1 g874(.A(KEYINPUT124), .B(new_n1036), .C1(new_n1048), .C2(new_n191), .ZN(new_n1061));
  OAI211_X1 g875(.A(KEYINPUT126), .B(new_n1058), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g876(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g877(.A(new_n1050), .B1(new_n1059), .B2(new_n1063), .ZN(G72));
  NAND2_X1  g878(.A1(G472), .A2(G902), .ZN(new_n1065));
  XOR2_X1   g879(.A(new_n1065), .B(KEYINPUT63), .Z(new_n1066));
  NAND3_X1  g880(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1067));
  OAI21_X1  g881(.A(new_n1066), .B1(new_n1067), .B2(new_n922), .ZN(new_n1068));
  INV_X1    g882(.A(new_n296), .ZN(new_n1069));
  NOR2_X1   g883(.A1(new_n1069), .A2(new_n196), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n972), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g885(.A1(new_n1069), .A2(new_n308), .ZN(new_n1072));
  INV_X1    g886(.A(KEYINPUT127), .ZN(new_n1073));
  AOI22_X1  g887(.A1(new_n1072), .A2(new_n1073), .B1(new_n290), .B2(new_n310), .ZN(new_n1074));
  OAI21_X1  g888(.A(new_n1074), .B1(new_n1073), .B2(new_n1072), .ZN(new_n1075));
  NAND4_X1  g889(.A1(new_n925), .A2(new_n949), .A3(new_n1066), .A4(new_n1075), .ZN(new_n1076));
  OAI21_X1  g890(.A(new_n1066), .B1(new_n1048), .B2(new_n922), .ZN(new_n1077));
  NAND2_X1  g891(.A1(new_n1077), .A2(new_n697), .ZN(new_n1078));
  AND3_X1   g892(.A1(new_n1071), .A2(new_n1076), .A3(new_n1078), .ZN(G57));
endmodule


