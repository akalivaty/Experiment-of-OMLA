//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950;
  XOR2_X1   g000(.A(G78gat), .B(G106gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G22gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT31), .B(G50gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT76), .ZN(new_n207));
  XOR2_X1   g006(.A(G197gat), .B(G204gat), .Z(new_n208));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209));
  NAND2_X1  g008(.A1(G211gat), .A2(G218gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT70), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n210), .ZN(new_n214));
  NOR2_X1   g013(.A1(G211gat), .A2(G218gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n213), .B(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n207), .B1(new_n218), .B2(KEYINPUT29), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT29), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(KEYINPUT76), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT77), .ZN(new_n224));
  INV_X1    g023(.A(G141gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(G148gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G141gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n226), .A2(new_n228), .B1(KEYINPUT2), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n231), .A2(KEYINPUT72), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n229), .B1(new_n231), .B2(KEYINPUT72), .ZN(new_n233));
  OR3_X1    g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  OR2_X1    g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n229), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT73), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT73), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n238), .A3(new_n229), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n237), .A2(new_n230), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT74), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n234), .A2(KEYINPUT74), .A3(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n223), .A2(new_n224), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n224), .B1(new_n223), .B2(new_n245), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n221), .B1(new_n241), .B2(KEYINPUT3), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n218), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(G228gat), .A3(G233gat), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n246), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n221), .B1(new_n211), .B2(new_n216), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n252), .B1(new_n216), .B2(new_n211), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n241), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G228gat), .A2(G233gat), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n206), .B1(new_n251), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n257), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n247), .A2(new_n250), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n259), .B(new_n205), .C1(new_n260), .C2(new_n246), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(KEYINPUT65), .B(KEYINPUT28), .Z(new_n263));
  XOR2_X1   g062(.A(KEYINPUT27), .B(G183gat), .Z(new_n264));
  OAI21_X1  g063(.A(new_n263), .B1(new_n264), .B2(G190gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT27), .B(G183gat), .ZN(new_n267));
  INV_X1    g066(.A(G190gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(KEYINPUT65), .A2(KEYINPUT28), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n265), .A2(new_n266), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G169gat), .ZN(new_n273));
  INV_X1    g072(.A(G176gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT26), .ZN(new_n276));
  NOR2_X1   g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI211_X1 g077(.A(KEYINPUT66), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT66), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(new_n277), .B2(new_n276), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT23), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n277), .B(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n266), .A2(KEYINPUT24), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n285), .A2(new_n275), .ZN(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n268), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(KEYINPUT24), .A3(new_n266), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n284), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT25), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n284), .A2(new_n286), .A3(KEYINPUT25), .A4(new_n289), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n272), .A2(new_n282), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G113gat), .ZN(new_n295));
  INV_X1    g094(.A(G120gat), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT1), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n295), .B2(new_n296), .ZN(new_n298));
  XNOR2_X1  g097(.A(G127gat), .B(G134gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT67), .B(G113gat), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n297), .B(new_n299), .C1(new_n302), .C2(new_n296), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n294), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n292), .A2(new_n293), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n282), .A2(new_n266), .A3(new_n270), .A4(new_n265), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n304), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G227gat), .A2(G233gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n311), .B(KEYINPUT64), .Z(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n305), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT32), .ZN(new_n315));
  XOR2_X1   g114(.A(G15gat), .B(G43gat), .Z(new_n316));
  XNOR2_X1  g115(.A(G71gat), .B(G99gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT68), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT33), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n314), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n319), .B1(new_n314), .B2(new_n320), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n315), .B(new_n318), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(KEYINPUT33), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n314), .A2(KEYINPUT32), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(KEYINPUT69), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n310), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(new_n311), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT34), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT34), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(new_n330), .A3(new_n312), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n326), .B(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n262), .A2(new_n334), .ZN(new_n335));
  XOR2_X1   g134(.A(G1gat), .B(G29gat), .Z(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(G85gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT5), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n241), .A2(new_n304), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n342), .B(KEYINPUT4), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G225gat), .A2(G233gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n304), .B1(new_n241), .B2(KEYINPUT3), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT75), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n220), .B1(new_n243), .B2(new_n244), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n350), .A2(new_n351), .A3(new_n347), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n344), .B(new_n345), .C1(new_n349), .C2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n342), .B1(new_n245), .B2(new_n304), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n354), .A2(new_n345), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n341), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n346), .A2(KEYINPUT75), .A3(new_n348), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n351), .B1(new_n350), .B2(new_n347), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n343), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT5), .B1(new_n360), .B2(new_n345), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n340), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n353), .A2(new_n341), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n355), .B1(new_n360), .B2(new_n345), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n339), .B(new_n363), .C1(new_n364), .C2(new_n341), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n357), .A2(new_n361), .A3(new_n340), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT6), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT30), .ZN(new_n371));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G226gat), .A2(G233gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(new_n308), .B2(new_n221), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n294), .A2(new_n375), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n217), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n375), .B1(new_n294), .B2(KEYINPUT29), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n308), .A2(new_n376), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n380), .A2(new_n218), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n374), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT71), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  AOI211_X1 g184(.A(KEYINPUT71), .B(new_n374), .C1(new_n379), .C2(new_n382), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n371), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n379), .A2(new_n374), .A3(new_n382), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n388), .B1(KEYINPUT30), .B2(new_n383), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT35), .B1(new_n335), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n323), .A2(new_n333), .A3(new_n325), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n333), .B1(new_n323), .B2(new_n325), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n323), .A2(new_n325), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(new_n332), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(KEYINPUT81), .A3(new_n395), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n398), .A2(new_n401), .A3(new_n391), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n368), .A2(KEYINPUT80), .A3(KEYINPUT6), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT80), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n365), .B2(new_n366), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n367), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT35), .B1(new_n258), .B2(new_n261), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n334), .A2(KEYINPUT36), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT36), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n412), .B1(new_n396), .B2(new_n397), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n379), .A2(new_n382), .A3(KEYINPUT37), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n415), .A2(new_n374), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT38), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT79), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n379), .A2(new_n382), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT37), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  AOI211_X1 g220(.A(KEYINPUT79), .B(KEYINPUT37), .C1(new_n379), .C2(new_n382), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n416), .B(new_n417), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n423), .B1(new_n385), .B2(new_n386), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n421), .A2(new_n422), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n417), .B1(new_n425), .B2(new_n416), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n427), .A2(new_n406), .A3(new_n367), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n357), .A2(new_n361), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n339), .A2(new_n429), .B1(new_n387), .B2(new_n389), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT39), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n431), .B1(new_n354), .B2(new_n345), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n360), .B2(new_n345), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n360), .A2(KEYINPUT39), .A3(new_n345), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n434), .A2(KEYINPUT78), .A3(new_n339), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT78), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n344), .B1(new_n349), .B2(new_n352), .ZN(new_n437));
  INV_X1    g236(.A(new_n345), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n431), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n439), .B2(new_n340), .ZN(new_n440));
  OAI211_X1 g239(.A(KEYINPUT40), .B(new_n433), .C1(new_n435), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n430), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT78), .B1(new_n434), .B2(new_n339), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n436), .A3(new_n340), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT40), .B1(new_n445), .B2(new_n433), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n262), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n414), .B1(new_n428), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n390), .B1(new_n367), .B2(new_n369), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n449), .A2(new_n262), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n410), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT96), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT94), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT92), .ZN(new_n454));
  XOR2_X1   g253(.A(G99gat), .B(G106gat), .Z(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT8), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(G99gat), .B2(G106gat), .ZN(new_n459));
  NOR2_X1   g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(G99gat), .A2(G106gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT8), .ZN(new_n463));
  OR2_X1    g262(.A1(G85gat), .A2(G92gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT91), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(G85gat), .A2(G92gat), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT7), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n456), .B1(new_n466), .B2(new_n472), .ZN(new_n473));
  AOI211_X1 g272(.A(new_n455), .B(new_n471), .C1(new_n461), .C2(new_n465), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n454), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OR3_X1    g274(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n477));
  AOI22_X1  g276(.A1(new_n476), .A2(new_n477), .B1(G29gat), .B2(G36gat), .ZN(new_n478));
  INV_X1    g277(.A(G43gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT83), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT83), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G43gat), .ZN(new_n482));
  INV_X1    g281(.A(G50gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n480), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(KEYINPUT84), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT84), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G50gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n487), .A3(new_n479), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT15), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT15), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n479), .A2(new_n483), .ZN(new_n491));
  NAND2_X1  g290(.A1(G43gat), .A2(G50gat), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n478), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n477), .ZN(new_n495));
  NAND2_X1  g294(.A1(G29gat), .A2(G36gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n493), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n494), .A2(new_n499), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n463), .A2(KEYINPUT91), .A3(new_n464), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT91), .B1(new_n463), .B2(new_n464), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n472), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n455), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n456), .B(new_n472), .C1(new_n501), .C2(new_n502), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(KEYINPUT92), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n475), .A2(new_n500), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT17), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n511), .A3(new_n499), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n484), .A2(new_n488), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n493), .B1(new_n513), .B2(new_n490), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n499), .B1(new_n514), .B2(new_n497), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT17), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n504), .A2(KEYINPUT92), .A3(new_n505), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT92), .B1(new_n504), .B2(new_n505), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n512), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT93), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n494), .A2(new_n511), .A3(new_n499), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n511), .B1(new_n494), .B2(new_n499), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n475), .A2(new_n506), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT93), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n510), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(G190gat), .B(G218gat), .Z(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n519), .A2(new_n520), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n524), .A2(KEYINPUT93), .A3(new_n525), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(new_n528), .A3(new_n510), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n453), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT90), .ZN(new_n537));
  XNOR2_X1  g336(.A(G134gat), .B(G162gat), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n537), .B(new_n538), .Z(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n528), .B1(new_n533), .B2(new_n510), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(KEYINPUT94), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT95), .B1(new_n535), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n539), .B1(new_n530), .B2(new_n453), .ZN(new_n544));
  AOI211_X1 g343(.A(new_n529), .B(new_n509), .C1(new_n531), .C2(new_n532), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT94), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT95), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n540), .B1(new_n530), .B2(new_n534), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n452), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  AOI211_X1 g351(.A(KEYINPUT96), .B(new_n550), .C1(new_n543), .C2(new_n548), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT87), .ZN(new_n555));
  INV_X1    g354(.A(G8gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(G15gat), .B(G22gat), .ZN(new_n557));
  AND2_X1   g356(.A1(KEYINPUT85), .A2(G1gat), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT16), .B1(KEYINPUT85), .B2(G1gat), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n556), .B1(new_n560), .B2(KEYINPUT86), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n560), .B1(G1gat), .B2(new_n557), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI221_X1 g362(.A(new_n560), .B1(KEYINPUT86), .B2(new_n556), .C1(G1gat), .C2(new_n557), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n555), .B1(new_n566), .B2(new_n515), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n516), .A2(new_n512), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n567), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n524), .A2(new_n555), .A3(new_n566), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT18), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n569), .A2(KEYINPUT18), .A3(new_n570), .A4(new_n571), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n500), .B(new_n565), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n570), .B(KEYINPUT13), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n574), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G113gat), .B(G141gat), .ZN(new_n580));
  INV_X1    g379(.A(G197gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT11), .B(G169gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n586), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n574), .A2(new_n588), .A3(new_n575), .A4(new_n578), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G57gat), .B(G64gat), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  OAI22_X1  g393(.A1(new_n592), .A2(new_n593), .B1(KEYINPUT88), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G71gat), .B(G78gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n565), .B1(new_n598), .B2(KEYINPUT21), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n597), .B(KEYINPUT21), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(new_n600), .B2(new_n565), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n601), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT89), .ZN(new_n607));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n505), .A3(new_n504), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT10), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n597), .B1(new_n474), .B2(new_n473), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n475), .A2(KEYINPUT10), .A3(new_n506), .A4(new_n598), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n620), .B1(new_n614), .B2(new_n616), .ZN(new_n622));
  OR2_X1    g421(.A1(new_n622), .A2(KEYINPUT97), .ZN(new_n623));
  XNOR2_X1  g422(.A(G120gat), .B(G148gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(KEYINPUT97), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n621), .A2(new_n623), .A3(new_n627), .A4(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n620), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n630), .B1(new_n617), .B2(new_n618), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n626), .B1(new_n631), .B2(new_n622), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NOR4_X1   g432(.A1(new_n554), .A2(new_n591), .A3(new_n613), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n451), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n370), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g438(.A1(new_n635), .A2(new_n391), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT42), .B1(new_n640), .B2(new_n556), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT16), .B(G8gat), .Z(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  MUX2_X1   g442(.A(KEYINPUT42), .B(new_n641), .S(new_n643), .Z(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n635), .A2(new_n645), .A3(new_n414), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n398), .A2(new_n401), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n635), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n646), .B1(new_n645), .B2(new_n648), .ZN(G1326gat));
  NOR2_X1   g448(.A1(new_n635), .A2(new_n262), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT43), .B(G22gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  NOR3_X1   g451(.A1(new_n591), .A2(new_n612), .A3(new_n633), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n451), .A2(new_n554), .A3(new_n653), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n654), .A2(G29gat), .A3(new_n370), .ZN(new_n655));
  XOR2_X1   g454(.A(new_n655), .B(KEYINPUT45), .Z(new_n656));
  NAND3_X1  g455(.A1(new_n451), .A2(KEYINPUT44), .A3(new_n554), .ZN(new_n657));
  INV_X1    g456(.A(new_n262), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n392), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT98), .B1(new_n449), .B2(new_n262), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n410), .B1(new_n448), .B2(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n663), .A2(new_n554), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n657), .B(new_n653), .C1(new_n664), .C2(KEYINPUT44), .ZN(new_n665));
  OAI21_X1  g464(.A(G29gat), .B1(new_n665), .B2(new_n370), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n656), .A2(new_n666), .ZN(G1328gat));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n668));
  OR3_X1    g467(.A1(new_n665), .A2(new_n668), .A3(new_n391), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n665), .B2(new_n391), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(G36gat), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n391), .A2(G36gat), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n654), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(KEYINPUT99), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n654), .A2(new_n676), .A3(new_n673), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n675), .A2(KEYINPUT46), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(KEYINPUT46), .B1(new_n675), .B2(new_n677), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n679), .A2(new_n680), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n671), .B(new_n678), .C1(new_n681), .C2(new_n682), .ZN(G1329gat));
  AND2_X1   g482(.A1(new_n480), .A2(new_n482), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n665), .B2(new_n414), .ZN(new_n685));
  OR3_X1    g484(.A1(new_n654), .A2(new_n647), .A3(new_n684), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT47), .Z(G1330gat));
  AND2_X1   g487(.A1(new_n485), .A2(new_n487), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(new_n665), .B2(new_n262), .ZN(new_n690));
  OR3_X1    g489(.A1(new_n654), .A2(new_n262), .A3(new_n689), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT48), .Z(G1331gat));
  NAND2_X1  g492(.A1(new_n549), .A2(new_n551), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT96), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n549), .A2(new_n452), .A3(new_n551), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n697), .A2(new_n591), .A3(new_n612), .A4(new_n633), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n663), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n370), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT102), .B(G57gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1332gat));
  NOR2_X1   g502(.A1(new_n700), .A2(new_n391), .ZN(new_n704));
  NOR2_X1   g503(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n705));
  AND2_X1   g504(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(new_n704), .B2(new_n705), .ZN(G1333gat));
  NOR3_X1   g507(.A1(new_n700), .A2(G71gat), .A3(new_n647), .ZN(new_n709));
  INV_X1    g508(.A(new_n700), .ZN(new_n710));
  INV_X1    g509(.A(new_n414), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n709), .B1(G71gat), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n658), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g515(.A1(new_n590), .A2(new_n612), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n663), .A2(new_n554), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n663), .A2(KEYINPUT51), .A3(new_n554), .A4(new_n717), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  INV_X1    g524(.A(new_n633), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n370), .A2(G85gat), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n590), .A2(new_n612), .A3(new_n726), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n657), .B(new_n729), .C1(new_n664), .C2(KEYINPUT44), .ZN(new_n730));
  OAI21_X1  g529(.A(G85gat), .B1(new_n730), .B2(new_n370), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(G1336gat));
  NAND3_X1  g531(.A1(new_n720), .A2(KEYINPUT104), .A3(new_n721), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n734), .A3(new_n719), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n391), .A2(G92gat), .A3(new_n726), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n733), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT105), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n733), .A2(new_n739), .A3(new_n735), .A4(new_n736), .ZN(new_n740));
  OAI21_X1  g539(.A(G92gat), .B1(new_n730), .B2(new_n391), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT52), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT52), .ZN(new_n744));
  INV_X1    g543(.A(new_n736), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n741), .B(new_n744), .C1(new_n722), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(G1337gat));
  XOR2_X1   g546(.A(KEYINPUT106), .B(G99gat), .Z(new_n748));
  NOR3_X1   g547(.A1(new_n647), .A2(new_n726), .A3(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT107), .Z(new_n750));
  NAND3_X1  g549(.A1(new_n724), .A2(new_n725), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n748), .B1(new_n730), .B2(new_n414), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(G1338gat));
  OAI21_X1  g552(.A(G106gat), .B1(new_n730), .B2(new_n262), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n262), .A2(G106gat), .A3(new_n726), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(new_n754), .B(new_n755), .C1(new_n722), .C2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n733), .A2(new_n735), .A3(new_n756), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n760), .B2(new_n755), .ZN(G1339gat));
  NAND3_X1  g560(.A1(new_n617), .A2(new_n630), .A3(new_n618), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n621), .A2(KEYINPUT54), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n627), .B1(new_n631), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n763), .A2(KEYINPUT55), .A3(new_n765), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n629), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(KEYINPUT108), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n772));
  INV_X1    g571(.A(new_n629), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n766), .B2(new_n767), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n772), .B1(new_n774), .B2(new_n769), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n590), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n576), .A2(new_n577), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n584), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n589), .A2(new_n633), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n697), .A2(new_n781), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n771), .A2(new_n775), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n589), .A2(new_n779), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n783), .A2(new_n695), .A3(new_n696), .A4(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n612), .B1(new_n782), .B2(new_n785), .ZN(new_n786));
  NOR4_X1   g585(.A1(new_n554), .A2(new_n590), .A3(new_n613), .A4(new_n633), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n637), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n789), .A2(new_n262), .A3(new_n402), .ZN(new_n790));
  OAI21_X1  g589(.A(G113gat), .B1(new_n790), .B2(new_n591), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n335), .A2(new_n390), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n590), .A2(new_n302), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT109), .Z(new_n795));
  OAI21_X1  g594(.A(new_n791), .B1(new_n793), .B2(new_n795), .ZN(G1340gat));
  OAI21_X1  g595(.A(G120gat), .B1(new_n790), .B2(new_n726), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n633), .A2(new_n296), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT110), .ZN(G1341gat));
  INV_X1    g599(.A(new_n793), .ZN(new_n801));
  AOI21_X1  g600(.A(G127gat), .B1(new_n801), .B2(new_n612), .ZN(new_n802));
  INV_X1    g601(.A(G127gat), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n790), .A2(new_n803), .A3(new_n613), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n802), .A2(new_n804), .ZN(G1342gat));
  NOR2_X1   g604(.A1(new_n697), .A2(G134gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  OR3_X1    g606(.A1(new_n807), .A2(KEYINPUT111), .A3(KEYINPUT56), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT111), .B1(new_n807), .B2(KEYINPUT56), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(KEYINPUT56), .ZN(new_n810));
  OAI21_X1  g609(.A(G134gat), .B1(new_n790), .B2(new_n697), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(G1343gat));
  XNOR2_X1  g611(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n262), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n784), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n552), .A2(new_n553), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n784), .A2(new_n819), .A3(new_n633), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n780), .A2(KEYINPUT112), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n820), .B(new_n821), .C1(new_n591), .C2(new_n770), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n822), .B1(new_n552), .B2(new_n553), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n818), .A2(new_n783), .B1(new_n823), .B2(KEYINPUT113), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT113), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n822), .B(new_n825), .C1(new_n552), .C2(new_n553), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n612), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n814), .B(new_n816), .C1(new_n827), .C2(new_n787), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n823), .A2(KEYINPUT113), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n785), .A3(new_n826), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n787), .B1(new_n830), .B2(new_n613), .ZN(new_n831));
  INV_X1    g630(.A(new_n816), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT114), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n658), .B1(new_n786), .B2(new_n787), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n815), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n828), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n711), .A2(new_n370), .A3(new_n390), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n591), .A2(new_n225), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n788), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g640(.A(KEYINPUT115), .B(new_n637), .C1(new_n786), .C2(new_n787), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n711), .A2(new_n390), .A3(new_n262), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n841), .A2(new_n590), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n225), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n839), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n813), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n813), .ZN(new_n849));
  AOI211_X1 g648(.A(KEYINPUT116), .B(new_n849), .C1(new_n839), .C2(new_n845), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n848), .A2(new_n850), .ZN(G1344gat));
  AND2_X1   g650(.A1(new_n842), .A2(new_n843), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n852), .A2(new_n841), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n227), .A3(new_n633), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT118), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n853), .A2(new_n856), .A3(new_n227), .A4(new_n633), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n227), .A2(KEYINPUT59), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n836), .A2(new_n837), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(new_n726), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n834), .A2(KEYINPUT57), .ZN(new_n862));
  INV_X1    g661(.A(new_n770), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n554), .A2(new_n863), .A3(new_n784), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n823), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n612), .B1(new_n865), .B2(KEYINPUT119), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n864), .A2(new_n867), .A3(new_n823), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n787), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n658), .A2(new_n815), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n633), .B(new_n862), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n227), .B1(new_n872), .B2(new_n837), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n861), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n875), .ZN(G1345gat));
  NAND4_X1  g675(.A1(new_n841), .A2(new_n612), .A3(new_n842), .A4(new_n843), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT120), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n852), .A2(new_n879), .A3(new_n612), .A4(new_n841), .ZN(new_n880));
  INV_X1    g679(.A(G155gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n878), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n836), .A2(G155gat), .A3(new_n612), .A4(new_n837), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n882), .A2(KEYINPUT121), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1346gat));
  OAI21_X1  g687(.A(G162gat), .B1(new_n860), .B2(new_n697), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n697), .A2(G162gat), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n853), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n891), .A2(KEYINPUT122), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(KEYINPUT122), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(G1347gat));
  NOR2_X1   g693(.A1(new_n637), .A2(new_n391), .ZN(new_n895));
  XOR2_X1   g694(.A(new_n895), .B(KEYINPUT123), .Z(new_n896));
  NOR3_X1   g695(.A1(new_n896), .A2(new_n658), .A3(new_n647), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n786), .A2(new_n787), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n273), .B1(new_n899), .B2(new_n590), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT124), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n898), .A2(new_n895), .ZN(new_n902));
  INV_X1    g701(.A(new_n335), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n273), .A3(new_n590), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n901), .A2(new_n906), .ZN(G1348gat));
  NAND3_X1  g706(.A1(new_n899), .A2(G176gat), .A3(new_n633), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n274), .B1(new_n904), .B2(new_n726), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(KEYINPUT125), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(KEYINPUT125), .B2(new_n909), .ZN(G1349gat));
  NAND3_X1  g710(.A1(new_n905), .A2(new_n267), .A3(new_n612), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT60), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n899), .A2(new_n612), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n912), .B(new_n913), .C1(new_n287), .C2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n287), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n904), .A2(new_n264), .A3(new_n613), .ZN(new_n918));
  OAI21_X1  g717(.A(KEYINPUT60), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n916), .A2(new_n919), .ZN(G1350gat));
  AOI21_X1  g719(.A(new_n268), .B1(new_n899), .B2(new_n554), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT61), .Z(new_n922));
  NAND3_X1  g721(.A1(new_n905), .A2(new_n268), .A3(new_n554), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(G1351gat));
  NOR2_X1   g723(.A1(new_n896), .A2(new_n711), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n862), .B(new_n925), .C1(new_n869), .C2(new_n870), .ZN(new_n926));
  OAI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n591), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n711), .A2(new_n262), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n898), .A2(new_n928), .A3(new_n895), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n590), .A2(new_n581), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(G1352gat));
  OR2_X1    g730(.A1(new_n726), .A2(G204gat), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT62), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n929), .A2(KEYINPUT62), .A3(new_n932), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n936), .B1(new_n935), .B2(new_n934), .ZN(new_n937));
  INV_X1    g736(.A(new_n925), .ZN(new_n938));
  OAI21_X1  g737(.A(G204gat), .B1(new_n871), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n937), .A2(new_n939), .ZN(G1353gat));
  OR3_X1    g739(.A1(new_n929), .A2(G211gat), .A3(new_n613), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n926), .A2(new_n613), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n943));
  OAI211_X1 g742(.A(KEYINPUT63), .B(G211gat), .C1(new_n926), .C2(new_n613), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n941), .B1(new_n943), .B2(new_n945), .ZN(G1354gat));
  AOI21_X1  g745(.A(new_n697), .B1(new_n926), .B2(KEYINPUT127), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n947), .B1(KEYINPUT127), .B2(new_n926), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G218gat), .ZN(new_n949));
  OR3_X1    g748(.A1(new_n929), .A2(G218gat), .A3(new_n697), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1355gat));
endmodule


