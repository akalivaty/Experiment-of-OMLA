//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT0), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G143), .B(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(new_n195), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n199), .A3(G125), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n200), .A2(KEYINPUT84), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n193), .B1(new_n188), .B2(KEYINPUT1), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(new_n198), .ZN(new_n205));
  OR2_X1    g019(.A1(new_n205), .A2(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n200), .A2(KEYINPUT84), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n201), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G953), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G224), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n208), .B(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT78), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(G104), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  NOR3_X1   g032(.A1(new_n218), .A2(KEYINPUT78), .A3(G107), .ZN(new_n219));
  AOI21_X1  g033(.A(KEYINPUT3), .B1(new_n218), .B2(G107), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n213), .B(new_n217), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n216), .A2(G104), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n218), .A2(G107), .ZN(new_n223));
  OAI21_X1  g037(.A(G101), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT2), .A2(G113), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n230));
  INV_X1    g044(.A(G113), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n228), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G116), .B(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(KEYINPUT5), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n238), .A2(KEYINPUT5), .A3(G119), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(new_n231), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n226), .A2(new_n236), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT67), .B1(new_n234), .B2(new_n235), .ZN(new_n243));
  INV_X1    g057(.A(new_n233), .ZN(new_n244));
  NOR3_X1   g058(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n227), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n235), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n246), .A2(KEYINPUT67), .A3(new_n247), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n253), .A3(G101), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n221), .A2(KEYINPUT4), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n214), .A2(new_n216), .A3(G104), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n256), .B1(new_n222), .B2(KEYINPUT3), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n213), .B1(new_n257), .B2(new_n217), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n254), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n242), .B1(new_n251), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT82), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n242), .B(new_n262), .C1(new_n251), .C2(new_n259), .ZN(new_n263));
  XNOR2_X1  g077(.A(G110), .B(G122), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(KEYINPUT83), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n261), .A2(KEYINPUT6), .A3(new_n263), .A4(new_n265), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n242), .B(new_n264), .C1(new_n251), .C2(new_n259), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n265), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n269), .B1(new_n260), .B2(KEYINPUT82), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT6), .B1(new_n270), .B2(new_n263), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n212), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT7), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n208), .A2(new_n273), .A3(new_n211), .ZN(new_n274));
  XOR2_X1   g088(.A(new_n264), .B(KEYINPUT8), .Z(new_n275));
  AOI21_X1  g089(.A(KEYINPUT85), .B1(new_n235), .B2(KEYINPUT5), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n235), .A2(KEYINPUT85), .A3(KEYINPUT5), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n240), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n226), .B(new_n236), .C1(new_n276), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n241), .A2(new_n236), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n225), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n275), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n206), .A2(new_n200), .B1(KEYINPUT7), .B2(new_n210), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n274), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(G902), .B1(new_n284), .B2(new_n267), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n272), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(G210), .B1(G237), .B2(G902), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n272), .A2(new_n287), .A3(new_n285), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(KEYINPUT86), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G214), .B1(G237), .B2(G902), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT86), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n272), .A2(new_n293), .A3(new_n287), .A4(new_n285), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT30), .ZN(new_n296));
  INV_X1    g110(.A(G137), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(KEYINPUT11), .A3(G134), .ZN(new_n298));
  INV_X1    g112(.A(G134), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G137), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G131), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT11), .ZN(new_n303));
  OAI211_X1 g117(.A(KEYINPUT64), .B(new_n303), .C1(new_n299), .C2(G137), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n297), .A2(G134), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT64), .B1(new_n306), .B2(new_n303), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n301), .B(new_n302), .C1(new_n305), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n300), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G131), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n205), .A3(new_n310), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n197), .A2(new_n199), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n301), .B1(new_n305), .B2(new_n307), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G131), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n312), .B1(new_n314), .B2(new_n308), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n311), .B1(new_n315), .B2(KEYINPUT65), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n197), .A2(new_n199), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n298), .A2(new_n300), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n303), .B1(new_n299), .B2(G137), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT64), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI211_X1 g135(.A(G131), .B(new_n318), .C1(new_n321), .C2(new_n304), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n304), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n302), .B1(new_n323), .B2(new_n301), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n317), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT65), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n296), .B1(new_n316), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n251), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT68), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT69), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT1), .B1(new_n189), .B2(G146), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n333), .A2(G128), .B1(new_n188), .B2(new_n190), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n202), .A2(new_n188), .A3(new_n190), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n203), .B(KEYINPUT69), .C1(new_n204), .C2(new_n198), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n336), .A2(new_n337), .A3(new_n308), .A4(new_n310), .ZN(new_n338));
  OAI211_X1 g152(.A(KEYINPUT68), .B(new_n317), .C1(new_n322), .C2(new_n324), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n331), .A2(KEYINPUT30), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n328), .A2(new_n329), .A3(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n331), .A2(new_n251), .A3(new_n338), .A4(new_n339), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(G237), .A2(G953), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G210), .ZN(new_n345));
  XOR2_X1   g159(.A(new_n345), .B(KEYINPUT27), .Z(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT26), .B(G101), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n346), .B(new_n347), .Z(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n351));
  INV_X1    g165(.A(new_n342), .ZN(new_n352));
  AND3_X1   g166(.A1(new_n308), .A2(new_n205), .A3(new_n310), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n325), .B2(new_n326), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n315), .A2(KEYINPUT65), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n251), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT28), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n251), .A2(new_n338), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT28), .B1(new_n358), .B2(new_n325), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n348), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n350), .A2(new_n351), .A3(new_n361), .ZN(new_n362));
  XOR2_X1   g176(.A(KEYINPUT71), .B(G902), .Z(new_n363));
  NOR2_X1   g177(.A1(new_n349), .A2(new_n351), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT70), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n339), .A2(new_n338), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n314), .A2(new_n308), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT68), .B1(new_n367), .B2(new_n317), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n365), .B(new_n329), .C1(new_n366), .C2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n329), .B1(new_n366), .B2(new_n368), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n342), .A2(new_n365), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT28), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n360), .B(new_n364), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n362), .A2(new_n363), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G472), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n341), .A2(new_n348), .A3(new_n342), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(KEYINPUT31), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT31), .ZN(new_n380));
  NAND4_X1  g194(.A1(new_n341), .A2(new_n380), .A3(new_n348), .A4(new_n342), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n329), .B1(new_n316), .B2(new_n327), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n374), .B1(new_n382), .B2(new_n342), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n349), .B1(new_n383), .B2(new_n359), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n379), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT32), .ZN(new_n386));
  NOR2_X1   g200(.A1(G472), .A2(G902), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n386), .B1(new_n385), .B2(new_n387), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n377), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G140), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT16), .B1(new_n391), .B2(G125), .ZN(new_n392));
  INV_X1    g206(.A(G125), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n393), .A2(KEYINPUT73), .A3(G140), .ZN(new_n394));
  XNOR2_X1  g208(.A(G125), .B(G140), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n395), .B2(KEYINPUT73), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n392), .B1(new_n396), .B2(KEYINPUT16), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n187), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT73), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(new_n391), .A3(G125), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n391), .A2(G125), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n393), .A2(G140), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(KEYINPUT16), .B(new_n400), .C1(new_n403), .C2(new_n399), .ZN(new_n404));
  INV_X1    g218(.A(new_n392), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G146), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n398), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n193), .A2(G119), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT23), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n193), .A2(G119), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT72), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G110), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n409), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT24), .B(G110), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n408), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n418), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n421), .B1(new_n414), .B2(G110), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n395), .A2(new_n187), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n407), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT74), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n407), .A2(KEYINPUT74), .A3(new_n422), .A4(new_n423), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n420), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT75), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(KEYINPUT22), .B(G137), .Z(new_n431));
  AND3_X1   g245(.A1(new_n209), .A2(G221), .A3(G234), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n420), .A2(new_n426), .A3(KEYINPUT75), .A4(new_n427), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n430), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n428), .A2(new_n434), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT76), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(KEYINPUT25), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n436), .A2(new_n363), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G217), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n441), .B1(new_n363), .B2(G234), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n436), .A2(new_n363), .A3(new_n437), .ZN(new_n445));
  INV_X1    g259(.A(new_n439), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n442), .A2(G902), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n436), .A2(new_n449), .A3(new_n437), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G237), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n209), .A3(G214), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n189), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n344), .A2(G143), .A3(G214), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n302), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT17), .ZN(new_n457));
  INV_X1    g271(.A(new_n455), .ZN(new_n458));
  AOI21_X1  g272(.A(G143), .B1(new_n344), .B2(G214), .ZN(new_n459));
  OAI21_X1  g273(.A(G131), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT17), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n454), .A2(new_n302), .A3(new_n455), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n398), .A2(new_n407), .A3(new_n457), .A4(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G113), .B(G122), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(new_n218), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n396), .A2(G146), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n423), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n454), .A2(KEYINPUT88), .A3(new_n455), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT18), .A3(G131), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT18), .A2(G131), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n454), .A2(KEYINPUT88), .A3(new_n471), .A4(new_n455), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n464), .A2(new_n466), .A3(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n454), .A2(new_n302), .A3(new_n455), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n456), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n460), .A2(KEYINPUT89), .A3(new_n462), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(KEYINPUT19), .B(new_n400), .C1(new_n403), .C2(new_n399), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT19), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n395), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n187), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n397), .B2(new_n187), .ZN(new_n484));
  OAI211_X1 g298(.A(KEYINPUT90), .B(new_n473), .C1(new_n479), .C2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n466), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n407), .A2(new_n477), .A3(new_n483), .A4(new_n478), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT90), .B1(new_n488), .B2(new_n473), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n474), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT20), .ZN(new_n491));
  NOR2_X1   g305(.A1(G475), .A2(G902), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT91), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT91), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n490), .A2(new_n495), .A3(new_n491), .A4(new_n492), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n490), .A2(new_n492), .ZN(new_n497));
  XOR2_X1   g311(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n494), .A2(new_n496), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n474), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n466), .B1(new_n464), .B2(new_n473), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G475), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n189), .A2(G128), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n193), .A2(G143), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n507), .A2(new_n508), .A3(new_n299), .ZN(new_n509));
  INV_X1    g323(.A(G122), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G116), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n238), .A2(G122), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G107), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n511), .A2(new_n512), .A3(new_n216), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(new_n507), .ZN(new_n518));
  XOR2_X1   g332(.A(KEYINPUT92), .B(KEYINPUT13), .Z(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n508), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n518), .B1(new_n520), .B2(new_n507), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n509), .B(new_n516), .C1(new_n521), .C2(new_n299), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n507), .A2(new_n508), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G134), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n509), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT93), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n512), .A2(new_n526), .A3(KEYINPUT14), .ZN(new_n527));
  INV_X1    g341(.A(new_n512), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT14), .B1(new_n510), .B2(G116), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT93), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n512), .A2(KEYINPUT14), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n515), .B(new_n525), .C1(new_n532), .C2(new_n216), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT9), .B(G234), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n534), .A2(new_n441), .A3(G953), .ZN(new_n535));
  AND3_X1   g349(.A1(new_n522), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n535), .B1(new_n522), .B2(new_n533), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n363), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT94), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n540), .B(new_n363), .C1(new_n536), .C2(new_n537), .ZN(new_n541));
  INV_X1    g355(.A(G478), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n542), .A2(KEYINPUT15), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n539), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n538), .B(KEYINPUT94), .C1(KEYINPUT15), .C2(new_n542), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(G952), .ZN(new_n547));
  AOI211_X1 g361(.A(G953), .B(new_n547), .C1(G234), .C2(G237), .ZN(new_n548));
  AOI211_X1 g362(.A(new_n209), .B(new_n363), .C1(G234), .C2(G237), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT21), .B(G898), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n501), .A2(new_n506), .A3(new_n546), .A4(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G221), .ZN(new_n554));
  INV_X1    g368(.A(new_n534), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(new_n502), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT77), .ZN(new_n557));
  INV_X1    g371(.A(G469), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT80), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n336), .A2(new_n337), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n221), .A2(KEYINPUT10), .A3(new_n224), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n561), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n563), .A2(KEYINPUT80), .A3(new_n336), .A4(new_n337), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n333), .A2(KEYINPUT79), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT79), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n188), .A2(new_n567), .A3(KEYINPUT1), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n193), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n203), .B1(new_n569), .B2(new_n198), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(new_n226), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT10), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n252), .A2(G101), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n258), .A2(new_n253), .B1(new_n197), .B2(new_n199), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n571), .A2(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n367), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n565), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n205), .B1(new_n224), .B2(new_n221), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n226), .B2(new_n570), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT81), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n367), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT12), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n571), .B1(new_n205), .B2(new_n226), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT12), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n584), .A2(new_n581), .A3(new_n585), .A4(new_n367), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n578), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(G110), .B(G140), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n209), .A2(G227), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n565), .A2(new_n576), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n367), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n594), .A2(new_n578), .A3(new_n590), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n558), .B1(new_n596), .B2(new_n502), .ZN(new_n597));
  INV_X1    g411(.A(new_n363), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n565), .A2(new_n577), .A3(new_n576), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n577), .B1(new_n565), .B2(new_n576), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n591), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n578), .A2(new_n583), .A3(new_n586), .A4(new_n590), .ZN(new_n602));
  AOI211_X1 g416(.A(G469), .B(new_n598), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n557), .B1(new_n597), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n553), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n295), .A2(new_n390), .A3(new_n451), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(G101), .ZN(G3));
  NAND2_X1  g421(.A1(new_n385), .A2(new_n387), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n357), .A2(new_n360), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n349), .A2(new_n610), .B1(new_n378), .B2(KEYINPUT31), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n598), .B1(new_n611), .B2(new_n381), .ZN(new_n612));
  INV_X1    g426(.A(G472), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT95), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n385), .A2(new_n363), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT95), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(G472), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n609), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n448), .A2(new_n450), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n604), .ZN(new_n620));
  INV_X1    g434(.A(new_n292), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n289), .B2(new_n290), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(KEYINPUT33), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n623), .A2(KEYINPUT33), .ZN(new_n625));
  OR4_X1    g439(.A1(new_n536), .A2(new_n537), .A3(new_n624), .A4(new_n625), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n623), .B(KEYINPUT33), .C1(new_n536), .C2(new_n537), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n598), .A2(new_n542), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n628), .A2(new_n629), .B1(new_n542), .B2(new_n538), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n501), .B2(new_n506), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n551), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n618), .A2(new_n620), .A3(new_n622), .A4(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n634), .B(KEYINPUT97), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT34), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(new_n218), .ZN(G6));
  INV_X1    g451(.A(new_n492), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n488), .A2(new_n473), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT90), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n641), .A2(new_n486), .A3(new_n485), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n638), .B1(new_n642), .B2(new_n474), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT98), .B1(new_n643), .B2(new_n498), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n497), .A2(new_n645), .A3(new_n499), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n490), .A2(new_n492), .A3(new_n498), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT99), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n490), .A2(new_n649), .A3(new_n492), .A4(new_n498), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n644), .A2(new_n646), .A3(new_n648), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n464), .A2(new_n473), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n486), .ZN(new_n653));
  AOI21_X1  g467(.A(G902), .B1(new_n653), .B2(new_n474), .ZN(new_n654));
  INV_X1    g468(.A(G475), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT100), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n505), .A2(new_n657), .A3(G475), .ZN(new_n658));
  AND4_X1   g472(.A1(new_n545), .A2(new_n656), .A3(new_n544), .A4(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n651), .A2(new_n659), .A3(new_n552), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(KEYINPUT101), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n651), .A2(new_n659), .A3(new_n662), .A4(new_n552), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n618), .A2(new_n620), .A3(new_n622), .A4(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT35), .B(G107), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G9));
  NOR2_X1   g481(.A1(new_n434), .A2(KEYINPUT36), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n430), .B2(new_n435), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n430), .A2(new_n435), .A3(new_n669), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n449), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n447), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n673), .B1(new_n674), .B2(new_n443), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n618), .A2(new_n295), .A3(new_n605), .A4(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n548), .B1(new_n549), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n651), .A2(new_n659), .A3(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n604), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n390), .A2(new_n683), .A3(new_n622), .A4(new_n675), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  NAND2_X1  g499(.A1(new_n291), .A2(new_n294), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(KEYINPUT38), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT38), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n291), .A2(new_n688), .A3(new_n294), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n601), .A2(new_n602), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(new_n558), .A3(new_n363), .ZN(new_n693));
  AOI21_X1  g507(.A(G902), .B1(new_n592), .B2(new_n595), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n693), .B1(new_n558), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n680), .B(KEYINPUT39), .Z(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n557), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT40), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n675), .A2(new_n621), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT40), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n695), .A2(new_n700), .A3(new_n557), .A4(new_n696), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n546), .B1(new_n501), .B2(new_n506), .ZN(new_n702));
  AND4_X1   g516(.A1(new_n698), .A2(new_n699), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n378), .B1(new_n373), .B2(new_n348), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n502), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(G472), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n388), .B2(new_n389), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n691), .A2(new_n703), .A3(new_n704), .A4(new_n708), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n701), .A2(new_n702), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(new_n708), .A3(new_n698), .A4(new_n699), .ZN(new_n711));
  OAI21_X1  g525(.A(KEYINPUT102), .B1(new_n711), .B2(new_n690), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G143), .ZN(G45));
  NAND2_X1  g528(.A1(new_n631), .A2(new_n681), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n604), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(new_n390), .A3(new_n622), .A4(new_n675), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G146), .ZN(G48));
  NAND2_X1  g532(.A1(new_n692), .A2(new_n363), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(G469), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT103), .B1(new_n721), .B2(new_n558), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n721), .A2(new_n724), .A3(new_n558), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n556), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n727), .A2(new_n728), .A3(new_n622), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n729), .A2(new_n451), .A3(new_n390), .A4(new_n633), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND4_X1  g546(.A1(new_n729), .A2(new_n664), .A3(new_n451), .A4(new_n390), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  AND3_X1   g548(.A1(new_n671), .A2(new_n449), .A3(new_n672), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n444), .B2(new_n447), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n553), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n556), .B1(new_n723), .B2(new_n726), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n390), .A2(new_n737), .A3(new_n622), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G119), .ZN(G21));
  NAND3_X1  g554(.A1(new_n727), .A2(new_n728), .A3(new_n552), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n622), .A2(new_n702), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n612), .A2(new_n613), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n372), .A2(new_n371), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n374), .B1(new_n745), .B2(new_n369), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n349), .B1(new_n746), .B2(new_n359), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n379), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT104), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n369), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n359), .B1(new_n751), .B2(KEYINPUT28), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n750), .B(new_n379), .C1(new_n752), .C2(new_n348), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n749), .A2(new_n381), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n744), .B1(new_n754), .B2(new_n387), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n743), .A2(new_n755), .A3(KEYINPUT105), .A4(new_n451), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT105), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n753), .A2(new_n381), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n750), .B1(new_n747), .B2(new_n379), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n387), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n744), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n761), .A3(new_n451), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n738), .A2(new_n552), .A3(new_n622), .A4(new_n702), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n756), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G122), .ZN(G24));
  NAND3_X1  g580(.A1(new_n760), .A2(new_n761), .A3(new_n675), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n680), .B(new_n630), .C1(new_n501), .C2(new_n506), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n738), .A2(new_n622), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n393), .ZN(G27));
  NAND2_X1  g585(.A1(new_n390), .A2(new_n451), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n686), .A2(new_n292), .A3(new_n695), .A4(new_n728), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT42), .B1(new_n774), .B2(new_n768), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT42), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n772), .A2(new_n773), .A3(new_n776), .A4(new_n715), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n302), .ZN(G33));
  NAND2_X1  g593(.A1(new_n608), .A2(KEYINPUT32), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n619), .B1(new_n782), .B2(new_n377), .ZN(new_n783));
  INV_X1    g597(.A(new_n682), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n621), .B(new_n556), .C1(new_n291), .C2(new_n294), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n695), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  NOR2_X1   g601(.A1(new_n618), .A2(new_n736), .ZN(new_n788));
  INV_X1    g602(.A(new_n630), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n501), .A2(KEYINPUT107), .A3(new_n506), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT107), .B1(new_n501), .B2(new_n506), .ZN(new_n791));
  OAI211_X1 g605(.A(KEYINPUT43), .B(new_n789), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n501), .A2(new_n506), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n630), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n792), .B1(KEYINPUT43), .B2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n788), .A2(KEYINPUT44), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT108), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n788), .A2(new_n798), .A3(KEYINPUT44), .A4(new_n795), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT44), .B1(new_n788), .B2(new_n795), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n621), .B1(new_n291), .B2(new_n294), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n592), .A2(new_n804), .A3(new_n595), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n804), .B1(new_n592), .B2(new_n595), .ZN(new_n806));
  OAI21_X1  g620(.A(G469), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(G469), .A2(G902), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(KEYINPUT46), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT106), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT106), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n807), .A2(new_n811), .A3(KEYINPUT46), .A4(new_n808), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT46), .ZN(new_n813));
  INV_X1    g627(.A(new_n806), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n592), .A2(new_n804), .A3(new_n595), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n813), .B(G469), .C1(new_n816), .C2(G902), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n810), .A2(new_n693), .A3(new_n812), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n728), .A3(new_n696), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n801), .A2(new_n803), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n800), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(KEYINPUT109), .B(G137), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(G39));
  NOR4_X1   g637(.A1(new_n803), .A2(new_n390), .A3(new_n451), .A4(new_n715), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n817), .A2(new_n812), .A3(new_n693), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n809), .A2(KEYINPUT106), .ZN(new_n826));
  OAI211_X1 g640(.A(KEYINPUT47), .B(new_n728), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT47), .B1(new_n818), .B2(new_n728), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n824), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G140), .ZN(G42));
  AND2_X1   g645(.A1(new_n795), .A2(new_n548), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n762), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n690), .A2(new_n621), .A3(new_n738), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT50), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n785), .A2(new_n727), .ZN(new_n843));
  INV_X1    g657(.A(new_n708), .ZN(new_n844));
  AND4_X1   g658(.A1(new_n451), .A2(new_n843), .A3(new_n548), .A4(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n506), .A3(new_n501), .A4(new_n630), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT116), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n834), .A2(new_n675), .A3(new_n755), .A4(new_n843), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n834), .A2(new_n835), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n828), .A2(new_n829), .ZN(new_n850));
  INV_X1    g664(.A(new_n727), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n850), .B1(new_n557), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n802), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n855));
  OR3_X1    g669(.A1(new_n842), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n855), .B1(new_n842), .B2(new_n854), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n834), .A2(new_n783), .A3(new_n843), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT48), .ZN(new_n859));
  INV_X1    g673(.A(new_n729), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT117), .B1(new_n849), .B2(new_n860), .ZN(new_n861));
  OR3_X1    g675(.A1(new_n849), .A2(KEYINPUT117), .A3(new_n860), .ZN(new_n862));
  AOI211_X1 g676(.A(new_n547), .B(G953), .C1(new_n845), .C2(new_n631), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n859), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n856), .A2(new_n857), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n546), .A2(new_n656), .A3(new_n658), .A4(new_n681), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(new_n695), .A3(new_n651), .A4(new_n557), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(new_n736), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n390), .A3(new_n802), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n760), .A2(new_n761), .A3(new_n675), .A4(new_n768), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n786), .B(new_n870), .C1(new_n773), .C2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n775), .ZN(new_n873));
  INV_X1    g687(.A(new_n777), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n606), .A2(new_n739), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n501), .A2(new_n506), .A3(new_n545), .A4(new_n544), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n551), .B1(new_n632), .B2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n618), .A2(new_n295), .A3(new_n620), .A4(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n783), .B(new_n729), .C1(new_n633), .C2(new_n664), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n876), .A2(new_n676), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n756), .A2(new_n764), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT110), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n875), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n869), .A2(new_n390), .A3(new_n802), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n774), .B2(new_n784), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n871), .A2(new_n773), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n887), .B(new_n888), .C1(new_n775), .C2(new_n777), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n879), .A2(new_n730), .A3(new_n733), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n606), .A2(new_n739), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n272), .A2(new_n287), .A3(new_n285), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n287), .B1(new_n272), .B2(new_n285), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n293), .ZN(new_n894));
  INV_X1    g708(.A(new_n294), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(new_n292), .A3(new_n605), .A4(new_n675), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n616), .B1(new_n615), .B2(G472), .ZN(new_n898));
  AOI211_X1 g712(.A(KEYINPUT95), .B(new_n613), .C1(new_n385), .C2(new_n363), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n608), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n891), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n890), .A2(new_n765), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT110), .B1(new_n889), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n885), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n597), .A2(new_n603), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n680), .B(KEYINPUT113), .Z(new_n907));
  NOR4_X1   g721(.A1(new_n675), .A2(new_n906), .A3(new_n556), .A4(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n908), .A2(new_n622), .A3(new_n708), .A4(new_n702), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n909), .A2(new_n717), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n684), .B1(new_n767), .B2(new_n769), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT52), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n910), .A2(new_n912), .A3(KEYINPUT52), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n866), .B1(new_n905), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n717), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n909), .A2(KEYINPUT52), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n911), .A2(KEYINPUT112), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT112), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n684), .B(new_n921), .C1(new_n767), .C2(new_n769), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n918), .B(new_n919), .C1(new_n920), .C2(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT114), .B1(new_n923), .B2(new_n913), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n920), .A2(new_n922), .ZN(new_n925));
  INV_X1    g739(.A(new_n919), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n925), .A2(new_n717), .A3(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT114), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n927), .A2(new_n914), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT111), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n885), .A2(new_n904), .A3(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT53), .B1(new_n905), .B2(KEYINPUT111), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n917), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT54), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT53), .B1(new_n905), .B2(new_n916), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n875), .A2(new_n883), .A3(KEYINPUT53), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n924), .B2(new_n929), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n936), .A2(new_n942), .ZN(new_n943));
  OAI22_X1  g757(.A1(new_n865), .A2(new_n943), .B1(G952), .B2(G953), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n727), .B(KEYINPUT49), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n945), .A2(new_n451), .A3(new_n292), .A4(new_n557), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n947));
  OR3_X1    g761(.A1(new_n946), .A2(new_n708), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n944), .B1(new_n691), .B2(new_n948), .ZN(G75));
  NOR2_X1   g763(.A1(new_n268), .A2(new_n271), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT118), .Z(new_n951));
  XOR2_X1   g765(.A(new_n212), .B(KEYINPUT55), .Z(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n598), .B(new_n288), .C1(new_n937), .C2(new_n939), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n956), .B2(KEYINPUT56), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT56), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n955), .A2(new_n958), .A3(new_n953), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n209), .A2(G952), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n957), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT119), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT119), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n957), .A2(new_n964), .A3(new_n959), .A4(new_n961), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n963), .A2(new_n965), .ZN(G51));
  XOR2_X1   g780(.A(new_n808), .B(KEYINPUT57), .Z(new_n967));
  INV_X1    g781(.A(new_n942), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n940), .A2(new_n941), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n692), .ZN(new_n971));
  INV_X1    g785(.A(new_n940), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n598), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n973), .A2(new_n807), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n960), .B1(new_n971), .B2(new_n974), .ZN(G54));
  INV_X1    g789(.A(new_n490), .ZN(new_n976));
  NAND2_X1  g790(.A1(KEYINPUT58), .A2(G475), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n976), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n961), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n973), .A2(new_n976), .A3(new_n977), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n979), .A2(new_n980), .ZN(G60));
  NAND2_X1  g795(.A1(G478), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT59), .Z(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n628), .B(new_n984), .C1(new_n968), .C2(new_n969), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n961), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n628), .B1(new_n943), .B2(new_n984), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n986), .A2(new_n987), .ZN(G63));
  NAND2_X1  g802(.A1(G217), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT60), .Z(new_n990));
  NAND4_X1  g804(.A1(new_n972), .A2(new_n671), .A3(new_n672), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n436), .A2(new_n437), .ZN(new_n992));
  INV_X1    g806(.A(new_n990), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n992), .B1(new_n940), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n991), .A2(new_n961), .A3(new_n994), .ZN(new_n995));
  XOR2_X1   g809(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(G66));
  NAND2_X1  g811(.A1(G224), .A2(G953), .ZN(new_n998));
  OAI22_X1  g812(.A1(new_n903), .A2(G953), .B1(new_n550), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(G898), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n951), .B1(new_n1000), .B2(G953), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n999), .B(new_n1001), .ZN(G69));
  AOI21_X1  g816(.A(new_n209), .B1(G227), .B2(G900), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n328), .A2(new_n340), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT121), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n480), .A2(new_n482), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1007), .B1(G900), .B2(G953), .ZN(new_n1008));
  OR3_X1    g822(.A1(new_n819), .A2(new_n772), .A3(new_n742), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1009), .A2(new_n830), .A3(new_n786), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1010), .A2(new_n778), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT123), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n918), .B1(new_n920), .B2(new_n922), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n821), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1012), .B1(new_n821), .B2(new_n1013), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1008), .B1(new_n1016), .B2(G953), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1003), .B1(new_n1017), .B2(KEYINPUT122), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n1013), .A2(KEYINPUT62), .A3(new_n713), .ZN(new_n1019));
  AOI21_X1  g833(.A(KEYINPUT62), .B1(new_n1013), .B2(new_n713), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n697), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n632), .A2(new_n877), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n783), .A2(new_n1022), .A3(new_n802), .A4(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n830), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1025), .B1(new_n800), .B2(new_n820), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n209), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n1007), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1017), .A2(new_n1029), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1018), .B(new_n1030), .Z(G72));
  INV_X1    g845(.A(KEYINPUT127), .ZN(new_n1032));
  NAND2_X1  g846(.A1(G472), .A2(G902), .ZN(new_n1033));
  XOR2_X1   g847(.A(new_n1033), .B(KEYINPUT63), .Z(new_n1034));
  OAI21_X1  g848(.A(new_n1034), .B1(new_n1016), .B2(new_n903), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n343), .A2(new_n348), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n960), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT126), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1034), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1039), .B1(new_n350), .B2(new_n378), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1038), .B1(new_n935), .B2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n884), .B1(new_n875), .B2(new_n883), .ZN(new_n1042));
  NOR3_X1   g856(.A1(new_n889), .A2(new_n903), .A3(KEYINPUT110), .ZN(new_n1043));
  OAI21_X1  g857(.A(KEYINPUT111), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g858(.A1(new_n1044), .A2(new_n866), .A3(new_n932), .A4(new_n930), .ZN(new_n1045));
  INV_X1    g859(.A(new_n917), .ZN(new_n1046));
  AND4_X1   g860(.A1(new_n1038), .A2(new_n1045), .A3(new_n1046), .A4(new_n1040), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1037), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n343), .A2(new_n348), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n1026), .B(new_n883), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1050), .A2(new_n1034), .ZN(new_n1051));
  INV_X1    g865(.A(KEYINPUT124), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g867(.A(KEYINPUT125), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n1050), .A2(KEYINPUT124), .A3(new_n1034), .ZN(new_n1055));
  AND3_X1   g869(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1054), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1032), .B1(new_n1048), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1060), .A2(KEYINPUT125), .ZN(new_n1061));
  NAND3_X1  g875(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n935), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1064));
  NAND3_X1  g878(.A1(new_n1045), .A2(new_n1046), .A3(new_n1040), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1065), .A2(KEYINPUT126), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g881(.A1(new_n1063), .A2(new_n1067), .A3(KEYINPUT127), .A4(new_n1037), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1059), .A2(new_n1068), .ZN(G57));
endmodule


