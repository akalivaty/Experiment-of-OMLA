//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT72), .ZN(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(KEYINPUT27), .B(G183gat), .Z(new_n207));
  INV_X1    g006(.A(KEYINPUT28), .ZN(new_n208));
  NOR3_X1   g007(.A1(new_n207), .A2(new_n208), .A3(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT27), .ZN(new_n212));
  OR2_X1    g011(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n211), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT68), .B1(new_n217), .B2(new_n208), .ZN(new_n218));
  AND2_X1   g017(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT27), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n216), .ZN(new_n222));
  AOI21_X1  g021(.A(G190gat), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT28), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n210), .B1(new_n218), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n229), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n227), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n226), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n228), .A2(KEYINPUT23), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(G169gat), .B2(G176gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n237), .A2(new_n239), .A3(KEYINPUT25), .A4(new_n230), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n213), .A2(new_n211), .A3(new_n214), .ZN(new_n241));
  NAND3_X1  g040(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT24), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n227), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n244), .B1(new_n227), .B2(new_n245), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n240), .B1(new_n243), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n237), .A2(new_n230), .A3(new_n239), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n227), .A2(new_n245), .ZN(new_n252));
  INV_X1    g051(.A(G183gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(new_n211), .A3(KEYINPUT64), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(G183gat), .B2(G190gat), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n252), .A2(new_n254), .A3(new_n256), .A4(new_n242), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT25), .B1(new_n251), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT67), .B1(new_n249), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT25), .ZN(new_n260));
  INV_X1    g059(.A(new_n257), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(new_n250), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n241), .B(new_n242), .C1(new_n246), .C2(new_n247), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n251), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT67), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  XOR2_X1   g066(.A(G113gat), .B(G120gat), .Z(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G134gat), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G113gat), .B(G120gat), .ZN(new_n272));
  INV_X1    g071(.A(G127gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(G134gat), .ZN(new_n274));
  INV_X1    g073(.A(G134gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(G127gat), .ZN(new_n276));
  OAI22_X1  g075(.A1(new_n272), .A2(KEYINPUT1), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g076(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n236), .A2(new_n267), .A3(KEYINPUT69), .A4(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n249), .A2(new_n258), .A3(KEYINPUT67), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n265), .B1(new_n262), .B2(new_n264), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n224), .B1(new_n223), .B2(KEYINPUT28), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT66), .B(G183gat), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n216), .B1(new_n284), .B2(KEYINPUT27), .ZN(new_n285));
  OAI211_X1 g084(.A(KEYINPUT68), .B(new_n208), .C1(new_n285), .C2(G190gat), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n209), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  OAI22_X1  g086(.A1(new_n281), .A2(new_n282), .B1(new_n287), .B2(new_n234), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n271), .A2(new_n277), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n280), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n288), .A2(new_n289), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n279), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G227gat), .A2(G233gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n206), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n236), .A2(new_n278), .A3(new_n267), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n278), .B1(new_n236), .B2(new_n267), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n300), .B2(new_n280), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n293), .B1(new_n301), .B2(new_n279), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT32), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n298), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n295), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n297), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT34), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n307), .A2(KEYINPUT74), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n279), .B(new_n308), .C1(new_n290), .C2(new_n291), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n311), .B1(new_n301), .B2(new_n279), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n293), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n307), .A2(KEYINPUT73), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n301), .A2(new_n279), .A3(new_n293), .ZN(new_n315));
  AND2_X1   g114(.A1(new_n307), .A2(KEYINPUT73), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n295), .B(KEYINPUT32), .C1(new_n206), .C2(new_n296), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n306), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT76), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n306), .A2(new_n318), .A3(new_n319), .A4(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n319), .ZN(new_n325));
  INV_X1    g124(.A(new_n296), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n205), .B1(new_n302), .B2(new_n326), .ZN(new_n327));
  AOI211_X1 g126(.A(new_n298), .B(new_n303), .C1(new_n292), .C2(new_n294), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n325), .B1(new_n329), .B2(new_n304), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT75), .B1(new_n330), .B2(new_n318), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n318), .B1(new_n306), .B2(new_n319), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n324), .A2(KEYINPUT36), .A3(new_n331), .A4(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n332), .B1(new_n321), .B2(new_n323), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(KEYINPUT36), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G78gat), .B(G106gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT31), .B(G50gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT22), .ZN(new_n342));
  INV_X1    g141(.A(G211gat), .ZN(new_n343));
  INV_X1    g142(.A(G218gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G204gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(G197gat), .ZN(new_n347));
  INV_X1    g146(.A(G197gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G204gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G211gat), .B(G218gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(KEYINPUT78), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT78), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n352), .B(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(KEYINPUT77), .A3(new_n350), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n341), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n355), .A2(new_n358), .A3(new_n341), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT84), .ZN(new_n363));
  NAND2_X1  g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT2), .ZN(new_n365));
  OR2_X1    g164(.A1(G141gat), .A2(G148gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(G141gat), .A2(G148gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n364), .ZN(new_n369));
  NOR2_X1   g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n363), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n367), .ZN(new_n373));
  NOR2_X1   g172(.A1(G141gat), .A2(G148gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G155gat), .B(G162gat), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n375), .A2(new_n376), .A3(KEYINPUT84), .A4(new_n365), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n372), .A2(new_n377), .B1(new_n371), .B2(new_n368), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n360), .A2(new_n361), .B1(new_n362), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n355), .A2(new_n358), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n362), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n378), .B1(new_n383), .B2(new_n379), .ZN(new_n384));
  INV_X1    g183(.A(G228gat), .ZN(new_n385));
  INV_X1    g184(.A(G233gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n381), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n361), .ZN(new_n390));
  INV_X1    g189(.A(new_n380), .ZN(new_n391));
  OAI22_X1  g190(.A1(new_n390), .A2(new_n359), .B1(KEYINPUT29), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n357), .A2(new_n350), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n353), .A2(new_n351), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n362), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n379), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n372), .A2(new_n377), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n368), .A2(new_n371), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n387), .B1(new_n392), .B2(new_n400), .ZN(new_n401));
  OR3_X1    g200(.A1(new_n389), .A2(new_n401), .A3(G22gat), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n340), .B1(new_n402), .B2(KEYINPUT88), .ZN(new_n403));
  OAI21_X1  g202(.A(G22gat), .B1(new_n389), .B2(new_n401), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n403), .B(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(G226gat), .A2(G233gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n249), .A2(new_n258), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n408), .B1(new_n226), .B2(new_n235), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n407), .B1(new_n409), .B2(KEYINPUT29), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n288), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n236), .A2(KEYINPUT80), .A3(new_n267), .ZN(new_n415));
  INV_X1    g214(.A(new_n407), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n390), .A2(new_n359), .ZN(new_n418));
  OAI211_X1 g217(.A(KEYINPUT81), .B(new_n407), .C1(new_n409), .C2(KEYINPUT29), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n412), .A2(new_n417), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n414), .A2(new_n415), .A3(new_n362), .A4(new_n407), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n409), .A2(new_n416), .ZN(new_n422));
  INV_X1    g221(.A(new_n418), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  XOR2_X1   g223(.A(G8gat), .B(G36gat), .Z(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT82), .ZN(new_n426));
  XOR2_X1   g225(.A(G64gat), .B(G92gat), .Z(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n420), .A2(new_n424), .A3(KEYINPUT30), .A4(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n420), .A2(new_n424), .A3(new_n428), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n428), .B1(new_n420), .B2(new_n424), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT5), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n399), .A2(new_n289), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n378), .A2(new_n278), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G225gat), .A2(G233gat), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n437), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n378), .B2(new_n278), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n278), .A2(new_n397), .A3(new_n444), .A4(new_n398), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n378), .A2(KEYINPUT85), .A3(new_n444), .A4(new_n278), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n289), .B1(new_n378), .B2(new_n379), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n441), .B1(new_n391), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n443), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n399), .A2(KEYINPUT3), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(new_n289), .A3(new_n380), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n442), .A2(KEYINPUT5), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n445), .B1(KEYINPUT86), .B2(new_n446), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n439), .A2(KEYINPUT86), .A3(KEYINPUT4), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n455), .B(new_n456), .C1(new_n457), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n453), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g260(.A(G1gat), .B(G29gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT0), .ZN(new_n463));
  XNOR2_X1  g262(.A(G57gat), .B(G85gat), .ZN(new_n464));
  XOR2_X1   g263(.A(new_n463), .B(new_n464), .Z(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n467), .A2(KEYINPUT6), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n460), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT87), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n453), .A2(new_n460), .A3(new_n471), .A4(new_n465), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT6), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n467), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n406), .B1(new_n436), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n428), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n420), .A2(new_n424), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(KEYINPUT37), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n412), .A2(new_n417), .A3(new_n419), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n483), .A2(new_n484), .A3(new_n423), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n484), .B1(new_n483), .B2(new_n423), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n423), .B1(new_n421), .B2(new_n422), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n482), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n490), .A2(KEYINPUT92), .A3(new_n475), .A4(new_n432), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n483), .A2(new_n423), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT90), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n483), .A2(new_n484), .A3(new_n423), .ZN(new_n495));
  INV_X1    g294(.A(new_n487), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n481), .B1(new_n497), .B2(KEYINPUT37), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n475), .A2(new_n432), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n492), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n480), .A2(KEYINPUT37), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n428), .B1(new_n480), .B2(KEYINPUT37), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(new_n502), .B2(KEYINPUT93), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT93), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n489), .B1(new_n420), .B2(new_n424), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(new_n428), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n478), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n491), .A2(new_n500), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n405), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(new_n403), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n455), .B1(new_n457), .B2(new_n459), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT39), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(new_n513), .A3(new_n442), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT89), .B1(new_n515), .B2(new_n466), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n514), .A2(new_n517), .A3(new_n465), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n512), .A2(new_n442), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n520), .B(KEYINPUT39), .C1(new_n442), .C2(new_n440), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n519), .A2(KEYINPUT40), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT40), .B1(new_n519), .B2(new_n521), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n522), .A2(new_n523), .A3(new_n474), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n431), .A2(new_n435), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n511), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n477), .B1(new_n509), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n324), .A2(new_n331), .A3(new_n334), .A4(new_n406), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n525), .A2(new_n475), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT35), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n511), .A2(KEYINPUT35), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n336), .A2(new_n532), .A3(new_n529), .ZN(new_n533));
  AOI22_X1  g332(.A1(new_n337), .A2(new_n527), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G183gat), .B(G211gat), .Z(new_n536));
  XNOR2_X1  g335(.A(G57gat), .B(G64gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT104), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT9), .ZN(new_n539));
  NAND2_X1  g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n537), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n538), .B2(new_n537), .ZN(new_n542));
  INV_X1    g341(.A(G71gat), .ZN(new_n543));
  INV_X1    g342(.A(G78gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT103), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT103), .B1(new_n543), .B2(new_n544), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT102), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n540), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT102), .B1(G71gat), .B2(G78gat), .ZN(new_n551));
  NOR4_X1   g350(.A1(new_n547), .A2(new_n548), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n542), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(KEYINPUT105), .A2(G57gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(G64gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n540), .B1(new_n545), .B2(new_n539), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT106), .B(KEYINPUT21), .Z(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(G127gat), .B(G155gat), .Z(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  XOR2_X1   g363(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n562), .B(new_n563), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n565), .ZN(new_n569));
  XNOR2_X1  g368(.A(G15gat), .B(G22gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT16), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(G1gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT101), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n572), .B(new_n573), .C1(G1gat), .C2(new_n570), .ZN(new_n574));
  INV_X1    g373(.A(G8gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n577), .B1(KEYINPUT21), .B2(new_n558), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n567), .A2(new_n569), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n567), .B2(new_n569), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n536), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n569), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n578), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n567), .A2(new_n569), .A3(new_n579), .ZN(new_n585));
  INV_X1    g384(.A(new_n536), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G43gat), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT15), .B1(new_n589), .B2(G50gat), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n590), .B1(new_n589), .B2(G50gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(G29gat), .A2(G36gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT96), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(G29gat), .A2(G36gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT14), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n591), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT14), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n595), .B(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n591), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n593), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n594), .A2(KEYINPUT100), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n596), .A2(KEYINPUT99), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n601), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT97), .B(G43gat), .ZN(new_n607));
  INV_X1    g406(.A(G50gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n609), .A2(KEYINPUT98), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n609), .A2(KEYINPUT98), .B1(new_n589), .B2(G50gat), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT15), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n597), .B1(new_n606), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT17), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT7), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(KEYINPUT107), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(KEYINPUT107), .ZN(new_n617));
  AND2_X1   g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT8), .ZN(new_n623));
  OAI22_X1  g422(.A1(new_n622), .A2(new_n623), .B1(G85gat), .B2(G92gat), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G99gat), .B(G106gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT108), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n630), .ZN(new_n632));
  AND2_X1   g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n632), .A2(new_n613), .B1(KEYINPUT41), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G190gat), .B(G218gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(KEYINPUT111), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n633), .A2(KEYINPUT41), .ZN(new_n640));
  XNOR2_X1  g439(.A(G134gat), .B(G162gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  NOR2_X1   g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n635), .A2(new_n637), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT109), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n635), .A2(KEYINPUT109), .A3(new_n637), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n638), .A2(KEYINPUT111), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n643), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n638), .B1(new_n646), .B2(new_n647), .ZN(new_n651));
  INV_X1    g450(.A(new_n642), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT110), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OR3_X1    g452(.A1(new_n651), .A2(KEYINPUT110), .A3(new_n652), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n588), .A2(new_n650), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n614), .A2(new_n576), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n577), .A2(new_n613), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G229gat), .A2(G233gat), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(KEYINPUT18), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(KEYINPUT18), .A3(new_n659), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n577), .B(new_n613), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n659), .B(KEYINPUT13), .Z(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT95), .B1(new_n661), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G113gat), .B(G141gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(G169gat), .B(G197gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT94), .B(KEYINPUT11), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT12), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g474(.A(KEYINPUT95), .B(new_n673), .C1(new_n661), .C2(new_n666), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(G230gat), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(new_n386), .ZN(new_n679));
  INV_X1    g478(.A(new_n558), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n630), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT10), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n630), .A2(new_n680), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n681), .A2(KEYINPUT10), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n679), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  AOI211_X1 g486(.A(new_n678), .B(new_n386), .C1(new_n682), .C2(new_n684), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(G120gat), .B(G148gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT112), .ZN(new_n691));
  XNOR2_X1  g490(.A(G176gat), .B(G204gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n689), .A2(new_n694), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n655), .A2(new_n677), .A3(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n535), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n475), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g500(.A1(new_n571), .A2(new_n575), .ZN(new_n702));
  NAND2_X1  g501(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n699), .A2(new_n525), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(KEYINPUT42), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n699), .A2(new_n525), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n706), .B1(new_n707), .B2(G8gat), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n705), .B1(new_n704), .B2(new_n708), .ZN(G1325gat));
  INV_X1    g508(.A(new_n699), .ZN(new_n710));
  INV_X1    g509(.A(new_n336), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n710), .A2(G15gat), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G15gat), .B1(new_n710), .B2(new_n337), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1326gat));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n511), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT43), .B(G22gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  NAND3_X1  g516(.A1(new_n654), .A2(new_n653), .A3(new_n650), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n531), .A2(new_n533), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n527), .A2(new_n337), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n588), .A2(new_n677), .A3(new_n697), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n724), .A2(G29gat), .A3(new_n476), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT45), .Z(new_n726));
  OR2_X1    g525(.A1(new_n722), .A2(KEYINPUT44), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n722), .A2(KEYINPUT44), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n723), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n476), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n726), .A2(new_n731), .ZN(G1328gat));
  OAI21_X1  g531(.A(G36gat), .B1(new_n730), .B2(new_n436), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n724), .A2(G36gat), .A3(new_n436), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT46), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1329gat));
  NOR2_X1   g535(.A1(new_n724), .A2(new_n711), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n737), .A2(new_n607), .ZN(new_n738));
  INV_X1    g537(.A(new_n337), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n607), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n730), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT47), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n743), .B(new_n738), .C1(new_n730), .C2(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(G1330gat));
  NAND4_X1  g544(.A1(new_n727), .A2(new_n511), .A3(new_n723), .A4(new_n728), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G50gat), .ZN(new_n747));
  AOI21_X1  g546(.A(KEYINPUT48), .B1(new_n747), .B2(KEYINPUT113), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n722), .A2(new_n608), .A3(new_n511), .A4(new_n723), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n747), .B(new_n749), .C1(KEYINPUT113), .C2(KEYINPUT48), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(G1331gat));
  INV_X1    g552(.A(new_n677), .ZN(new_n754));
  INV_X1    g553(.A(new_n697), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n534), .A2(new_n655), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n475), .B(KEYINPUT114), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g559(.A(new_n436), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n762), .A2(KEYINPUT115), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(KEYINPUT115), .ZN(new_n764));
  OR2_X1    g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n765), .B1(new_n763), .B2(new_n764), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(G1333gat));
  AOI21_X1  g567(.A(new_n543), .B1(new_n756), .B2(new_n739), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n711), .A2(G71gat), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n769), .B1(new_n756), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n511), .ZN(new_n773));
  XOR2_X1   g572(.A(KEYINPUT116), .B(G78gat), .Z(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1335gat));
  NOR2_X1   g574(.A1(new_n754), .A2(new_n588), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n755), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n729), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G85gat), .B1(new_n779), .B2(new_n476), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n527), .A2(new_n337), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n332), .B(KEYINPUT75), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n784), .A2(new_n529), .A3(new_n324), .A4(new_n406), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n532), .A2(new_n529), .ZN(new_n786));
  AOI22_X1  g585(.A1(new_n785), .A2(KEYINPUT35), .B1(new_n786), .B2(new_n336), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n782), .B(new_n718), .C1(new_n783), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n776), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n722), .A2(new_n782), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n781), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n777), .B1(new_n722), .B2(new_n782), .ZN(new_n792));
  OAI21_X1  g591(.A(KEYINPUT117), .B1(new_n534), .B2(new_n719), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(KEYINPUT51), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  OR3_X1    g595(.A1(new_n755), .A2(G85gat), .A3(new_n476), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n780), .B1(new_n796), .B2(new_n797), .ZN(G1336gat));
  NOR3_X1   g597(.A1(new_n755), .A2(new_n436), .A3(G92gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n727), .A2(new_n525), .A3(new_n728), .A4(new_n778), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(new_n801), .B2(G92gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n801), .A2(G92gat), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n793), .A2(new_n805), .A3(new_n788), .A4(new_n776), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT51), .B1(new_n806), .B2(KEYINPUT120), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT119), .B1(KEYINPUT120), .B2(KEYINPUT51), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n792), .B2(new_n793), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n799), .B(KEYINPUT118), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n804), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n803), .B1(new_n812), .B2(new_n813), .ZN(G1337gat));
  OAI21_X1  g613(.A(G99gat), .B1(new_n779), .B2(new_n337), .ZN(new_n815));
  OR3_X1    g614(.A1(new_n711), .A2(G99gat), .A3(new_n755), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n796), .B2(new_n816), .ZN(G1338gat));
  NAND4_X1  g616(.A1(new_n727), .A2(new_n511), .A3(new_n728), .A4(new_n778), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT53), .B1(new_n818), .B2(G106gat), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT121), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n755), .A2(G106gat), .A3(new_n406), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n820), .B1(new_n795), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n821), .ZN(new_n823));
  AOI211_X1 g622(.A(KEYINPUT121), .B(new_n823), .C1(new_n791), .C2(new_n794), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n819), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n807), .A2(new_n809), .A3(new_n823), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n818), .A2(G106gat), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT53), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(G1339gat));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n687), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n685), .A2(new_n686), .A3(new_n679), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n693), .B1(new_n687), .B2(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n834), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n837), .A2(new_n695), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n677), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n666), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n841), .B(new_n673), .C1(new_n660), .C2(KEYINPUT18), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n658), .A2(new_n659), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n663), .A2(new_n664), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n672), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n755), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n719), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n839), .B1(KEYINPUT122), .B2(new_n846), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n846), .A2(KEYINPUT122), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n850), .A3(new_n718), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n588), .B1(new_n848), .B2(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n655), .A2(new_n754), .A3(new_n697), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n854), .A2(new_n436), .A3(new_n758), .ZN(new_n855));
  INV_X1    g654(.A(new_n528), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858), .B2(new_n754), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n854), .A2(new_n406), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n336), .A2(new_n475), .A3(new_n436), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n754), .A2(G113gat), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(G1340gat));
  INV_X1    g663(.A(new_n862), .ZN(new_n865));
  OAI21_X1  g664(.A(G120gat), .B1(new_n865), .B2(new_n755), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n755), .A2(G120gat), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT123), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n866), .B1(new_n857), .B2(new_n868), .ZN(G1341gat));
  INV_X1    g668(.A(new_n588), .ZN(new_n870));
  OAI21_X1  g669(.A(G127gat), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n588), .A2(new_n273), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n857), .B2(new_n872), .ZN(G1342gat));
  OAI21_X1  g672(.A(G134gat), .B1(new_n865), .B2(new_n719), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n855), .A2(new_n275), .A3(new_n856), .A4(new_n718), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT56), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(G1343gat));
  NAND2_X1  g678(.A1(new_n837), .A2(KEYINPUT124), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n835), .A2(new_n881), .A3(new_n836), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n880), .A2(new_n695), .A3(new_n838), .A4(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n677), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n719), .B1(new_n884), .B2(new_n847), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n588), .B1(new_n885), .B2(new_n851), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n511), .B1(new_n886), .B2(new_n853), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n889), .B(new_n511), .C1(new_n852), .C2(new_n853), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n739), .A2(new_n476), .A3(new_n525), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n888), .A2(new_n754), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G141gat), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n739), .A2(new_n406), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n855), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n677), .A2(G141gat), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT125), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n893), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT58), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n893), .B(new_n900), .C1(new_n895), .C2(new_n897), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1344gat));
  OR3_X1    g701(.A1(new_n895), .A2(G148gat), .A3(new_n755), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n695), .A2(new_n838), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n881), .B1(new_n835), .B2(new_n836), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT124), .B(KEYINPUT55), .C1(new_n833), .C2(new_n834), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n847), .B1(new_n908), .B2(new_n754), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n851), .B1(new_n909), .B2(new_n718), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n853), .B1(new_n910), .B2(new_n870), .ZN(new_n911));
  OAI211_X1 g710(.A(KEYINPUT126), .B(new_n889), .C1(new_n911), .C2(new_n406), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT57), .B(new_n511), .C1(new_n852), .C2(new_n853), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT126), .B1(new_n887), .B2(new_n889), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n697), .B(new_n891), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n904), .B1(new_n916), .B2(G148gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n888), .A2(new_n890), .A3(new_n891), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n755), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n904), .A2(G148gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n903), .B1(new_n917), .B2(new_n921), .ZN(G1345gat));
  OAI21_X1  g721(.A(G155gat), .B1(new_n918), .B2(new_n870), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n870), .A2(G155gat), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n895), .B2(new_n924), .ZN(G1346gat));
  OAI21_X1  g724(.A(G162gat), .B1(new_n918), .B2(new_n719), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n719), .A2(G162gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n895), .B2(new_n927), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n436), .A2(new_n475), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n854), .A2(new_n856), .A3(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n754), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n336), .A2(new_n525), .A3(new_n757), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n860), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n754), .A2(G169gat), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(G1348gat));
  INV_X1    g735(.A(G176gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n931), .A2(new_n937), .A3(new_n697), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n860), .A2(new_n755), .A3(new_n933), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n939), .B2(new_n937), .ZN(G1349gat));
  NOR3_X1   g739(.A1(new_n860), .A2(new_n870), .A3(new_n933), .ZN(new_n941));
  INV_X1    g740(.A(new_n284), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n870), .A2(new_n207), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n930), .A2(new_n944), .ZN(new_n945));
  OR3_X1    g744(.A1(new_n943), .A2(KEYINPUT60), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT60), .B1(new_n943), .B2(new_n945), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1350gat));
  NAND3_X1  g747(.A1(new_n931), .A2(new_n211), .A3(new_n718), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n718), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(G190gat), .ZN(new_n952));
  AOI211_X1 g751(.A(KEYINPUT61), .B(new_n211), .C1(new_n934), .C2(new_n718), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(G1351gat));
  NAND3_X1  g753(.A1(new_n854), .A2(new_n894), .A3(new_n929), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n956), .A2(new_n348), .A3(new_n754), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT127), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n739), .A2(new_n436), .A3(new_n758), .ZN(new_n959));
  OAI211_X1 g758(.A(new_n754), .B(new_n959), .C1(new_n914), .C2(new_n915), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n958), .B1(new_n961), .B2(new_n348), .ZN(G1352gat));
  NOR3_X1   g761(.A1(new_n955), .A2(G204gat), .A3(new_n755), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT62), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n697), .B(new_n959), .C1(new_n914), .C2(new_n915), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n964), .B1(new_n346), .B2(new_n966), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n956), .A2(new_n343), .A3(new_n588), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n588), .B(new_n959), .C1(new_n914), .C2(new_n915), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(G1354gat));
  NAND3_X1  g771(.A1(new_n956), .A2(new_n344), .A3(new_n718), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n718), .B(new_n959), .C1(new_n914), .C2(new_n915), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n973), .B1(new_n975), .B2(new_n344), .ZN(G1355gat));
endmodule


