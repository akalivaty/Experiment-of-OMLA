//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n559, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT66), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G221), .A3(G220), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n463), .A2(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n464), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(new_n468), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n465), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n471), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  AND2_X1   g056(.A1(new_n466), .A2(new_n468), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n482), .A2(G2105), .A3(new_n464), .ZN(new_n483));
  INV_X1    g058(.A(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n467), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n483), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(G136), .B2(new_n470), .ZN(G162));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  AND2_X1   g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n482), .A2(new_n490), .A3(new_n464), .A4(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n464), .A2(new_n466), .A3(new_n468), .A4(new_n491), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT69), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(KEYINPUT70), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n467), .A2(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(new_n495), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n492), .A2(new_n494), .A3(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n473), .A2(new_n468), .A3(G138), .A4(new_n467), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT4), .A2(G138), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n469), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n489), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n508), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n470), .A2(new_n511), .B1(new_n506), .B2(new_n505), .ZN(new_n512));
  AND4_X1   g087(.A1(new_n464), .A2(new_n466), .A3(new_n468), .A4(new_n491), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(new_n490), .B1(new_n499), .B2(new_n502), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT71), .A4(new_n494), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(new_n515), .ZN(G164));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT6), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n520), .A2(G543), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n520), .A2(new_n522), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G88), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n528), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(new_n521), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n525), .A2(new_n530), .A3(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND2_X1  g109(.A1(new_n524), .A2(G51), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n529), .A2(G89), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n528), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n535), .A2(new_n536), .A3(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND2_X1  g118(.A1(new_n524), .A2(G52), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n529), .A2(G90), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n521), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n524), .A2(G43), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n529), .A2(G81), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n521), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT73), .Z(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g133(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n559));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n528), .A2(KEYINPUT77), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n526), .A2(new_n565), .A3(new_n527), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n563), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  OR3_X1    g144(.A1(new_n567), .A2(KEYINPUT78), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g145(.A(KEYINPUT78), .B1(new_n567), .B2(new_n569), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n570), .A2(G651), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT79), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n574));
  AND2_X1   g149(.A1(G53), .A2(G543), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n520), .A2(new_n574), .A3(new_n522), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT75), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(KEYINPUT9), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n520), .A2(new_n579), .A3(new_n522), .A4(new_n575), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n580), .A2(KEYINPUT9), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n578), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n570), .A2(new_n583), .A3(new_n571), .A4(G651), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n529), .A2(G91), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n573), .A2(new_n582), .A3(new_n584), .A4(new_n585), .ZN(G299));
  NAND2_X1  g161(.A1(new_n524), .A2(G49), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n529), .A2(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n528), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(new_n521), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n520), .A2(G48), .A3(G543), .A4(new_n522), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n520), .A2(G86), .A3(new_n522), .A4(new_n528), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(new_n524), .A2(G47), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n529), .A2(G85), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n596), .B(new_n597), .C1(new_n521), .C2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT80), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n529), .A2(G92), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G54), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n604), .B1(new_n523), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n605), .B2(new_n523), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(new_n564), .B2(new_n566), .ZN(new_n609));
  AND2_X1   g184(.A1(G79), .A2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(G651), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(KEYINPUT82), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n607), .A2(new_n614), .A3(new_n611), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n603), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n601), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n601), .B1(new_n616), .B2(G868), .ZN(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G299), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n619), .B2(G168), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(new_n619), .B2(G168), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n616), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g203(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT13), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n633));
  AOI22_X1  g208(.A1(new_n631), .A2(new_n632), .B1(new_n633), .B2(G2100), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n632), .B2(new_n631), .ZN(new_n635));
  OR3_X1    g210(.A1(new_n635), .A2(new_n633), .A3(G2100), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(new_n633), .B2(G2100), .ZN(new_n637));
  INV_X1    g212(.A(G123), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n467), .A2(G111), .ZN(new_n639));
  OAI21_X1  g214(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n640));
  OAI22_X1  g215(.A1(new_n483), .A2(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(G135), .B2(new_n470), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT84), .B(G2096), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n636), .A2(new_n637), .A3(new_n644), .ZN(G156));
  XOR2_X1   g220(.A(G1341), .B(G1348), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT86), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n649), .B(new_n655), .Z(new_n656));
  XOR2_X1   g231(.A(G2443), .B(G2446), .Z(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n659), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n660), .A2(G14), .A3(new_n661), .ZN(G401));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT17), .Z(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n665), .B2(new_n663), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT87), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n665), .A3(new_n663), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT18), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n669), .A2(new_n665), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n674), .B1(new_n664), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2096), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT88), .B(G2100), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1956), .B(G2474), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NOR3_X1   g261(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n685), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT20), .Z(new_n689));
  AOI211_X1 g264(.A(new_n687), .B(new_n689), .C1(new_n682), .C2(new_n686), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT89), .ZN(new_n691));
  XOR2_X1   g266(.A(G1981), .B(G1986), .Z(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n691), .B(new_n696), .ZN(G229));
  MUX2_X1   g272(.A(G23), .B(G288), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT33), .B(G1976), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G22), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(G1971), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  MUX2_X1   g280(.A(G6), .B(G305), .S(G16), .Z(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n700), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n710), .A2(new_n711), .ZN(new_n713));
  MUX2_X1   g288(.A(G24), .B(G290), .S(G16), .Z(new_n714));
  INV_X1    g289(.A(G1986), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G25), .ZN(new_n718));
  INV_X1    g293(.A(G95), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n719), .A2(new_n467), .A3(KEYINPUT90), .ZN(new_n720));
  AOI21_X1  g295(.A(KEYINPUT90), .B1(new_n719), .B2(new_n467), .ZN(new_n721));
  OAI221_X1 g296(.A(G2104), .B1(G107), .B2(new_n467), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G119), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n483), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G131), .B2(new_n470), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n718), .B1(new_n725), .B2(new_n717), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n712), .A2(new_n713), .A3(new_n716), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT36), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n717), .A2(G32), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT26), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n734), .A2(new_n735), .B1(G105), .B2(new_n478), .ZN(new_n736));
  INV_X1    g311(.A(G141), .ZN(new_n737));
  INV_X1    g312(.A(G129), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n736), .B1(new_n737), .B2(new_n469), .C1(new_n483), .C2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT93), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n740), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n731), .B1(new_n744), .B2(new_n717), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT27), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1996), .ZN(new_n747));
  NOR2_X1   g322(.A1(G27), .A2(G29), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G164), .B2(G29), .ZN(new_n749));
  INV_X1    g324(.A(G2078), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n717), .A2(G33), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT25), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n473), .A2(new_n468), .A3(G127), .ZN(new_n755));
  NAND2_X1  g330(.A1(G115), .A2(G2104), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n467), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n754), .B(new_n757), .C1(G139), .C2(new_n470), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n752), .B1(new_n758), .B2(new_n717), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT92), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G2072), .ZN(new_n761));
  NOR2_X1   g336(.A1(G286), .A2(new_n701), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(KEYINPUT94), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT94), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G16), .B2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n763), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G1966), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n701), .A2(G5), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G171), .B2(new_n701), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(G1961), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT31), .B(G11), .ZN(new_n771));
  INV_X1    g346(.A(G28), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n772), .B2(KEYINPUT30), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(KEYINPUT95), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(KEYINPUT30), .B2(new_n772), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(KEYINPUT95), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n771), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n642), .B2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G2084), .ZN(new_n779));
  INV_X1    g354(.A(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n780), .B2(KEYINPUT24), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(KEYINPUT24), .B2(new_n780), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n480), .B2(new_n717), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n778), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G1961), .B2(new_n769), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n761), .A2(new_n767), .A3(new_n770), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n779), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT96), .Z(new_n788));
  OAI22_X1  g363(.A1(new_n760), .A2(G2072), .B1(new_n766), .B2(G1966), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n747), .A2(new_n751), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n701), .A2(G20), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT23), .Z(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G299), .B2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1956), .ZN(new_n798));
  NOR2_X1   g373(.A1(G29), .A2(G35), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G162), .B2(G29), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G2090), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n701), .A2(G19), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n555), .B2(new_n701), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1341), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n717), .A2(G26), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT28), .ZN(new_n810));
  INV_X1    g385(.A(G128), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n467), .A2(G116), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n483), .A2(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G140), .B2(new_n470), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n810), .B1(new_n815), .B2(new_n717), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G2067), .ZN(new_n817));
  NOR4_X1   g392(.A1(new_n804), .A2(new_n805), .A3(new_n808), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n701), .A2(G4), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n616), .B2(new_n701), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(G1348), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(G1348), .ZN(new_n822));
  AND4_X1   g397(.A1(new_n798), .A2(new_n818), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n730), .A2(new_n793), .A3(new_n794), .A4(new_n823), .ZN(G150));
  INV_X1    g399(.A(G150), .ZN(G311));
  XOR2_X1   g400(.A(KEYINPUT100), .B(G860), .Z(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n616), .A2(G559), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT99), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n524), .A2(G55), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n529), .A2(G93), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n831), .B(new_n832), .C1(new_n521), .C2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(new_n554), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n554), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n830), .B(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n827), .B1(new_n840), .B2(KEYINPUT39), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(KEYINPUT39), .B2(new_n840), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n834), .A2(new_n827), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(G145));
  XNOR2_X1  g420(.A(new_n743), .B(new_n815), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT70), .B1(new_n496), .B2(new_n498), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n501), .A2(new_n495), .A3(new_n500), .ZN(new_n848));
  OAI22_X1  g423(.A1(new_n847), .A2(new_n848), .B1(new_n493), .B2(KEYINPUT69), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n493), .A2(KEYINPUT69), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT101), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n492), .A2(new_n494), .A3(new_n503), .A4(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(KEYINPUT102), .B1(new_n854), .B2(new_n512), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n856));
  AOI211_X1 g431(.A(new_n856), .B(new_n509), .C1(new_n851), .C2(new_n853), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n846), .B(new_n858), .Z(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n758), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n725), .B(new_n631), .ZN(new_n861));
  INV_X1    g436(.A(G130), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n467), .A2(KEYINPUT104), .A3(G118), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT104), .B1(new_n467), .B2(G118), .ZN(new_n864));
  OR2_X1    g439(.A1(G106), .A2(G2105), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(G2104), .A3(new_n865), .ZN(new_n866));
  OAI22_X1  g441(.A1(new_n483), .A2(new_n862), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT103), .ZN(new_n868));
  INV_X1    g443(.A(G142), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n868), .B1(new_n469), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n470), .A2(KEYINPUT103), .A3(G142), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n861), .B(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT105), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n860), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n642), .B(new_n480), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G162), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n877), .B1(new_n860), .B2(new_n874), .ZN(new_n880));
  INV_X1    g455(.A(new_n873), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n860), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g459(.A1(new_n834), .A2(new_n619), .ZN(new_n885));
  XNOR2_X1  g460(.A(G303), .B(G305), .ZN(new_n886));
  XNOR2_X1  g461(.A(G290), .B(G288), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT107), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n888), .B2(new_n887), .ZN(new_n890));
  INV_X1    g465(.A(new_n887), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n891), .A2(KEYINPUT107), .A3(new_n886), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT42), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n625), .B(new_n839), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n573), .A2(new_n584), .A3(new_n585), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n616), .A2(new_n896), .A3(new_n582), .ZN(new_n897));
  INV_X1    g472(.A(new_n603), .ZN(new_n898));
  INV_X1    g473(.A(new_n615), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n614), .B1(new_n607), .B2(new_n611), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(G299), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n895), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n903), .A2(KEYINPUT41), .ZN(new_n906));
  XOR2_X1   g481(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n897), .B2(new_n902), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n905), .B1(new_n895), .B2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n894), .B(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n885), .B1(new_n911), .B2(new_n619), .ZN(G295));
  OAI21_X1  g487(.A(new_n885), .B1(new_n911), .B2(new_n619), .ZN(G331));
  INV_X1    g488(.A(KEYINPUT110), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n915));
  INV_X1    g490(.A(new_n837), .ZN(new_n916));
  OAI21_X1  g491(.A(G171), .B1(new_n916), .B2(new_n835), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n836), .A2(G301), .A3(new_n837), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(G168), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G168), .B1(new_n917), .B2(new_n918), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n906), .B2(new_n908), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n904), .B1(new_n920), .B2(new_n921), .ZN(new_n924));
  INV_X1    g499(.A(new_n893), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n893), .B(KEYINPUT108), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n923), .A2(new_n924), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT109), .A4(new_n925), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n928), .A2(new_n931), .A3(new_n879), .A4(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(G37), .B1(new_n926), .B2(new_n927), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n903), .A2(new_n907), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n937), .B(new_n922), .C1(KEYINPUT41), .C2(new_n904), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(new_n924), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(new_n929), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n936), .A2(new_n940), .A3(KEYINPUT43), .A4(new_n932), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n915), .B1(new_n935), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n936), .A2(new_n940), .A3(new_n934), .A4(new_n932), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n915), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n914), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT44), .B1(new_n944), .B2(new_n945), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n942), .A2(new_n949), .A3(KEYINPUT110), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n948), .A2(new_n950), .ZN(G397));
  INV_X1    g526(.A(KEYINPUT127), .ZN(new_n952));
  NAND2_X1  g527(.A1(G160), .A2(G40), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n852), .B1(new_n514), .B2(new_n494), .ZN(new_n954));
  AND4_X1   g529(.A1(new_n852), .A2(new_n492), .A3(new_n494), .A4(new_n503), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n512), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n856), .ZN(new_n957));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n509), .B1(new_n851), .B2(new_n853), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT102), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n957), .A2(new_n958), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G2067), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n815), .B(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT111), .ZN(new_n966));
  INV_X1    g541(.A(G1996), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n743), .B(new_n967), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n725), .B(new_n727), .Z(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(G290), .B(new_n715), .ZN(new_n973));
  AOI211_X1 g548(.A(new_n953), .B(new_n963), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G8), .ZN(new_n975));
  INV_X1    g550(.A(G1966), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n962), .B1(new_n959), .B2(G1384), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n978));
  INV_X1    g553(.A(new_n953), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n510), .A2(new_n515), .A3(new_n958), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(new_n962), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n978), .B1(new_n977), .B2(new_n979), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n976), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(G1384), .B1(new_n854), .B2(new_n512), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n953), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n981), .A2(new_n989), .A3(KEYINPUT50), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n981), .B2(KEYINPUT50), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n988), .B(new_n779), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n975), .B1(new_n985), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(G286), .A2(G8), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n993), .A2(KEYINPUT51), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n985), .A2(new_n992), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(G8), .A3(G168), .ZN(new_n998));
  XOR2_X1   g573(.A(new_n994), .B(KEYINPUT123), .Z(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(new_n993), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g575(.A(KEYINPUT122), .B(KEYINPUT51), .Z(new_n1001));
  AOI21_X1  g576(.A(new_n996), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n984), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(G2078), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1003), .A2(new_n982), .A3(new_n980), .A4(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n1007));
  INV_X1    g582(.A(G1961), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n962), .A2(G1384), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n957), .A2(new_n960), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n953), .B1(new_n981), .B2(new_n962), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n750), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT124), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1013), .A2(new_n1014), .A3(new_n1004), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1014), .B1(new_n1013), .B2(new_n1004), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1006), .B(new_n1009), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT125), .B1(new_n1017), .B2(G171), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1013), .A2(new_n1004), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT124), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1013), .A2(new_n1014), .A3(new_n1004), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT125), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(G301), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n979), .A2(new_n1005), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1027), .B1(new_n858), .B2(new_n1010), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1008), .A2(new_n1007), .B1(new_n1028), .B2(new_n963), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1026), .B1(new_n1030), .B2(G171), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1018), .A2(new_n1025), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G305), .A2(G1981), .ZN(new_n1033));
  INV_X1    g608(.A(G1981), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1033), .A2(KEYINPUT49), .A3(new_n1035), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n959), .A2(new_n953), .A3(G1384), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(new_n975), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n587), .A2(new_n588), .A3(G1976), .A4(new_n589), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT114), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1042), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1043), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1971), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n986), .A2(new_n987), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n979), .B1(new_n981), .B2(KEYINPUT50), .ZN(new_n1055));
  NOR3_X1   g630(.A1(new_n1054), .A2(new_n1055), .A3(G2090), .ZN(new_n1056));
  OAI21_X1  g631(.A(G8), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(G303), .A2(G8), .ZN(new_n1058));
  NOR2_X1   g633(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT113), .B(KEYINPUT55), .Z(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1057), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n988), .B(new_n803), .C1(new_n990), .C2(new_n991), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(G8), .B1(new_n1066), .B2(new_n1053), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1052), .B(new_n1064), .C1(new_n1063), .C2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(G301), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1029), .B(G301), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1026), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1002), .A2(new_n1032), .A3(new_n1069), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT126), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1017), .A2(G171), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1071), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1068), .B1(new_n1077), .B2(new_n1026), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT126), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n1032), .A4(new_n1002), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n573), .A2(new_n1081), .A3(new_n584), .A4(new_n585), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n1083));
  AND3_X1   g658(.A1(G299), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(G299), .B1(new_n1083), .B2(new_n1082), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1011), .A2(new_n1012), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1956), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1090), .B(new_n1088), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT61), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n986), .A2(new_n979), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1041), .A2(KEYINPUT120), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT58), .B(G1341), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1101));
  OAI22_X1  g676(.A1(new_n1099), .A2(new_n1100), .B1(new_n1101), .B2(G1996), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1102), .A2(KEYINPUT59), .A3(new_n555), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT59), .B1(new_n1102), .B2(new_n555), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n1094), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1099), .A2(new_n964), .ZN(new_n1106));
  INV_X1    g681(.A(G1348), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1007), .A2(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(KEYINPUT60), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT60), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT121), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n901), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1111), .A2(new_n1116), .A3(new_n1114), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1092), .A2(KEYINPUT61), .A3(new_n1093), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1105), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1092), .B1(new_n1109), .B2(new_n901), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1093), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1075), .A2(new_n1080), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1063), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1101), .A2(new_n704), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n975), .B1(new_n1127), .B2(new_n1065), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1052), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(G288), .A2(G1976), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1043), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT115), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(new_n1132), .A3(new_n1035), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1130), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1035), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT115), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1133), .A2(new_n1042), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1129), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT116), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1129), .A2(new_n1138), .A3(KEYINPUT116), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(KEYINPUT118), .B(KEYINPUT63), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1068), .B2(new_n998), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n1067), .B2(new_n1063), .ZN(new_n1147));
  AOI211_X1 g722(.A(new_n975), .B(G286), .C1(new_n985), .C2(new_n992), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1128), .A2(new_n1126), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1052), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1143), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n993), .A2(new_n999), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1001), .B1(new_n1153), .B2(new_n1148), .ZN(new_n1154));
  INV_X1    g729(.A(new_n996), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1154), .A2(KEYINPUT62), .A3(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1076), .A2(new_n1068), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1152), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n974), .B1(new_n1125), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n963), .A2(new_n953), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n971), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT48), .ZN(new_n1165));
  NOR2_X1   g740(.A1(G290), .A2(G1986), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1164), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1168), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n969), .A2(new_n727), .A3(new_n725), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n815), .A2(new_n964), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1169), .B1(new_n1163), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1163), .A2(new_n967), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT46), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n966), .A2(new_n744), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1163), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT47), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n952), .B1(new_n1162), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1180), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1141), .A2(new_n1142), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1183), .B1(new_n1158), .B2(new_n1184), .ZN(new_n1185));
  AOI22_X1  g760(.A1(new_n1074), .A2(KEYINPUT126), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1185), .B1(new_n1186), .B2(new_n1080), .ZN(new_n1187));
  OAI211_X1 g762(.A(KEYINPUT127), .B(new_n1182), .C1(new_n1187), .C2(new_n974), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1181), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g764(.A1(G229), .A2(G227), .A3(new_n460), .A4(G401), .ZN(new_n1191));
  NAND3_X1  g765(.A1(new_n883), .A2(new_n946), .A3(new_n1191), .ZN(G225));
  INV_X1    g766(.A(G225), .ZN(G308));
endmodule


