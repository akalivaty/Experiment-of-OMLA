//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  INV_X1    g0008(.A(G50), .ZN(new_n209));
  INV_X1    g0009(.A(G226), .ZN(new_n210));
  INV_X1    g0010(.A(G116), .ZN(new_n211));
  INV_X1    g0011(.A(G270), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G58), .B2(G232), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT65), .B(G244), .Z(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G77), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G87), .A2(G250), .ZN(new_n218));
  NAND4_X1  g0018(.A1(new_n214), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n201), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n208), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(new_n201), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(KEYINPUT64), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n232), .B1(new_n208), .B2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(G13), .ZN(new_n234));
  NAND4_X1  g0034(.A1(new_n234), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n236), .B(G250), .C1(G257), .C2(G264), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT0), .ZN(new_n238));
  NAND3_X1  g0038(.A1(new_n223), .A2(new_n231), .A3(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(new_n239), .ZN(G361));
  XOR2_X1   g0040(.A(G238), .B(G244), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT2), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n210), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G264), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G270), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G358));
  XOR2_X1   g0049(.A(KEYINPUT68), .B(KEYINPUT69), .Z(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G97), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G68), .A2(G77), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n203), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT67), .ZN(new_n257));
  XNOR2_X1  g0057(.A(G50), .B(G58), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n254), .B(new_n259), .ZN(G351));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G223), .A3(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G222), .ZN(new_n265));
  OAI221_X1 g0065(.A(new_n262), .B1(new_n202), .B2(new_n261), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  OAI211_X1 g0075(.A(G1), .B(G13), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n270), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n273), .B1(new_n277), .B2(new_n210), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n278), .A2(KEYINPUT70), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(KEYINPUT70), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n268), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G169), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(G20), .B1(new_n225), .B2(G50), .ZN(new_n284));
  INV_X1    g0084(.A(G150), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n229), .A2(new_n274), .ZN(new_n286));
  XOR2_X1   g0086(.A(KEYINPUT8), .B(G58), .Z(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT71), .B1(new_n274), .B2(G20), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT71), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(new_n229), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n284), .B1(new_n285), .B2(new_n286), .C1(new_n288), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n228), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n269), .A2(G13), .A3(G20), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n209), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n295), .B1(new_n269), .B2(G20), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G50), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n296), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT72), .B(G179), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n302), .B1(new_n281), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n283), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT9), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G190), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n281), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n281), .A2(G200), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n302), .A2(new_n307), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n308), .A2(new_n310), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT10), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n311), .B2(KEYINPUT74), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n315), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n306), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n300), .A2(G77), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT73), .ZN(new_n321));
  INV_X1    g0121(.A(new_n295), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT15), .B(G87), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n292), .A2(new_n323), .B1(new_n229), .B2(new_n202), .ZN(new_n324));
  INV_X1    g0124(.A(new_n286), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(new_n287), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n321), .B1(G77), .B2(new_n297), .C1(new_n322), .C2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n261), .A2(G238), .A3(G1698), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n261), .A2(G232), .A3(new_n263), .ZN(new_n329));
  INV_X1    g0129(.A(G107), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(new_n261), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n267), .ZN(new_n332));
  INV_X1    g0132(.A(new_n277), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n215), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n273), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n282), .ZN(new_n336));
  OR2_X1    g0136(.A1(new_n335), .A2(new_n304), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n327), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n261), .A2(G232), .A3(G1698), .ZN(new_n340));
  NAND2_X1  g0140(.A1(G33), .A2(G97), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n340), .B(new_n341), .C1(new_n264), .C2(new_n210), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n272), .B1(new_n342), .B2(new_n267), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT13), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n333), .A2(G238), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n344), .B1(new_n343), .B2(new_n345), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT14), .B1(new_n348), .B2(new_n282), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(G179), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT14), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n351), .B(G169), .C1(new_n346), .C2(new_n347), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n325), .A2(G50), .ZN(new_n354));
  XNOR2_X1  g0154(.A(new_n354), .B(KEYINPUT75), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n292), .A2(new_n202), .B1(new_n229), .B2(G68), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n295), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT11), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n300), .A2(G68), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n357), .B2(new_n358), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n297), .A2(G68), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT12), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n359), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n339), .B1(new_n353), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n348), .A2(G190), .ZN(new_n367));
  OAI21_X1  g0167(.A(G200), .B1(new_n346), .B2(new_n347), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n319), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G58), .A2(G68), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n229), .B1(new_n225), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(G159), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n286), .A2(new_n373), .ZN(new_n374));
  OR3_X1    g0174(.A1(new_n372), .A2(new_n374), .A3(KEYINPUT77), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT77), .B1(new_n372), .B2(new_n374), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT3), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n274), .ZN(new_n379));
  NAND2_X1  g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n379), .A2(KEYINPUT7), .A3(new_n229), .A4(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n379), .A2(KEYINPUT76), .A3(new_n380), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT76), .B1(new_n379), .B2(new_n380), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n229), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n382), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(KEYINPUT16), .B(new_n377), .C1(new_n387), .C2(new_n201), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT16), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n379), .A2(new_n229), .A3(new_n380), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(new_n386), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n201), .B1(new_n391), .B2(new_n381), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n372), .A2(new_n374), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n388), .A2(new_n394), .A3(new_n295), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n288), .A2(new_n297), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n300), .B2(new_n288), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n261), .A2(G226), .A3(G1698), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n261), .A2(G223), .A3(new_n263), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G33), .A2(G87), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n267), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n276), .A2(G232), .A3(new_n270), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n404), .A3(new_n273), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G200), .ZN(new_n406));
  AOI211_X1 g0206(.A(new_n403), .B(new_n272), .C1(new_n401), .C2(new_n267), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(G190), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n395), .A2(new_n397), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT17), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n402), .A2(new_n303), .A3(new_n404), .A4(new_n273), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n407), .B2(G169), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n395), .B2(new_n397), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n413), .B(KEYINPUT18), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n327), .B1(G200), .B2(new_n335), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n335), .A2(new_n309), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n410), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n370), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(KEYINPUT3), .A2(G33), .ZN(new_n420));
  NOR2_X1   g0220(.A1(KEYINPUT3), .A2(G33), .ZN(new_n421));
  OAI211_X1 g0221(.A(G264), .B(G1698), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT82), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n261), .A2(KEYINPUT82), .A3(G264), .A4(G1698), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n261), .A2(G257), .A3(new_n263), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n420), .A2(new_n421), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G303), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n424), .A2(new_n425), .A3(new_n426), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n267), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT5), .B(G41), .ZN(new_n431));
  INV_X1    g0231(.A(G45), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(G1), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(G270), .A3(new_n276), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n431), .A2(G274), .A3(new_n433), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n430), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n269), .A2(G33), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n322), .A2(new_n297), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G116), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n298), .A2(new_n211), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n294), .A2(new_n228), .B1(G20), .B2(new_n211), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G283), .ZN(new_n445));
  INV_X1    g0245(.A(G97), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n445), .B(new_n229), .C1(G33), .C2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT20), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n444), .A2(KEYINPUT20), .A3(new_n447), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n442), .B(new_n443), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n439), .A2(G169), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT21), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n282), .B1(new_n430), .B2(new_n438), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT21), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n437), .B1(new_n267), .B2(new_n429), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G179), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(KEYINPUT83), .B1(new_n458), .B2(new_n450), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n454), .A2(KEYINPUT21), .B1(G179), .B2(new_n456), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT83), .ZN(new_n461));
  INV_X1    g0261(.A(new_n450), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n453), .B1(new_n459), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G200), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n456), .A2(new_n465), .ZN(new_n466));
  AOI211_X1 g0266(.A(new_n450), .B(new_n466), .C1(G190), .C2(new_n456), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n229), .B(G87), .C1(new_n420), .C2(new_n421), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT22), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT22), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n261), .A2(new_n471), .A3(new_n229), .A4(G87), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n274), .A2(new_n211), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n229), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n229), .A2(G107), .ZN(new_n476));
  XNOR2_X1  g0276(.A(new_n476), .B(KEYINPUT23), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(KEYINPUT24), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT24), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n470), .A2(new_n472), .B1(new_n229), .B2(new_n474), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n477), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n295), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n441), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(new_n330), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n297), .A2(G107), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n487), .B(KEYINPUT25), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g0289(.A(G257), .B(G1698), .C1(new_n420), .C2(new_n421), .ZN(new_n490));
  OAI211_X1 g0290(.A(G250), .B(new_n263), .C1(new_n420), .C2(new_n421), .ZN(new_n491));
  INV_X1    g0291(.A(G294), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n490), .B(new_n491), .C1(new_n274), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n267), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT84), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n436), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n267), .B1(new_n433), .B2(new_n431), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(G264), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n493), .A2(KEYINPUT84), .A3(new_n267), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n496), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G169), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n493), .A2(new_n267), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n498), .A2(G264), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n436), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G179), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n489), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT85), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n489), .A2(new_n508), .A3(KEYINPUT85), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g0313(.A(G244), .B(G1698), .C1(new_n420), .C2(new_n421), .ZN(new_n514));
  OAI211_X1 g0314(.A(G238), .B(new_n263), .C1(new_n420), .C2(new_n421), .ZN(new_n515));
  INV_X1    g0315(.A(new_n474), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT79), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT79), .A4(new_n516), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n267), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n433), .A2(G274), .ZN(new_n523));
  XNOR2_X1  g0323(.A(new_n523), .B(KEYINPUT78), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n276), .B(G250), .C1(G1), .C2(new_n432), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(KEYINPUT80), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n276), .B1(new_n519), .B2(new_n520), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT80), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n529), .A2(new_n530), .A3(new_n526), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n303), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n289), .A2(new_n291), .A3(G97), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n261), .A2(new_n229), .A3(G68), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n229), .B1(new_n341), .B2(new_n534), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(G87), .B2(new_n206), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT81), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT81), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n535), .A2(new_n541), .A3(new_n536), .A4(new_n538), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n295), .A3(new_n542), .ZN(new_n543));
  OR2_X1    g0343(.A1(new_n484), .A2(new_n323), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n323), .A2(new_n298), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n522), .A2(KEYINPUT80), .A3(new_n527), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n530), .B1(new_n529), .B2(new_n526), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n282), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n532), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(G244), .B(new_n263), .C1(new_n420), .C2(new_n421), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n263), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n445), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n267), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n498), .A2(G257), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n436), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G200), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n391), .A2(new_n381), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G107), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT6), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n446), .A2(new_n330), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(new_n205), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n330), .A2(KEYINPUT6), .A3(G97), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n229), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n286), .A2(new_n202), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n563), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(new_n295), .B1(new_n446), .B2(new_n298), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n441), .A2(G97), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n558), .A2(G190), .A3(new_n436), .A4(new_n559), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n561), .A2(new_n573), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n560), .A2(new_n282), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n298), .A2(new_n446), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n330), .B1(new_n391), .B2(new_n381), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n579), .A2(new_n568), .A3(new_n570), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n578), .B(new_n574), .C1(new_n580), .C2(new_n322), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n558), .A2(new_n303), .A3(new_n436), .A4(new_n559), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n483), .A2(new_n486), .A3(new_n488), .ZN(new_n585));
  INV_X1    g0385(.A(new_n500), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT84), .B1(new_n493), .B2(new_n267), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n588), .A2(KEYINPUT86), .A3(new_n309), .A4(new_n499), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n496), .A2(new_n309), .A3(new_n499), .A4(new_n500), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT86), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n465), .B1(new_n503), .B2(new_n505), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n585), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(G190), .B1(new_n528), .B2(new_n531), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n548), .A2(G200), .A3(new_n549), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n441), .A2(G87), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n543), .A2(new_n545), .A3(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  AND4_X1   g0401(.A1(new_n551), .A2(new_n584), .A3(new_n595), .A4(new_n601), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n419), .A2(new_n468), .A3(new_n513), .A4(new_n602), .ZN(G372));
  NAND2_X1  g0403(.A1(new_n548), .A2(new_n549), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n546), .B1(new_n604), .B2(new_n303), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n529), .A2(new_n526), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n282), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n599), .B1(new_n604), .B2(G190), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(G200), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n605), .A2(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n576), .A2(new_n583), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n585), .B2(new_n594), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n478), .A2(KEYINPUT24), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n481), .A2(new_n480), .A3(new_n477), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n485), .B1(new_n616), .B2(new_n295), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n617), .A2(new_n488), .B1(new_n502), .B2(new_n507), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n453), .B1(new_n460), .B2(new_n462), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT87), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n458), .A2(new_n450), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT87), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n509), .A2(new_n621), .A3(new_n622), .A4(new_n453), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n611), .A2(new_n613), .A3(new_n620), .A4(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n605), .A2(new_n608), .ZN(new_n625));
  INV_X1    g0425(.A(new_n583), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n551), .A2(new_n601), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n625), .B1(new_n627), .B2(KEYINPUT26), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT26), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n611), .A2(new_n629), .A3(new_n626), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n624), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n419), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n410), .A2(new_n369), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n414), .B1(new_n633), .B2(new_n366), .ZN(new_n634));
  INV_X1    g0434(.A(new_n318), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n635), .A2(new_n316), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n306), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n632), .A2(new_n638), .ZN(G369));
  NOR2_X1   g0439(.A1(new_n234), .A2(G20), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n269), .ZN(new_n641));
  OR2_X1    g0441(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(KEYINPUT27), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G213), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(G343), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n462), .A2(new_n647), .ZN(new_n648));
  MUX2_X1   g0448(.A(new_n468), .B(new_n619), .S(new_n648), .Z(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n511), .A2(new_n512), .B1(new_n489), .B2(new_n646), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n595), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n618), .A2(new_n646), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n458), .A2(KEYINPUT83), .A3(new_n450), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n461), .B1(new_n460), .B2(new_n462), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n657), .A2(new_n658), .B1(new_n452), .B2(new_n451), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n646), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI22_X1  g0461(.A1(new_n661), .A2(new_n652), .B1(new_n509), .B2(new_n646), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n656), .A2(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n236), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G1), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n226), .B2(new_n666), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT28), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n631), .A2(KEYINPUT90), .A3(new_n647), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT90), .B1(new_n631), .B2(new_n647), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT29), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT30), .ZN(new_n674));
  INV_X1    g0474(.A(new_n457), .ZN(new_n675));
  INV_X1    g0475(.A(new_n504), .ZN(new_n676));
  AOI211_X1 g0476(.A(new_n676), .B(new_n503), .C1(new_n548), .C2(new_n549), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT88), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n675), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n604), .A2(new_n678), .A3(new_n504), .A4(new_n494), .ZN(new_n680));
  INV_X1    g0480(.A(new_n560), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n674), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n681), .A2(new_n304), .A3(new_n506), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n606), .A2(KEYINPUT89), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n606), .A2(KEYINPUT89), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n684), .A2(new_n685), .A3(new_n439), .A4(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n504), .B(new_n494), .C1(new_n528), .C2(new_n531), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n457), .B1(new_n688), .B2(KEYINPUT88), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(KEYINPUT30), .A3(new_n681), .A4(new_n680), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n683), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(new_n646), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n468), .A2(new_n602), .A3(new_n513), .A4(new_n647), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT31), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(new_n695), .A3(new_n646), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n694), .A2(G330), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT29), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n627), .A2(new_n629), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT91), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n611), .A2(KEYINPUT26), .A3(new_n626), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n627), .A2(KEYINPUT91), .A3(new_n629), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n625), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n489), .A2(new_n508), .A3(KEYINPUT85), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT85), .B1(new_n489), .B2(new_n508), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(KEYINPUT92), .B1(new_n708), .B2(new_n464), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n596), .A2(new_n600), .A3(new_n610), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n595), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n584), .A2(KEYINPUT93), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT93), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n612), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n711), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT92), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n513), .A2(new_n716), .A3(new_n659), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n709), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n704), .A2(new_n705), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n698), .B1(new_n719), .B2(new_n647), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n673), .A2(new_n697), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n670), .B1(new_n721), .B2(G1), .ZN(G364));
  INV_X1    g0522(.A(new_n650), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n269), .B1(new_n640), .B2(G45), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n665), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(G330), .B2(new_n649), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n383), .A2(new_n384), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n664), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n227), .A2(new_n432), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n731), .B(new_n732), .C1(new_n259), .C2(new_n432), .ZN(new_n733));
  INV_X1    g0533(.A(G355), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n236), .A2(new_n261), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n733), .B1(G116), .B2(new_n236), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n228), .B1(G20), .B2(new_n282), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n726), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n229), .A2(new_n465), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n745), .A2(G179), .A3(G190), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n747), .A2(KEYINPUT94), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(KEYINPUT94), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n330), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n745), .A2(new_n303), .A3(new_n309), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n745), .A2(new_n303), .A3(G190), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n209), .A2(new_n753), .B1(new_n755), .B2(new_n201), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n751), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n229), .B1(new_n758), .B2(G190), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT95), .Z(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G97), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n303), .A2(G200), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(G20), .A3(G190), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n229), .A2(G190), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n764), .A2(new_n224), .B1(new_n766), .B2(new_n202), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n745), .A2(new_n309), .A3(G179), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n427), .B(new_n767), .C1(G87), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n765), .A2(new_n758), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n373), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT32), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n757), .A2(new_n762), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(G283), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT96), .ZN(new_n775));
  INV_X1    g0575(.A(new_n768), .ZN(new_n776));
  INV_X1    g0576(.A(G303), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n427), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n750), .A2(new_n774), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n775), .B2(new_n778), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n752), .A2(G326), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n759), .A2(new_n492), .ZN(new_n782));
  INV_X1    g0582(.A(new_n770), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G329), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n766), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT33), .B(G317), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n782), .B(new_n786), .C1(new_n754), .C2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n780), .A2(new_n781), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(G322), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n764), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n773), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n743), .B1(new_n792), .B2(new_n740), .ZN(new_n793));
  INV_X1    g0593(.A(new_n739), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n742), .B(new_n793), .C1(new_n649), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n728), .A2(new_n795), .ZN(G396));
  INV_X1    g0596(.A(new_n697), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT98), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n338), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n327), .A2(new_n337), .A3(KEYINPUT98), .A4(new_n336), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n799), .A2(new_n800), .B1(new_n415), .B2(new_n416), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n327), .A2(new_n646), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n801), .A2(new_n802), .B1(new_n339), .B2(new_n646), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n631), .A2(new_n647), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT90), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n631), .A2(KEYINPUT90), .A3(new_n647), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n631), .A2(new_n647), .A3(new_n801), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  OR3_X1    g0611(.A1(new_n797), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n743), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(KEYINPUT99), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n797), .B1(new_n809), .B2(new_n811), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT99), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n812), .A2(new_n816), .A3(new_n743), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n740), .A2(new_n737), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n202), .ZN(new_n820));
  INV_X1    g0620(.A(new_n750), .ZN(new_n821));
  INV_X1    g0621(.A(new_n764), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n821), .A2(G87), .B1(G294), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n427), .B1(new_n770), .B2(new_n785), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(new_n752), .B2(G303), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n823), .A2(new_n762), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n766), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n827), .A2(G116), .B1(G283), .B2(new_n754), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT97), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n826), .B(new_n829), .C1(new_n330), .C2(new_n776), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G137), .A2(new_n752), .B1(new_n754), .B2(G150), .ZN(new_n831));
  INV_X1    g0631(.A(G143), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n831), .B1(new_n832), .B2(new_n764), .C1(new_n373), .C2(new_n766), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n833), .B(KEYINPUT34), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n730), .B1(new_n224), .B2(new_n759), .C1(new_n835), .C2(new_n770), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n821), .B2(G68), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n834), .B(new_n837), .C1(new_n209), .C2(new_n776), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n830), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n743), .B1(new_n839), .B2(new_n740), .ZN(new_n840));
  OAI211_X1 g0640(.A(new_n820), .B(new_n840), .C1(new_n804), .C2(new_n738), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n818), .A2(new_n841), .ZN(G384));
  NAND2_X1  g0642(.A1(new_n566), .A2(new_n567), .ZN(new_n843));
  XOR2_X1   g0643(.A(new_n843), .B(KEYINPUT100), .Z(new_n844));
  INV_X1    g0644(.A(KEYINPUT35), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n846), .A2(G116), .A3(new_n230), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT101), .Z(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n845), .B2(new_n844), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT36), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n371), .A2(G77), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n226), .A2(new_n851), .B1(G50), .B2(new_n201), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(G1), .A3(new_n234), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT102), .Z(new_n855));
  INV_X1    g0655(.A(KEYINPUT104), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n409), .A2(KEYINPUT17), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n409), .A2(KEYINPUT17), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT18), .ZN(new_n859));
  AOI211_X1 g0659(.A(new_n859), .B(new_n412), .C1(new_n395), .C2(new_n397), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n395), .A2(new_n397), .ZN(new_n861));
  INV_X1    g0661(.A(new_n412), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT18), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI22_X1  g0663(.A1(new_n857), .A2(new_n858), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n644), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n409), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n395), .A2(new_n397), .B1(new_n412), .B2(new_n644), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n869), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT37), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(new_n872), .A3(new_n409), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n864), .A2(new_n867), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n856), .B1(new_n874), .B2(KEYINPUT38), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n377), .B1(new_n387), .B2(new_n201), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n389), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n295), .A3(new_n388), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n644), .B1(new_n878), .B2(new_n397), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n864), .A2(new_n879), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n878), .A2(new_n397), .B1(new_n412), .B2(new_n644), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n881), .B2(new_n868), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n873), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n866), .B1(new_n414), .B2(new_n410), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n870), .A2(new_n873), .ZN(new_n887));
  OAI211_X1 g0687(.A(KEYINPUT104), .B(new_n885), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n875), .A2(new_n884), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n353), .A2(new_n365), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n890), .B(new_n369), .C1(new_n364), .C2(new_n647), .ZN(new_n891));
  INV_X1    g0691(.A(new_n369), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n365), .B(new_n646), .C1(new_n892), .C2(new_n353), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n803), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n889), .A2(new_n694), .A3(new_n696), .A4(new_n894), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n694), .A2(new_n696), .A3(new_n894), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n880), .A2(KEYINPUT38), .A3(new_n883), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT38), .B1(new_n880), .B2(new_n883), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(KEYINPUT40), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n895), .A2(KEYINPUT40), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n694), .A2(new_n696), .ZN(new_n902));
  INV_X1    g0702(.A(new_n419), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n901), .B(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(G330), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT105), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n414), .A2(new_n865), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n875), .A2(new_n888), .A3(new_n909), .A4(new_n884), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT39), .B1(new_n897), .B2(new_n898), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n353), .A2(new_n365), .A3(new_n647), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n908), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n799), .A2(new_n647), .A3(new_n800), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT103), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n917), .A2(KEYINPUT103), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n810), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n891), .A2(new_n893), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n920), .B(new_n921), .C1(new_n897), .C2(new_n898), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n719), .A2(new_n647), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(KEYINPUT29), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n807), .A2(new_n698), .A3(new_n808), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n903), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n638), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n924), .B(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n907), .B(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n640), .A2(new_n269), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n855), .B1(new_n932), .B2(new_n933), .ZN(G367));
  AOI21_X1  g0734(.A(new_n730), .B1(G97), .B2(new_n746), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT46), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n768), .A2(G116), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n935), .B1(new_n936), .B2(new_n937), .C1(new_n330), .C2(new_n759), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n822), .A2(G303), .B1(G294), .B2(new_n754), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n939), .B1(new_n774), .B2(new_n766), .C1(new_n785), .C2(new_n753), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n937), .A2(new_n936), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT107), .Z(new_n942));
  NOR3_X1   g0742(.A1(new_n938), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(G317), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(new_n770), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n760), .A2(new_n201), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n427), .B1(new_n768), .B2(G58), .ZN(new_n947));
  INV_X1    g0747(.A(G137), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n947), .B1(new_n948), .B2(new_n770), .C1(new_n753), .C2(new_n832), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n946), .B(new_n949), .C1(G150), .C2(new_n822), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n755), .A2(new_n373), .B1(new_n209), .B2(new_n766), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT108), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n950), .B(new_n952), .C1(new_n202), .C2(new_n747), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n945), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT47), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n743), .B1(new_n955), .B2(new_n740), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n600), .A2(new_n647), .ZN(new_n957));
  MUX2_X1   g0757(.A(new_n611), .B(new_n625), .S(new_n957), .Z(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(new_n794), .ZN(new_n959));
  INV_X1    g0759(.A(new_n731), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n741), .B1(new_n236), .B2(new_n323), .C1(new_n248), .C2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n956), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n712), .A2(new_n714), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n581), .A2(new_n646), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n626), .A2(new_n646), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n662), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n662), .A2(new_n968), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT44), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n656), .ZN(new_n975));
  INV_X1    g0775(.A(new_n656), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n970), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OR3_X1    g0778(.A1(new_n654), .A2(KEYINPUT106), .A3(new_n660), .ZN(new_n979));
  INV_X1    g0779(.A(new_n652), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n660), .ZN(new_n981));
  OAI21_X1  g0781(.A(KEYINPUT106), .B1(new_n654), .B2(new_n660), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n979), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(new_n650), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n721), .B1(new_n978), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n665), .B(KEYINPUT41), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n725), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n981), .A2(KEYINPUT42), .A3(new_n965), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n583), .B1(new_n965), .B2(new_n513), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n647), .ZN(new_n990));
  OAI21_X1  g0790(.A(KEYINPUT42), .B1(new_n981), .B2(new_n965), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n656), .A2(new_n967), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n994));
  AND3_X1   g0794(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n993), .B1(new_n992), .B2(new_n994), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OR3_X1    g0798(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n998), .B1(new_n995), .B2(new_n996), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n962), .B1(new_n987), .B2(new_n1001), .ZN(G387));
  OAI22_X1  g0802(.A1(new_n764), .A2(new_n209), .B1(new_n766), .B2(new_n201), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n821), .B2(G97), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n760), .A2(new_n323), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G159), .B2(new_n752), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n754), .A2(new_n287), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n730), .B1(new_n285), .B2(new_n770), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G77), .B2(new_n768), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n822), .A2(G317), .B1(new_n827), .B2(G303), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n785), .B2(new_n755), .C1(new_n790), .C2(new_n753), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT48), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n776), .A2(new_n492), .B1(new_n759), .B2(new_n774), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT109), .Z(new_n1015));
  AND2_X1   g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT49), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(KEYINPUT49), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n730), .B1(G326), .B2(new_n783), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n747), .A2(new_n211), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1010), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n740), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1023), .B(new_n726), .C1(new_n654), .C2(new_n794), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n667), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n287), .A2(new_n209), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1025), .B1(new_n1026), .B2(KEYINPUT50), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1027), .A2(new_n1028), .A3(new_n432), .A4(new_n255), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n731), .B(new_n1029), .C1(new_n244), .C2(new_n432), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(G107), .B2(new_n236), .C1(new_n667), .C2(new_n735), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1024), .B1(new_n741), .B2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n983), .B(new_n723), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1032), .B1(new_n725), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n721), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n984), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1033), .A2(new_n721), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n665), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1034), .A2(new_n1038), .ZN(G393));
  INV_X1    g0839(.A(new_n977), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n976), .B1(new_n970), .B2(new_n973), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT110), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n725), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n261), .B1(new_n783), .B2(G322), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n211), .B2(new_n759), .C1(new_n776), .C2(new_n774), .ZN(new_n1046));
  AOI211_X1 g0846(.A(new_n1046), .B(new_n751), .C1(G294), .C2(new_n827), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n753), .A2(new_n944), .B1(new_n764), .B2(new_n785), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT52), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1047), .B(new_n1049), .C1(new_n777), .C2(new_n755), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n730), .B1(new_n832), .B2(new_n770), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n760), .A2(new_n202), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n287), .B2(new_n827), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n209), .B2(new_n755), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT111), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1051), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n821), .A2(G87), .B1(G68), .B2(new_n768), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n1055), .C2(new_n1054), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n822), .A2(G159), .B1(G150), .B2(new_n752), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT51), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1050), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n743), .B1(new_n1061), .B2(new_n740), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n741), .B1(new_n446), .B2(new_n236), .C1(new_n254), .C2(new_n960), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n794), .C2(new_n967), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n666), .B1(new_n978), .B2(new_n1037), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n978), .B2(new_n1037), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1044), .A2(new_n1064), .A3(new_n1066), .ZN(G390));
  NAND2_X1  g0867(.A1(new_n819), .A2(new_n288), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n427), .B1(new_n770), .B2(new_n492), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1069), .B(new_n1052), .C1(G87), .C2(new_n768), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n755), .A2(new_n330), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n753), .A2(new_n774), .B1(new_n446), .B2(new_n766), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1071), .B(new_n1072), .C1(G116), .C2(new_n822), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1070), .B(new_n1073), .C1(new_n201), .C2(new_n750), .ZN(new_n1074));
  XOR2_X1   g0874(.A(KEYINPUT54), .B(G143), .Z(new_n1075));
  AOI22_X1  g0875(.A1(new_n761), .A2(G159), .B1(new_n827), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n948), .B2(new_n755), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1077), .A2(KEYINPUT113), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(KEYINPUT113), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n764), .A2(new_n835), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n752), .A2(G128), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1081), .B(new_n261), .C1(new_n209), .C2(new_n747), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1080), .B(new_n1082), .C1(G125), .C2(new_n783), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1078), .A2(new_n1079), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n768), .A2(G150), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT114), .Z(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT53), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1074), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n743), .B1(new_n1088), .B2(new_n740), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1068), .B(new_n1089), .C1(new_n912), .C2(new_n738), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT115), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n921), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n719), .A2(new_n647), .A3(new_n801), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n916), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n889), .A2(new_n913), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n914), .B1(new_n920), .B2(new_n921), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1094), .A2(new_n1095), .B1(new_n1096), .B2(new_n912), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n694), .A2(new_n894), .A3(G330), .A4(new_n696), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1098), .B1(new_n1096), .B2(new_n912), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1091), .B1(new_n1102), .B2(new_n724), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT116), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n1091), .B(KEYINPUT116), .C1(new_n1102), .C2(new_n724), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n694), .A2(G330), .A3(new_n696), .A4(new_n804), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n1092), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1109), .A2(new_n916), .A3(new_n1093), .A4(new_n1098), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n920), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n697), .A2(new_n894), .B1(new_n1108), .B2(new_n1092), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(G330), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n902), .A2(new_n903), .A3(new_n1114), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n928), .A2(new_n929), .A3(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1113), .A2(new_n1116), .A3(KEYINPUT112), .ZN(new_n1117));
  AOI21_X1  g0917(.A(KEYINPUT112), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1102), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1100), .A2(new_n1113), .A3(new_n1101), .A4(new_n1116), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n665), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1107), .A2(new_n1121), .ZN(G378));
  INV_X1    g0922(.A(KEYINPUT118), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n302), .A2(new_n865), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n319), .A2(new_n1124), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n635), .A2(new_n316), .B1(new_n283), .B2(new_n305), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1124), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT55), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1125), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT56), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1129), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n319), .A2(new_n1124), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT55), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT56), .B1(new_n1137), .B2(new_n1130), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1123), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1138), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(KEYINPUT56), .A3(new_n1130), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(KEYINPUT118), .A3(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1139), .B(new_n1142), .C1(new_n901), .C2(new_n1114), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n895), .A2(KEYINPUT40), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n896), .A2(new_n900), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n1134), .A2(new_n1138), .A3(new_n1123), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1146), .A2(G330), .A3(new_n1147), .ZN(new_n1148));
  AND3_X1   g0948(.A1(new_n1143), .A2(new_n1148), .A3(new_n923), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n923), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n725), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1140), .A2(new_n737), .A3(new_n1141), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n819), .A2(new_n209), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n760), .A2(new_n285), .B1(new_n766), .B2(new_n948), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n822), .A2(G128), .B1(G125), .B2(new_n752), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n835), .B2(new_n755), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(new_n768), .C2(new_n1075), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1157), .B(KEYINPUT59), .ZN(new_n1158));
  AOI21_X1  g0958(.A(G41), .B1(new_n783), .B2(G124), .ZN(new_n1159));
  AOI21_X1  g0959(.A(G33), .B1(new_n746), .B2(G159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n275), .B1(new_n770), .B2(new_n774), .C1(new_n776), .C2(new_n202), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n730), .B(new_n1162), .C1(G58), .C2(new_n746), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n946), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n822), .A2(G107), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n755), .A2(new_n446), .B1(new_n323), .B2(new_n766), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G116), .B2(new_n752), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT58), .ZN(new_n1169));
  AOI21_X1  g0969(.A(G41), .B1(new_n730), .B2(G33), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1161), .B(new_n1169), .C1(G50), .C2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT117), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n743), .B1(new_n1172), .B2(new_n740), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1152), .A2(new_n1153), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1151), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1113), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1116), .B1(new_n1102), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n1150), .B2(new_n1149), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n666), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1143), .A2(new_n1148), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n924), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1143), .A2(new_n1148), .A3(new_n923), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1182), .A2(new_n1183), .B1(new_n1120), .B2(new_n1116), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(KEYINPUT57), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1175), .B1(new_n1180), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G375));
  OAI21_X1  g0987(.A(new_n730), .B1(new_n776), .B2(new_n373), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n746), .A2(G58), .B1(G128), .B2(new_n783), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n285), .B2(new_n766), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1188), .B(new_n1190), .C1(G50), .C2(new_n761), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT120), .Z(new_n1192));
  AOI22_X1  g0992(.A1(new_n822), .A2(G137), .B1(new_n754), .B2(new_n1075), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n835), .C2(new_n753), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n770), .A2(new_n777), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n750), .A2(new_n202), .B1(new_n330), .B2(new_n766), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G116), .B2(new_n754), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n427), .B1(new_n776), .B2(new_n446), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1198), .B(new_n1005), .C1(G294), .C2(new_n752), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1197), .B(new_n1199), .C1(new_n774), .C2(new_n764), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1194), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n743), .B1(new_n1201), .B2(new_n740), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n921), .B2(new_n738), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n201), .B2(new_n819), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1113), .B2(new_n725), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n986), .B(KEYINPUT119), .Z(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1205), .B1(new_n1207), .B2(new_n1208), .ZN(G381));
  INV_X1    g1009(.A(new_n1103), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1121), .A2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G375), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1034), .A2(new_n1038), .A3(new_n795), .A4(new_n728), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(G381), .A2(new_n1213), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(G390), .A2(G387), .A3(G384), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .ZN(G407));
  NAND2_X1  g1016(.A1(new_n645), .A2(G213), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1212), .A2(new_n1218), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT121), .Z(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(G213), .A3(G407), .ZN(G409));
  AND2_X1   g1021(.A1(new_n1151), .A2(new_n1174), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n665), .B1(new_n1184), .B2(KEYINPUT57), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1224));
  OAI211_X1 g1024(.A(G378), .B(new_n1222), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1184), .A2(new_n1206), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1121), .B(new_n1210), .C1(new_n1226), .C2(new_n1175), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT123), .ZN(new_n1229));
  XOR2_X1   g1029(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1229), .B1(new_n1231), .B2(new_n1208), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n419), .B1(new_n673), .B2(new_n720), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n904), .A2(G330), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n638), .A3(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1109), .A2(new_n1098), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(new_n920), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1237), .A3(new_n1110), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1235), .B1(new_n1237), .B2(new_n1110), .ZN(new_n1239));
  OAI211_X1 g1039(.A(KEYINPUT123), .B(new_n1238), .C1(new_n1239), .C2(new_n1230), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n666), .B1(new_n1208), .B2(KEYINPUT60), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1232), .A2(new_n1240), .A3(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1242), .A2(G384), .A3(new_n1205), .ZN(new_n1243));
  AOI21_X1  g1043(.A(G384), .B1(new_n1242), .B2(new_n1205), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1228), .A2(new_n1217), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT62), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1218), .A2(G2897), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1218), .A2(KEYINPUT125), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1245), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1242), .A2(new_n1205), .ZN(new_n1252));
  INV_X1    g1052(.A(G384), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1242), .A2(G384), .A3(new_n1205), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1254), .A2(new_n1249), .A3(new_n1255), .A4(new_n1250), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1211), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1184), .A2(new_n1206), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1222), .A2(new_n1259), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1186), .A2(G378), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1251), .A2(new_n1257), .B1(new_n1261), .B2(new_n1218), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT62), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1228), .A2(new_n1264), .A3(new_n1217), .A4(new_n1245), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1247), .A2(new_n1262), .A3(new_n1263), .A4(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(G390), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G393), .A2(G396), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1268), .A2(new_n1213), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT127), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1269), .B1(new_n1270), .B2(G387), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n962), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1035), .B1(new_n1042), .B2(new_n1033), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n986), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n724), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1001), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1272), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1268), .A2(new_n1213), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1267), .B1(new_n1271), .B2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1278), .B1(new_n1277), .B2(KEYINPUT127), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1269), .A2(G387), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1281), .A2(G390), .A3(new_n1282), .ZN(new_n1283));
  AND2_X1   g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1266), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(KEYINPUT61), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1228), .A2(KEYINPUT63), .A3(new_n1217), .A4(new_n1245), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1254), .A2(new_n1255), .A3(new_n1250), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1248), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n1256), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1228), .A2(new_n1217), .ZN(new_n1292));
  AND3_X1   g1092(.A1(new_n1291), .A2(KEYINPUT126), .A3(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(KEYINPUT126), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1288), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1246), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(KEYINPUT124), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT124), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1246), .A2(new_n1299), .A3(new_n1296), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1285), .B1(new_n1295), .B2(new_n1301), .ZN(G405));
  OAI21_X1  g1102(.A(new_n1225), .B1(new_n1186), .B2(new_n1211), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(new_n1303), .B(new_n1245), .ZN(new_n1304));
  XNOR2_X1  g1104(.A(new_n1304), .B(new_n1284), .ZN(G402));
endmodule


