//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT67), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  NOR3_X1   g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT69), .B1(new_n460), .B2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n464), .A2(new_n468), .B1(new_n473), .B2(G101), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G125), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n465), .A2(new_n466), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT70), .Z(G160));
  INV_X1    g056(.A(new_n464), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(new_n479), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT72), .Z(new_n485));
  OAI221_X1 g060(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n479), .C2(G112), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n482), .A2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  XOR2_X1   g064(.A(new_n489), .B(KEYINPUT71), .Z(new_n490));
  NAND2_X1  g065(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND2_X1  g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n465), .A2(new_n466), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n464), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n459), .A2(G2104), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n499), .A2(new_n500), .A3(G138), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT67), .B(G2105), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(G114), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n504), .B1(new_n505), .B2(G2105), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n497), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n511), .A2(G62), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT73), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n516), .A2(new_n521), .ZN(G166));
  XOR2_X1   g097(.A(KEYINPUT5), .B(G543), .Z(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT74), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n524), .A2(G63), .A3(G651), .ZN(new_n525));
  INV_X1    g100(.A(new_n514), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n512), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n525), .B(new_n527), .C1(KEYINPUT75), .C2(new_n531), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n531), .A2(KEYINPUT75), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n532), .A2(new_n533), .ZN(G168));
  AOI22_X1  g109(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n517), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  INV_X1    g112(.A(G52), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n512), .A2(new_n537), .B1(new_n514), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  AOI22_X1  g115(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n517), .ZN(new_n542));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n512), .A2(new_n543), .B1(new_n514), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g123(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n549));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n523), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n512), .ZN(new_n556));
  AOI22_X1  g131(.A1(G651), .A2(new_n555), .B1(new_n556), .B2(G91), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n510), .A2(G53), .A3(G543), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT9), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  INV_X1    g136(.A(G168), .ZN(G286));
  INV_X1    g137(.A(G166), .ZN(G303));
  NAND3_X1  g138(.A1(new_n556), .A2(KEYINPUT77), .A3(G87), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT77), .ZN(new_n565));
  INV_X1    g140(.A(G87), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n512), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n564), .A2(new_n567), .B1(G49), .B2(new_n526), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(G288));
  INV_X1    g145(.A(G86), .ZN(new_n571));
  INV_X1    g146(.A(G48), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n512), .A2(new_n571), .B1(new_n514), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n517), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(G85), .A2(new_n556), .B1(new_n526), .B2(G47), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n579), .B2(new_n517), .ZN(G290));
  AND3_X1   g155(.A1(new_n511), .A2(new_n510), .A3(G92), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n581), .B(KEYINPUT10), .ZN(new_n582));
  NAND2_X1  g157(.A1(G79), .A2(G543), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT78), .ZN(new_n584));
  INV_X1    g159(.A(G66), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n523), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(new_n526), .B2(G54), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n588), .A2(KEYINPUT79), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n588), .A2(KEYINPUT79), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  MUX2_X1   g167(.A(new_n592), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g168(.A(new_n592), .B(G301), .S(G868), .Z(G321));
  INV_X1    g169(.A(G299), .ZN(new_n595));
  OAI21_X1  g170(.A(KEYINPUT80), .B1(new_n595), .B2(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(G286), .A2(G868), .ZN(new_n597));
  MUX2_X1   g172(.A(KEYINPUT80), .B(new_n596), .S(new_n597), .Z(G297));
  MUX2_X1   g173(.A(KEYINPUT80), .B(new_n596), .S(new_n597), .Z(G280));
  XOR2_X1   g174(.A(KEYINPUT81), .B(G559), .Z(new_n600));
  OAI21_X1  g175(.A(new_n591), .B1(G860), .B2(new_n600), .ZN(G148));
  NAND2_X1  g176(.A1(new_n591), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(KEYINPUT82), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(KEYINPUT82), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n604), .B(new_n605), .C1(G868), .C2(new_n546), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AOI22_X1  g182(.A1(G123), .A2(new_n483), .B1(new_n488), .B2(G135), .ZN(new_n608));
  INV_X1    g183(.A(G111), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT84), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n502), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n610), .B2(new_n611), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(G2096), .Z(new_n615));
  NAND2_X1  g190(.A1(new_n473), .A2(new_n477), .ZN(new_n616));
  XNOR2_X1  g191(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT13), .Z(new_n619));
  INV_X1    g194(.A(G2100), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(new_n619), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(KEYINPUT85), .Z(G156));
  XOR2_X1   g198(.A(G1341), .B(G1348), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT89), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n625), .B(new_n626), .Z(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT88), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2430), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(KEYINPUT14), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n627), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT87), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G14), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n635), .A2(new_n639), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT90), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT17), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2084), .B(G2090), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n648), .B1(new_n645), .B2(new_n647), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n646), .B2(new_n647), .ZN(new_n651));
  INV_X1    g226(.A(new_n647), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n652), .A2(new_n648), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  NOR3_X1   g230(.A1(new_n649), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(new_n620), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT91), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n660));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT93), .ZN(new_n670));
  OR3_X1    g245(.A1(new_n662), .A2(new_n665), .A3(new_n668), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  INV_X1    g255(.A(G29), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G35), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G162), .B2(new_n681), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT29), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G2090), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT102), .Z(new_n686));
  XOR2_X1   g261(.A(KEYINPUT31), .B(G11), .Z(new_n687));
  XOR2_X1   g262(.A(KEYINPUT100), .B(G28), .Z(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(KEYINPUT30), .ZN(new_n689));
  AOI21_X1  g264(.A(G29), .B1(new_n688), .B2(KEYINPUT30), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n681), .A2(G32), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n488), .A2(G141), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n483), .A2(G129), .ZN(new_n694));
  NAND3_X1  g269(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT26), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n473), .A2(G105), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n693), .A2(new_n694), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n692), .B1(new_n698), .B2(G29), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT27), .B(G1996), .ZN(new_n700));
  OAI221_X1 g275(.A(new_n691), .B1(new_n681), .B2(new_n614), .C1(new_n699), .C2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n681), .A2(G33), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n703), .A2(new_n479), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT25), .ZN(new_n706));
  AOI211_X1 g281(.A(new_n704), .B(new_n706), .C1(G139), .C2(new_n488), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n702), .B1(new_n707), .B2(new_n681), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(G2072), .ZN(new_n709));
  NOR2_X1   g284(.A1(G27), .A2(G29), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G164), .B2(G29), .ZN(new_n711));
  AOI211_X1 g286(.A(new_n701), .B(new_n709), .C1(G2078), .C2(new_n711), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(G2078), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n699), .A2(new_n700), .ZN(new_n714));
  AOI211_X1 g289(.A(new_n713), .B(new_n714), .C1(G2072), .C2(new_n708), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G21), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G168), .B2(new_n716), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(G1966), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(KEYINPUT101), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(G4), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n591), .B2(new_n716), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G1348), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n712), .A2(new_n715), .A3(new_n720), .A4(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n546), .A2(new_n716), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n716), .B2(G19), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G171), .A2(new_n716), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G5), .B2(new_n716), .ZN(new_n729));
  INV_X1    g304(.A(G1961), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n727), .A2(G1341), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n681), .A2(G26), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT28), .Z(new_n733));
  OAI221_X1 g308(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n479), .C2(G116), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT98), .ZN(new_n735));
  AOI22_X1  g310(.A1(G128), .A2(new_n483), .B1(new_n488), .B2(G140), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n733), .B1(new_n737), .B2(G29), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT99), .B(G2067), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT24), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(G34), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(G34), .ZN(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G160), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(G29), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n740), .B1(G2084), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n731), .A2(new_n749), .ZN(new_n750));
  OAI22_X1  g325(.A1(new_n727), .A2(G1341), .B1(new_n729), .B2(new_n730), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n718), .A2(G1966), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n748), .B2(G2084), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n724), .A2(new_n750), .A3(new_n751), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n716), .A2(G20), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT23), .Z(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G299), .B2(G16), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT103), .ZN(new_n758));
  INV_X1    g333(.A(G1956), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI221_X1 g335(.A(new_n760), .B1(G1348), .B2(new_n722), .C1(KEYINPUT101), .C2(new_n719), .ZN(new_n761));
  INV_X1    g336(.A(new_n684), .ZN(new_n762));
  INV_X1    g337(.A(G2090), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND3_X1   g339(.A1(new_n686), .A2(new_n754), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(G16), .A2(G24), .ZN(new_n766));
  XOR2_X1   g341(.A(G290), .B(KEYINPUT94), .Z(new_n767));
  AOI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(G16), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT95), .ZN(new_n769));
  INV_X1    g344(.A(G1986), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n716), .A2(G23), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G288), .B2(G16), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT33), .B(G1976), .Z(new_n775));
  OR2_X1    g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n716), .A2(G22), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n716), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(G1971), .Z(new_n780));
  NOR2_X1   g355(.A1(G6), .A2(G16), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n576), .B2(G16), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT32), .B(G1981), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n776), .A2(new_n777), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(KEYINPUT34), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n681), .A2(G25), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n483), .A2(G119), .ZN(new_n788));
  OAI221_X1 g363(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n479), .C2(G107), .ZN(new_n789));
  AND2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n488), .A2(G131), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n787), .B1(new_n793), .B2(new_n681), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT35), .B(G1991), .Z(new_n795));
  XOR2_X1   g370(.A(new_n794), .B(new_n795), .Z(new_n796));
  AOI211_X1 g371(.A(KEYINPUT96), .B(new_n796), .C1(new_n785), .C2(KEYINPUT34), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n771), .A2(new_n786), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT97), .B(KEYINPUT36), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n765), .A2(new_n801), .ZN(G150));
  INV_X1    g377(.A(G150), .ZN(G311));
  NAND2_X1  g378(.A1(new_n524), .A2(G67), .ZN(new_n804));
  NAND2_X1  g379(.A1(G80), .A2(G543), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n517), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G93), .ZN(new_n807));
  INV_X1    g382(.A(G55), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n512), .A2(new_n807), .B1(new_n514), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G860), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT37), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n591), .A2(G559), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT38), .ZN(new_n815));
  INV_X1    g390(.A(new_n810), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n542), .B2(new_n545), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n546), .A2(new_n810), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n815), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT39), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT104), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n811), .B1(new_n820), .B2(new_n821), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n813), .B1(new_n823), .B2(new_n824), .ZN(G145));
  XNOR2_X1  g400(.A(new_n491), .B(G160), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(new_n614), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n737), .B(new_n508), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n698), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n707), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT105), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n792), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n488), .A2(G142), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n483), .A2(G130), .ZN(new_n834));
  OAI221_X1 g409(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n479), .C2(G118), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n832), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n618), .ZN(new_n838));
  INV_X1    g413(.A(new_n836), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n832), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n618), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n830), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n830), .A2(new_n843), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n827), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(KEYINPUT106), .B(G37), .ZN(new_n848));
  INV_X1    g423(.A(new_n827), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT107), .B1(new_n830), .B2(new_n843), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n849), .A2(new_n850), .A3(new_n844), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n830), .A2(KEYINPUT107), .A3(new_n843), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n847), .B(new_n848), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g429(.A1(new_n816), .A2(G868), .ZN(new_n855));
  XOR2_X1   g430(.A(G166), .B(KEYINPUT108), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G288), .ZN(new_n857));
  XNOR2_X1  g432(.A(G290), .B(new_n576), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT42), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n819), .B(new_n602), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n588), .B(G299), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT41), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n862), .B2(new_n861), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n860), .B1(new_n866), .B2(KEYINPUT109), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(KEYINPUT109), .B2(new_n866), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT109), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n860), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n855), .B1(new_n871), .B2(G868), .ZN(G295));
  AOI21_X1  g447(.A(new_n855), .B1(new_n871), .B2(G868), .ZN(G331));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n817), .A2(G301), .A3(new_n818), .ZN(new_n875));
  AOI21_X1  g450(.A(G301), .B1(new_n817), .B2(new_n818), .ZN(new_n876));
  OAI21_X1  g451(.A(G286), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n819), .A2(G171), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n817), .A2(G301), .A3(new_n818), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(G168), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n877), .A2(new_n880), .A3(new_n863), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n862), .B1(new_n877), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n859), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n859), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n877), .A2(new_n880), .A3(new_n863), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n877), .A2(new_n880), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n884), .B(new_n885), .C1(new_n886), .C2(new_n862), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n883), .A2(new_n887), .A3(new_n888), .A4(new_n848), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT110), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n883), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT43), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n889), .A2(KEYINPUT110), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n874), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n892), .A2(new_n888), .ZN(new_n897));
  AND4_X1   g472(.A1(KEYINPUT43), .A2(new_n883), .A3(new_n887), .A4(new_n848), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT44), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(G397));
  INV_X1    g475(.A(G1384), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n508), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT112), .ZN(new_n906));
  XNOR2_X1  g481(.A(KEYINPUT111), .B(G40), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n478), .B2(new_n479), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n468), .A2(new_n464), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n473), .A2(G101), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n906), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n499), .A2(new_n500), .A3(G125), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n475), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n907), .B1(new_n915), .B2(new_n502), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(KEYINPUT112), .A3(new_n474), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n905), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G1996), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT46), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n737), .A2(G2067), .ZN(new_n924));
  INV_X1    g499(.A(G2067), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n735), .A2(new_n925), .A3(new_n736), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n920), .B1(new_n928), .B2(new_n698), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n923), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT47), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n698), .B(new_n921), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n793), .A2(new_n795), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n926), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n920), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n792), .B(new_n795), .Z(new_n937));
  NOR2_X1   g512(.A1(new_n933), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n938), .A2(new_n919), .ZN(new_n939));
  XOR2_X1   g514(.A(new_n939), .B(KEYINPUT126), .Z(new_n940));
  NOR3_X1   g515(.A1(new_n919), .A2(G1986), .A3(G290), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT48), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n931), .B(new_n936), .C1(new_n940), .C2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G8), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n495), .B1(new_n502), .B2(new_n493), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n506), .B1(new_n946), .B2(new_n464), .ZN(new_n947));
  AOI21_X1  g522(.A(G1384), .B1(new_n947), .B2(new_n503), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n945), .B1(new_n918), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G1981), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n576), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT49), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n576), .A2(new_n950), .ZN(new_n954));
  OR3_X1    g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n953), .B1(new_n952), .B2(new_n954), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n949), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(G288), .A2(G1976), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n949), .B1(new_n959), .B2(new_n952), .ZN(new_n960));
  AOI21_X1  g535(.A(G1976), .B1(new_n568), .B2(new_n569), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT115), .ZN(new_n962));
  OR3_X1    g537(.A1(new_n961), .A2(new_n962), .A3(KEYINPUT52), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n962), .B1(new_n961), .B2(KEYINPUT52), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n568), .A2(new_n569), .A3(G1976), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n963), .A2(new_n964), .A3(new_n949), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n949), .A2(new_n965), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT52), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n966), .A2(new_n968), .A3(new_n957), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(G303), .A2(G8), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT55), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  XOR2_X1   g548(.A(KEYINPUT113), .B(G1971), .Z(new_n974));
  AND2_X1   g549(.A1(new_n918), .A2(new_n904), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n902), .A2(new_n903), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n974), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n902), .A2(KEYINPUT50), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n508), .A2(new_n980), .A3(new_n901), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n918), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n763), .A2(KEYINPUT114), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n763), .A2(KEYINPUT114), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n973), .B(G8), .C1(new_n978), .C2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n960), .B1(new_n970), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT117), .ZN(new_n988));
  OAI21_X1  g563(.A(G8), .B1(new_n985), .B2(new_n978), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n972), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n969), .A2(new_n990), .A3(new_n986), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n975), .A2(KEYINPUT116), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n918), .A2(new_n904), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT116), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n976), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(G1966), .B1(new_n992), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n982), .A2(G2084), .ZN(new_n997));
  OAI211_X1 g572(.A(G8), .B(G168), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n991), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n988), .B1(new_n999), .B2(KEYINPUT63), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT63), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n991), .B2(new_n998), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n987), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n992), .A2(new_n995), .ZN(new_n1004));
  INV_X1    g579(.A(G1966), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n997), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n945), .B1(new_n1006), .B2(G168), .ZN(new_n1007));
  OAI21_X1  g582(.A(G286), .B1(new_n996), .B2(new_n997), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT51), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT62), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1013), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1012), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT62), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n975), .A2(new_n977), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1018), .B1(new_n1019), .B2(G2078), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n982), .A2(KEYINPUT120), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n917), .A2(new_n913), .B1(new_n902), .B2(KEYINPUT50), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(new_n981), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1018), .A2(G2078), .ZN(new_n1026));
  OAI221_X1 g601(.A(new_n1020), .B1(new_n1025), .B2(G1961), .C1(new_n1004), .C2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(G171), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n991), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1014), .A2(new_n1017), .A3(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n988), .B(new_n1001), .C1(new_n991), .C2(new_n998), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1003), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1023), .B1(new_n1022), .B2(new_n981), .ZN(new_n1033));
  AND4_X1   g608(.A1(new_n1023), .A2(new_n918), .A3(new_n979), .A4(new_n981), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G1348), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n916), .A2(KEYINPUT112), .A3(new_n474), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT112), .B1(new_n916), .B2(new_n474), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1037), .B(new_n948), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1037), .B1(new_n918), .B2(new_n948), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n925), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1035), .A2(new_n1036), .B1(new_n1043), .B2(KEYINPUT119), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n948), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT118), .ZN(new_n1046));
  AOI21_X1  g621(.A(G2067), .B1(new_n1046), .B2(new_n1040), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT121), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1043), .A2(KEYINPUT119), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1021), .A2(new_n1024), .A3(new_n1036), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1051), .A2(new_n1049), .A3(KEYINPUT121), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT60), .B1(new_n1050), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(KEYINPUT124), .A3(new_n592), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1052), .B1(new_n1048), .B2(new_n1047), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1043), .A2(KEYINPUT119), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT60), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(new_n1053), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1061), .B1(new_n1060), .B2(new_n1053), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT124), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n591), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g640(.A(KEYINPUT124), .B(new_n1061), .C1(new_n1060), .C2(new_n1053), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1056), .B(new_n1062), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n975), .A2(new_n977), .A3(new_n1068), .ZN(new_n1069));
  AND2_X1   g644(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1070));
  NOR2_X1   g645(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n982), .A2(new_n759), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT61), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1076), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT61), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n1074), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT58), .B(G1341), .Z(new_n1081));
  NAND3_X1  g656(.A1(new_n1046), .A2(new_n1040), .A3(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n977), .A2(new_n921), .A3(new_n918), .A4(new_n904), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1082), .A2(KEYINPUT122), .A3(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT122), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n546), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT59), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1088), .B(new_n546), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1089));
  AOI221_X4 g664(.A(KEYINPUT123), .B1(new_n1077), .B2(new_n1080), .C1(new_n1087), .C2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1067), .A2(new_n1095), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1050), .A2(new_n1054), .A3(new_n592), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1074), .B1(new_n1097), .B2(new_n1076), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1100));
  INV_X1    g675(.A(G40), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n480), .A2(new_n1101), .A3(new_n1026), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n977), .A2(new_n904), .A3(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1020), .B(new_n1103), .C1(new_n1025), .C2(G1961), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1028), .B1(G171), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1027), .A2(G171), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1106), .B1(new_n1104), .B2(G171), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n991), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1100), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1100), .A2(new_n1107), .A3(new_n1110), .A4(KEYINPUT125), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1032), .B1(new_n1099), .B2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(G290), .B(new_n770), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n919), .B1(new_n938), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n944), .B1(new_n1116), .B2(new_n1118), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n1121));
  OAI21_X1  g695(.A(G319), .B1(new_n641), .B2(new_n642), .ZN(new_n1122));
  NOR2_X1   g696(.A1(G227), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g697(.A(KEYINPUT127), .B1(new_n679), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g698(.A1(new_n679), .A2(KEYINPUT127), .A3(new_n1123), .ZN(new_n1125));
  OAI21_X1  g699(.A(new_n853), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g700(.A1(new_n1121), .A2(new_n1126), .ZN(G308));
  OAI221_X1 g701(.A(new_n853), .B1(new_n1124), .B2(new_n1125), .C1(new_n894), .C2(new_n895), .ZN(G225));
endmodule


