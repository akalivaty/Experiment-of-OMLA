//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI21_X1  g031(.A(KEYINPUT65), .B1(new_n452), .B2(G2106), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n457), .B1(G567), .B2(new_n454), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n452), .A2(KEYINPUT65), .A3(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT66), .Z(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n465), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n472), .A2(KEYINPUT3), .A3(new_n473), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n477), .A2(G137), .A3(new_n478), .A4(new_n464), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n478), .A3(new_n464), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n477), .A2(G2105), .A3(new_n464), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n478), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND4_X1  g065(.A1(new_n477), .A2(KEYINPUT4), .A3(G138), .A4(new_n464), .ZN(new_n491));
  NAND2_X1  g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n477), .A2(G126), .A3(new_n464), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n478), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n467), .ZN(new_n497));
  AND2_X1   g072(.A1(new_n478), .A2(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT4), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n493), .A2(new_n496), .A3(new_n499), .ZN(G164));
  OR2_X1    g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  XOR2_X1   g091(.A(KEYINPUT68), .B(G88), .Z(new_n517));
  OAI22_X1  g092(.A1(new_n510), .A2(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n506), .A2(new_n518), .ZN(G166));
  NAND3_X1  g094(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT69), .ZN(new_n521));
  INV_X1    g096(.A(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(new_n507), .B2(new_n508), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G51), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(new_n516), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n521), .B(new_n524), .C1(new_n525), .C2(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n529), .A2(new_n525), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n505), .ZN(new_n534));
  INV_X1    g109(.A(G52), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n510), .A2(new_n535), .B1(new_n516), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n505), .ZN(new_n540));
  INV_X1    g115(.A(new_n516), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n541), .A2(G81), .B1(G43), .B2(new_n523), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT71), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n523), .A2(new_n551), .A3(G53), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT9), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n503), .A2(G65), .ZN(new_n554));
  INV_X1    g129(.A(G78), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT74), .B1(new_n555), .B2(new_n522), .ZN(new_n556));
  OR3_X1    g131(.A1(new_n555), .A2(new_n522), .A3(KEYINPUT74), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT73), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n503), .A2(new_n509), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G91), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n560), .A2(new_n565), .ZN(G299));
  XNOR2_X1  g141(.A(G171), .B(KEYINPUT75), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  OR2_X1    g145(.A1(new_n503), .A2(G74), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(new_n523), .B2(G49), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n561), .A2(G87), .A3(new_n563), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G288));
  OAI21_X1  g149(.A(G61), .B1(new_n513), .B2(new_n512), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(KEYINPUT76), .A2(G73), .A3(G543), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(G48), .B2(new_n523), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n561), .A2(G86), .A3(new_n563), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n541), .A2(G85), .B1(G47), .B2(new_n523), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n584), .A2(KEYINPUT77), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n584), .A2(KEYINPUT77), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n585), .A2(new_n586), .B1(new_n505), .B2(new_n587), .ZN(G290));
  XNOR2_X1  g163(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n564), .A2(G92), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n503), .A2(G66), .ZN(new_n592));
  INV_X1    g167(.A(G79), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n522), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(G54), .B2(new_n523), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n590), .B1(new_n564), .B2(G92), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  MUX2_X1   g175(.A(G301), .B(new_n599), .S(new_n600), .Z(G321));
  XNOR2_X1  g176(.A(G321), .B(KEYINPUT79), .ZN(G284));
  NAND2_X1  g177(.A1(G299), .A2(new_n600), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n600), .B2(G168), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(new_n600), .B2(G168), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n606), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT80), .ZN(new_n609));
  MUX2_X1   g184(.A(new_n543), .B(new_n609), .S(G868), .Z(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n485), .A2(G123), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n478), .A2(G111), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n483), .A2(G135), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n615), .A2(KEYINPUT82), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n615), .A2(KEYINPUT82), .ZN(new_n617));
  OAI221_X1 g192(.A(new_n612), .B1(new_n613), .B2(new_n614), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND2_X1  g194(.A1(new_n497), .A2(new_n474), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n619), .A2(new_n624), .ZN(G156));
  XOR2_X1   g200(.A(KEYINPUT15), .B(G2435), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2438), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2430), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT84), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n627), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n630), .A2(KEYINPUT14), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G1341), .B(G1348), .Z(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n632), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2451), .B(G2454), .Z(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n636), .A2(new_n639), .ZN(new_n641));
  AND3_X1   g216(.A1(new_n640), .A2(G14), .A3(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT18), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(KEYINPUT17), .ZN(new_n649));
  INV_X1    g224(.A(new_n643), .ZN(new_n650));
  INV_X1    g225(.A(new_n644), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n650), .A2(new_n646), .A3(new_n651), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(new_n645), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n648), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2096), .B(G2100), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n664), .A2(new_n662), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n659), .A2(new_n664), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n667));
  OAI221_X1 g242(.A(new_n663), .B1(new_n665), .B2(new_n659), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  AOI21_X1  g243(.A(new_n668), .B1(new_n666), .B2(new_n667), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1991), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1981), .B(G1986), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G229));
  AND2_X1   g250(.A1(new_n572), .A2(new_n573), .ZN(new_n676));
  INV_X1    g251(.A(G16), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n677), .B2(G23), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT33), .B(G1976), .Z(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  MUX2_X1   g257(.A(G6), .B(G305), .S(G16), .Z(new_n683));
  XOR2_X1   g258(.A(KEYINPUT32), .B(G1981), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n677), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n677), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(G1971), .Z(new_n689));
  NAND4_X1  g264(.A1(new_n682), .A2(new_n685), .A3(new_n686), .A4(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT34), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(KEYINPUT34), .ZN(new_n692));
  MUX2_X1   g267(.A(G24), .B(G290), .S(G16), .Z(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(G1986), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n483), .A2(G131), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n485), .A2(G119), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n478), .A2(G107), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n695), .B(new_n696), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G29), .ZN(new_n700));
  INV_X1    g275(.A(G29), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G25), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT86), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT35), .B(G1991), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n691), .A2(new_n692), .A3(new_n694), .A4(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT36), .Z(new_n708));
  INV_X1    g283(.A(G1956), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n677), .A2(G20), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT95), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT23), .ZN(new_n712));
  INV_X1    g287(.A(G299), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n677), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G168), .A2(new_n677), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n677), .B2(G21), .ZN(new_n717));
  INV_X1    g292(.A(G1966), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n709), .A2(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n709), .B2(new_n715), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n701), .A2(G32), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n483), .A2(G141), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT91), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT26), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n474), .A2(G105), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G129), .B2(new_n485), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n721), .B1(new_n730), .B2(new_n701), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT27), .B(G1996), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT25), .Z(new_n735));
  INV_X1    g310(.A(G139), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n497), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n735), .B1(new_n736), .B2(new_n482), .C1(new_n737), .C2(new_n478), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT89), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  MUX2_X1   g315(.A(G33), .B(new_n740), .S(G29), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2072), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n701), .A2(G26), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT28), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n483), .A2(G140), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n485), .A2(G128), .ZN(new_n746));
  OR2_X1    g321(.A1(G104), .A2(G2105), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n747), .B(G2104), .C1(G116), .C2(new_n478), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n745), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n744), .B1(new_n750), .B2(new_n701), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT88), .B(G2067), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n733), .A2(new_n742), .A3(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G34), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n755), .B2(KEYINPUT24), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(KEYINPUT24), .B2(new_n755), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n480), .B2(new_n701), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G2084), .ZN(new_n759));
  NOR2_X1   g334(.A1(G5), .A2(G16), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT92), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G171), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1961), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n759), .B(new_n764), .C1(new_n701), .C2(new_n618), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT31), .B(G11), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT30), .B(G28), .Z(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(G29), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n544), .A2(G16), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G16), .B2(G19), .ZN(new_n770));
  INV_X1    g345(.A(G1341), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n772), .B1(new_n771), .B2(new_n770), .C1(new_n717), .C2(new_n718), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n720), .A2(new_n754), .A3(new_n765), .A4(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n741), .A2(G2072), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT90), .ZN(new_n777));
  NOR2_X1   g352(.A1(G29), .A2(G35), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G162), .B2(G29), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G2090), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT94), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n677), .A2(G4), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n598), .B2(new_n677), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT87), .B(G1348), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n701), .A2(G27), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G164), .B2(new_n701), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2078), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n781), .B2(G2090), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n783), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  NOR4_X1   g367(.A1(new_n708), .A2(new_n775), .A3(new_n777), .A4(new_n792), .ZN(G311));
  INV_X1    g368(.A(G311), .ZN(G150));
  NAND2_X1  g369(.A1(new_n598), .A2(G559), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT38), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n797), .A2(new_n505), .ZN(new_n798));
  INV_X1    g373(.A(G55), .ZN(new_n799));
  INV_X1    g374(.A(G93), .ZN(new_n800));
  OAI22_X1  g375(.A1(new_n510), .A2(new_n799), .B1(new_n516), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n543), .B(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n796), .B(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(KEYINPUT39), .ZN(new_n805));
  INV_X1    g380(.A(G860), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(KEYINPUT39), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n805), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n802), .A2(new_n806), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT37), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(G145));
  XNOR2_X1  g386(.A(new_n740), .B(new_n729), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n699), .B(new_n622), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n494), .A2(new_n495), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n499), .B1(new_n815), .B2(G2105), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n491), .A2(new_n492), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(new_n478), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(new_n749), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n483), .A2(G142), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n485), .A2(G130), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n478), .A2(G118), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n821), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n820), .B(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n814), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n480), .B(new_n489), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(new_n618), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n814), .A2(new_n826), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n827), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(G37), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n829), .B1(new_n827), .B2(new_n830), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT96), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n827), .A2(new_n830), .ZN(new_n836));
  INV_X1    g411(.A(new_n829), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT96), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n838), .A2(new_n839), .A3(new_n832), .A4(new_n831), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g417(.A1(new_n713), .A2(new_n598), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n599), .A2(G299), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT98), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT41), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n843), .A2(new_n844), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT98), .B1(new_n849), .B2(KEYINPUT41), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n609), .B(new_n803), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT99), .B(KEYINPUT41), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n849), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT100), .B1(new_n845), .B2(new_n854), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n851), .A2(new_n852), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n845), .A2(KEYINPUT97), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n845), .A2(KEYINPUT97), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n858), .B1(new_n862), .B2(new_n852), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n676), .B(KEYINPUT101), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(G290), .ZN(new_n865));
  XNOR2_X1  g440(.A(G305), .B(G166), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(KEYINPUT102), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n866), .B(KEYINPUT102), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT42), .ZN(new_n870));
  OAI21_X1  g445(.A(G868), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(new_n870), .B2(new_n863), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n874), .B(new_n875), .C1(G868), .C2(new_n802), .ZN(G295));
  OAI211_X1 g451(.A(new_n874), .B(new_n875), .C1(G868), .C2(new_n802), .ZN(G331));
  NAND2_X1  g452(.A1(G168), .A2(new_n567), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(G168), .B2(G171), .ZN(new_n879));
  INV_X1    g454(.A(new_n803), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n878), .B(new_n803), .C1(G168), .C2(G171), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(KEYINPUT104), .A3(new_n880), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n845), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n857), .A2(new_n848), .A3(new_n856), .A4(new_n850), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n881), .A2(new_n883), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n886), .A2(KEYINPUT105), .A3(new_n845), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n869), .ZN(new_n895));
  INV_X1    g470(.A(new_n869), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n889), .A2(new_n892), .A3(new_n896), .A4(new_n893), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n895), .A2(new_n832), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n849), .A2(new_n847), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n849), .B2(new_n854), .ZN(new_n903));
  OAI22_X1  g478(.A1(new_n861), .A2(new_n891), .B1(new_n886), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n904), .B2(new_n869), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n899), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT106), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n898), .A2(KEYINPUT43), .B1(new_n901), .B2(new_n905), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n910), .A2(new_n911), .A3(KEYINPUT44), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n900), .B1(new_n905), .B2(new_n897), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n901), .A2(new_n832), .A3(new_n895), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT44), .ZN(new_n915));
  OAI22_X1  g490(.A1(new_n909), .A2(new_n912), .B1(new_n913), .B2(new_n915), .ZN(G397));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(G164), .B2(G1384), .ZN(new_n918));
  AND4_X1   g493(.A1(G40), .A2(new_n470), .A3(new_n479), .A4(new_n475), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G1996), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n729), .B(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G2067), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n749), .B(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n705), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n699), .A2(new_n926), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n923), .A2(new_n925), .A3(new_n927), .A4(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(G290), .B(G1986), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n921), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n932), .B(KEYINPUT107), .Z(new_n933));
  INV_X1    g508(.A(KEYINPUT118), .ZN(new_n934));
  INV_X1    g509(.A(G1384), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n819), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n816), .B2(new_n818), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n936), .A2(KEYINPUT50), .B1(new_n939), .B2(KEYINPUT109), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n819), .A2(new_n937), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n920), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G2084), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n819), .A2(KEYINPUT45), .A3(new_n935), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n918), .A2(new_n919), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n718), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(new_n948), .A3(G168), .ZN(new_n949));
  AND2_X1   g524(.A1(KEYINPUT51), .A2(G8), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(G168), .B1(new_n945), .B2(new_n948), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT51), .B1(new_n949), .B2(G8), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n934), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n954), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n945), .A2(new_n948), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(G286), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n958), .A2(new_n949), .A3(new_n950), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n959), .A3(KEYINPUT118), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n955), .A2(KEYINPUT62), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT123), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT123), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n955), .A2(new_n960), .A3(new_n963), .A4(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT62), .B1(new_n955), .B2(new_n960), .ZN(new_n966));
  XOR2_X1   g541(.A(KEYINPUT112), .B(G1981), .Z(new_n967));
  NAND3_X1  g542(.A1(new_n581), .A2(new_n582), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G61), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n969), .B1(new_n501), .B2(new_n502), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n578), .A2(new_n579), .ZN(new_n971));
  OAI21_X1  g546(.A(G651), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n523), .A2(G48), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n503), .A2(new_n509), .A3(G86), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G1981), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n968), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT49), .ZN(new_n980));
  INV_X1    g555(.A(G8), .ZN(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n816), .B2(new_n818), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(new_n982), .B2(new_n919), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT49), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n977), .A2(new_n978), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n980), .A2(new_n983), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n819), .A2(new_n919), .A3(new_n935), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n676), .A2(G1976), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(G8), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT52), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(G288), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n983), .A2(new_n988), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n986), .A2(new_n990), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT115), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n986), .A2(new_n990), .A3(new_n996), .A4(new_n993), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n999));
  NAND3_X1  g574(.A1(G303), .A2(G8), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n999), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(G166), .B2(new_n981), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n941), .A2(new_n919), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n982), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G2090), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT108), .B(G1971), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1007), .A2(new_n1008), .B1(new_n947), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1003), .B1(new_n1010), .B2(new_n981), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n940), .A2(new_n943), .A3(new_n1008), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n947), .A2(new_n1009), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1003), .B(KEYINPUT111), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(G8), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n998), .A2(new_n1011), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n947), .B2(G2078), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n940), .A2(new_n943), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n763), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n918), .A2(new_n946), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1018), .A2(G2078), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n919), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1025), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1019), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1017), .A2(new_n567), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n966), .A2(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n965), .A2(KEYINPUT124), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT124), .B1(new_n965), .B2(new_n1030), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1014), .A2(G8), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1003), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G286), .A2(new_n981), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n957), .A2(KEYINPUT63), .A3(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1035), .A2(new_n1016), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n994), .B(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n957), .A2(new_n1036), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n998), .A2(new_n1011), .A3(new_n1016), .A4(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT63), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1038), .A2(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1016), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n986), .A2(new_n991), .A3(new_n676), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n968), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n983), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1033), .B1(new_n1044), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1040), .A2(new_n1037), .A3(new_n1016), .A4(new_n1035), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1050), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(new_n1055), .A3(KEYINPUT116), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n987), .A2(G2067), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(new_n1020), .B2(new_n786), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(new_n599), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT57), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1060), .B1(new_n560), .B2(new_n565), .ZN(new_n1061));
  AND4_X1   g636(.A1(new_n1060), .A2(new_n553), .A3(new_n565), .A4(new_n559), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n709), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT56), .B(G2072), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n918), .A2(new_n946), .A3(new_n919), .A4(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1059), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1063), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1070), .B2(new_n1069), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1067), .A2(KEYINPUT61), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1058), .A2(KEYINPUT60), .A3(new_n599), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT58), .B(G1341), .Z(new_n1076));
  NAND2_X1  g651(.A1(new_n987), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n947), .B2(G1996), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n544), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(KEYINPUT59), .A3(new_n544), .ZN(new_n1082));
  AND4_X1   g657(.A1(new_n1074), .A2(new_n1075), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n1058), .A2(KEYINPUT60), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n599), .B1(new_n1058), .B2(KEYINPUT60), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1063), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1069), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n1067), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT61), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1084), .A2(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1073), .B1(new_n1083), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n955), .A2(new_n1017), .A3(new_n960), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(G301), .B(new_n1019), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n920), .A2(KEYINPUT120), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n920), .A2(KEYINPUT120), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1022), .A2(new_n1023), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1021), .A2(new_n1097), .A3(new_n1019), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G171), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1094), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT54), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1028), .A2(new_n567), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1098), .A2(new_n567), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(KEYINPUT54), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1104), .A2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1051), .A2(new_n1056), .B1(new_n1093), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n1031), .A2(new_n1032), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1093), .A2(new_n1109), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n933), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n921), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(new_n730), .B2(new_n925), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT46), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n921), .A2(new_n922), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT47), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n923), .A2(new_n925), .A3(new_n928), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n750), .A2(new_n924), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1118), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  OR3_X1    g702(.A1(new_n1118), .A2(G1986), .A3(G290), .ZN(new_n1128));
  XNOR2_X1  g703(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n921), .A2(new_n930), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  OR2_X1    g705(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1127), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1124), .A2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT126), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1117), .A2(new_n1134), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g710(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1137));
  NAND2_X1  g711(.A1(new_n841), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g712(.A(KEYINPUT127), .B1(new_n1138), .B2(new_n910), .ZN(new_n1139));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n1140));
  NAND4_X1  g714(.A1(new_n907), .A2(new_n1140), .A3(new_n841), .A4(new_n1137), .ZN(new_n1141));
  AND2_X1   g715(.A1(new_n1139), .A2(new_n1141), .ZN(G308));
  NAND3_X1  g716(.A1(new_n907), .A2(new_n841), .A3(new_n1137), .ZN(G225));
endmodule


