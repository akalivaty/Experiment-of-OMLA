//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G131), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT66), .A2(G134), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT66), .A2(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G137), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n188), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT11), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n189), .A2(G137), .A3(new_n190), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n194), .A2(G137), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT11), .B1(new_n191), .B2(new_n192), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT67), .B(G131), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n196), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT65), .A2(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(G143), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT68), .A2(G128), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT68), .A2(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT64), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(KEYINPUT64), .A2(G143), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n207), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  INV_X1    g034(.A(new_n209), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT65), .A2(G146), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n211), .A2(new_n215), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n220), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(G146), .A3(new_n216), .ZN(new_n228));
  AND4_X1   g042(.A1(new_n225), .A2(new_n210), .A3(new_n228), .A4(G128), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT69), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n210), .A2(new_n228), .A3(new_n225), .A4(G128), .ZN(new_n232));
  AOI21_X1  g046(.A(G146), .B1(new_n227), .B2(new_n216), .ZN(new_n233));
  AOI21_X1  g047(.A(G143), .B1(new_n208), .B2(new_n209), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n214), .B1(new_n210), .B2(KEYINPUT1), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n231), .B(new_n232), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n205), .A2(new_n230), .A3(new_n237), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT2), .B(G113), .Z(new_n239));
  XNOR2_X1  g053(.A(G116), .B(G119), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n239), .A2(new_n240), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(G131), .B1(new_n201), .B2(new_n202), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT66), .A2(G134), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT66), .A2(G134), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n197), .B1(new_n247), .B2(G137), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n199), .B1(new_n247), .B2(G137), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n204), .B(new_n248), .C1(new_n249), .C2(new_n197), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n244), .A2(new_n250), .ZN(new_n251));
  AND2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n233), .B2(new_n234), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n210), .A2(new_n228), .A3(new_n252), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n238), .A2(new_n243), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G237), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(KEYINPUT27), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G101), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n238), .A2(KEYINPUT30), .A3(new_n259), .ZN(new_n268));
  INV_X1    g082(.A(new_n243), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n232), .B1(new_n235), .B2(new_n236), .ZN(new_n271));
  INV_X1    g085(.A(new_n196), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n271), .A2(new_n250), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n257), .B1(new_n250), .B2(new_n244), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n268), .A2(new_n269), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT70), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n268), .A2(new_n275), .A3(new_n278), .A4(new_n269), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n267), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT31), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n238), .A2(new_n243), .A3(new_n259), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT28), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n260), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n266), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n277), .A2(new_n279), .ZN(new_n292));
  INV_X1    g106(.A(new_n267), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n281), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n187), .B1(new_n291), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT32), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n280), .A2(new_n281), .B1(new_n289), .B2(new_n288), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n293), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT31), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT32), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(new_n301), .A3(new_n187), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n243), .B1(new_n238), .B2(new_n259), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT28), .B1(new_n283), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT71), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n238), .A2(new_n259), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n269), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n260), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT28), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n266), .A2(KEYINPUT29), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n306), .A2(new_n311), .A3(new_n287), .A4(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(KEYINPUT72), .A3(new_n314), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n288), .A2(new_n289), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n319), .A2(KEYINPUT29), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n292), .A2(new_n260), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n289), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n317), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G472), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n303), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(G221), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT9), .B(G234), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n327), .B1(new_n329), .B2(new_n314), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT10), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT81), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n210), .A2(new_n228), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G128), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(new_n219), .B2(KEYINPUT1), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n232), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G107), .ZN(new_n338));
  AND2_X1   g152(.A1(KEYINPUT80), .A2(G104), .ZN(new_n339));
  NOR2_X1   g153(.A1(KEYINPUT80), .A2(G104), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n342));
  INV_X1    g156(.A(G101), .ZN(new_n343));
  OR2_X1    g157(.A1(KEYINPUT80), .A2(G104), .ZN(new_n344));
  NAND2_X1  g158(.A1(KEYINPUT80), .A2(G104), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(G107), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n338), .A3(G104), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n342), .A2(new_n343), .A3(new_n346), .A4(new_n348), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n338), .A2(G104), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n343), .B1(new_n341), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AND4_X1   g166(.A1(new_n332), .A2(new_n337), .A3(new_n349), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n344), .A2(new_n345), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n347), .B1(new_n354), .B2(new_n338), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n346), .A2(new_n348), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n351), .B1(new_n357), .B2(new_n343), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n332), .B1(new_n358), .B2(new_n337), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n331), .B1(new_n353), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n230), .A2(new_n237), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n349), .A2(new_n362), .A3(new_n352), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n362), .B1(new_n349), .B2(new_n352), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(new_n365), .A3(KEYINPUT10), .ZN(new_n366));
  INV_X1    g180(.A(new_n251), .ZN(new_n367));
  OAI21_X1  g181(.A(G101), .B1(new_n355), .B2(new_n356), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(KEYINPUT4), .A3(new_n349), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n370), .B(G101), .C1(new_n355), .C2(new_n356), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n258), .A3(new_n371), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n360), .A2(new_n366), .A3(new_n367), .A4(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT83), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n372), .ZN(new_n376));
  OAI21_X1  g190(.A(G128), .B1(new_n233), .B2(new_n225), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n229), .B1(new_n333), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n349), .A2(new_n352), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT81), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n358), .A2(new_n332), .A3(new_n337), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n376), .B1(new_n382), .B2(new_n331), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n383), .A2(KEYINPUT83), .A3(new_n367), .A4(new_n366), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n375), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT12), .ZN(new_n386));
  INV_X1    g200(.A(new_n271), .ZN(new_n387));
  AOI22_X1  g201(.A1(new_n380), .A2(new_n381), .B1(new_n387), .B2(new_n379), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n386), .B1(new_n388), .B2(new_n367), .ZN(new_n389));
  OAI22_X1  g203(.A1(new_n353), .A2(new_n359), .B1(new_n271), .B2(new_n358), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT12), .A3(new_n251), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G140), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n262), .A2(G227), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n394), .B(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(new_n375), .B2(new_n384), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n383), .A2(new_n366), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n251), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n393), .A2(new_n396), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G469), .B1(new_n400), .B2(G902), .ZN(new_n401));
  INV_X1    g215(.A(G469), .ZN(new_n402));
  AOI221_X4 g216(.A(new_n396), .B1(new_n391), .B2(new_n389), .C1(new_n375), .C2(new_n384), .ZN(new_n403));
  INV_X1    g217(.A(new_n396), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n385), .B2(new_n399), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n402), .B(new_n314), .C1(new_n403), .C2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n330), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(G210), .B1(G237), .B2(G902), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT87), .ZN(new_n409));
  INV_X1    g223(.A(G125), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n387), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n257), .A2(G125), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G224), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(G953), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n413), .B(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n369), .A2(new_n269), .A3(new_n371), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G110), .B(G122), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(KEYINPUT85), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n379), .A2(KEYINPUT82), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n349), .A2(new_n362), .A3(new_n352), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n240), .A2(KEYINPUT5), .ZN(new_n425));
  INV_X1    g239(.A(G116), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n426), .A2(KEYINPUT5), .A3(G119), .ZN(new_n427));
  INV_X1    g241(.A(G113), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n241), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n423), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT84), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT84), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n423), .A2(new_n433), .A3(new_n424), .A4(new_n430), .ZN(new_n434));
  AOI211_X1 g248(.A(new_n419), .B(new_n422), .C1(new_n432), .C2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n419), .B1(new_n432), .B2(new_n434), .ZN(new_n437));
  XOR2_X1   g251(.A(new_n421), .B(KEYINPUT86), .Z(new_n438));
  OAI22_X1  g252(.A1(new_n435), .A2(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n438), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n432), .A2(new_n434), .ZN(new_n441));
  OAI211_X1 g255(.A(KEYINPUT6), .B(new_n440), .C1(new_n441), .C2(new_n419), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n417), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT7), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n413), .B1(new_n444), .B2(new_n415), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n411), .A2(KEYINPUT7), .A3(new_n416), .A4(new_n412), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n379), .A2(new_n430), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n379), .A2(new_n430), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n421), .B(KEYINPUT8), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n445), .A2(new_n446), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n314), .B1(new_n435), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n409), .B1(new_n443), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n436), .B1(new_n437), .B2(new_n421), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n437), .A2(new_n438), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n442), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n417), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n409), .ZN(new_n459));
  INV_X1    g273(.A(new_n452), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G214), .B1(G237), .B2(G902), .ZN(new_n463));
  INV_X1    g277(.A(G478), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(KEYINPUT15), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(G217), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n328), .A2(new_n467), .A3(G953), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n213), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT68), .A2(G128), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(G143), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n227), .A2(G128), .A3(new_n216), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n247), .ZN(new_n474));
  INV_X1    g288(.A(G122), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(G116), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n426), .A2(G122), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n338), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n477), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n479), .A2(G107), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n474), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n217), .A2(new_n218), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(KEYINPUT13), .A3(G128), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT13), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n473), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n485), .A3(new_n472), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n481), .B1(new_n486), .B2(G134), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n476), .A2(KEYINPUT14), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n479), .A2(new_n488), .A3(G107), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n476), .B(new_n477), .C1(KEYINPUT14), .C2(new_n338), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n472), .A2(new_n473), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n191), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n491), .B1(new_n493), .B2(new_n474), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n469), .B1(new_n487), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n474), .ZN(new_n496));
  INV_X1    g310(.A(new_n491), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n486), .A2(G134), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n498), .B(new_n468), .C1(new_n499), .C2(new_n481), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT95), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n495), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(KEYINPUT95), .B(new_n469), .C1(new_n487), .C2(new_n494), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n314), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT96), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n502), .A2(KEYINPUT96), .A3(new_n314), .A4(new_n503), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n466), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n465), .B1(new_n504), .B2(new_n505), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G475), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n227), .A2(KEYINPUT88), .A3(new_n216), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n261), .A2(new_n262), .A3(G214), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G214), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n515), .A2(G237), .A3(G953), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n516), .B(new_n220), .C1(new_n226), .C2(KEYINPUT88), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(KEYINPUT18), .A2(G131), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n514), .A2(new_n517), .A3(KEYINPUT18), .A4(G131), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n522));
  XNOR2_X1  g336(.A(G125), .B(G140), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n522), .B1(new_n523), .B2(new_n207), .ZN(new_n524));
  INV_X1    g338(.A(G140), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G125), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n410), .A2(G140), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(KEYINPUT89), .A3(G146), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n221), .A2(new_n222), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n523), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n524), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n520), .A2(new_n521), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT90), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n520), .A2(new_n521), .A3(new_n535), .A4(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n513), .A2(G143), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT88), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n227), .A2(new_n539), .A3(new_n216), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n538), .A2(new_n540), .B1(new_n512), .B2(new_n513), .ZN(new_n541));
  INV_X1    g355(.A(new_n204), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT91), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n518), .A2(new_n544), .A3(new_n204), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n541), .A2(new_n542), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n543), .A2(new_n545), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT16), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n525), .A3(G125), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n528), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n207), .ZN(new_n552));
  OAI211_X1 g366(.A(G146), .B(new_n550), .C1(new_n528), .C2(new_n549), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n518), .A2(new_n204), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(KEYINPUT17), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(G113), .B(G122), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT93), .B(G104), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT94), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n537), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n534), .A2(new_n536), .B1(new_n548), .B2(new_n556), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n562), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n511), .B1(new_n564), .B2(new_n314), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n523), .A2(KEYINPUT19), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n523), .A2(KEYINPUT19), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT92), .B(new_n530), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n553), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n523), .B(KEYINPUT19), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT92), .B1(new_n570), .B2(new_n530), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n537), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n562), .B1(new_n575), .B2(new_n560), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT20), .ZN(new_n577));
  NOR2_X1   g391(.A1(G475), .A2(G902), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n537), .A2(new_n557), .A3(new_n561), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n560), .B1(new_n537), .B2(new_n574), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n578), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT20), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n565), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(G234), .A2(G237), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(G952), .A3(new_n262), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT21), .B(G898), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(G902), .A3(G953), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n586), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n590), .B(KEYINPUT97), .Z(new_n591));
  AND3_X1   g405(.A1(new_n510), .A2(new_n584), .A3(new_n591), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n462), .A2(new_n463), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT78), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT25), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT22), .B(G137), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n596), .B(new_n597), .Z(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT23), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(KEYINPUT74), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT74), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(KEYINPUT23), .ZN(new_n603));
  INV_X1    g417(.A(G119), .ZN(new_n604));
  OAI22_X1  g418(.A1(new_n601), .A2(new_n603), .B1(new_n604), .B2(G128), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n470), .A2(KEYINPUT23), .A3(G119), .A4(new_n471), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(G128), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n212), .A2(new_n213), .A3(new_n604), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT73), .B1(new_n335), .B2(G119), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT73), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(new_n604), .A3(G128), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT24), .B(G110), .Z(new_n615));
  AOI22_X1  g429(.A1(new_n608), .A2(G110), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT75), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n616), .A2(new_n617), .A3(new_n554), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n616), .B2(new_n554), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n553), .A2(new_n531), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n608), .A2(G110), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n614), .A2(new_n615), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(KEYINPUT76), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n608), .A2(G110), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n614), .A2(new_n615), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n554), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT75), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n616), .A2(new_n617), .A3(new_n554), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n624), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT76), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n599), .B1(new_n625), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n598), .B1(new_n631), .B2(new_n632), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n634), .A2(G902), .A3(new_n635), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n594), .B(new_n595), .C1(new_n636), .C2(KEYINPUT77), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n467), .B1(G234), .B2(new_n314), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT25), .B1(new_n636), .B2(new_n594), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n631), .A2(new_n632), .ZN(new_n640));
  AOI211_X1 g454(.A(KEYINPUT76), .B(new_n624), .C1(new_n630), .C2(new_n629), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n598), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n635), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n314), .A3(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT77), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT78), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n637), .B(new_n638), .C1(new_n639), .C2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n634), .A2(new_n635), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT79), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n638), .A2(G902), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n326), .A2(new_n407), .A3(new_n593), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G101), .ZN(G3));
  AOI21_X1  g469(.A(G902), .B1(new_n297), .B2(new_n299), .ZN(new_n656));
  INV_X1    g470(.A(G472), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n295), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n653), .A2(new_n407), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT33), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n502), .A2(new_n661), .A3(new_n503), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n495), .A2(new_n500), .A3(KEYINPUT33), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n662), .A2(G478), .A3(new_n314), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n504), .A2(new_n464), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n584), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n463), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n458), .A2(new_n460), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(new_n408), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n443), .A2(new_n408), .A3(new_n452), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n672), .A2(new_n591), .A3(new_n674), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n660), .A2(new_n669), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT34), .B(G104), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  NAND3_X1  g492(.A1(new_n579), .A2(new_n583), .A3(KEYINPUT98), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT98), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n565), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(new_n508), .B2(new_n509), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n660), .A2(new_n675), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT35), .B(G107), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G9));
  INV_X1    g504(.A(new_n638), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n691), .B1(new_n646), .B2(new_n595), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n594), .B1(new_n636), .B2(KEYINPUT77), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n595), .B1(new_n644), .B2(KEYINPUT78), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n631), .B(KEYINPUT99), .Z(new_n696));
  NOR2_X1   g510(.A1(new_n599), .A2(KEYINPUT36), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n696), .B(new_n697), .Z(new_n698));
  AOI22_X1  g512(.A1(new_n692), .A2(new_n695), .B1(new_n650), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n658), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n407), .A3(new_n593), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT37), .B(G110), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G12));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n506), .A2(new_n507), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n465), .ZN(new_n706));
  INV_X1    g520(.A(new_n509), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n565), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n589), .A2(G900), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n586), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n708), .A2(new_n682), .A3(new_n679), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT100), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT100), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n686), .A2(new_n713), .A3(new_n710), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n672), .A2(new_n674), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n704), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n699), .B1(new_n303), .B2(new_n325), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n452), .B1(new_n456), .B2(new_n457), .ZN(new_n719));
  INV_X1    g533(.A(new_n408), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n463), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n673), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n712), .A2(new_n722), .A3(new_n714), .A4(KEYINPUT101), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n717), .A2(new_n407), .A3(new_n718), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G128), .ZN(G30));
  XNOR2_X1  g539(.A(new_n710), .B(KEYINPUT39), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n407), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT40), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n321), .A2(new_n266), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n314), .B1(new_n309), .B2(new_n266), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n303), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n462), .B(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n699), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n706), .A2(new_n707), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n582), .A2(KEYINPUT20), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n684), .B1(new_n680), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n736), .A2(new_n670), .A3(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n728), .A2(new_n733), .A3(new_n735), .A4(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(new_n482), .Z(G45));
  NAND2_X1  g557(.A1(new_n668), .A2(new_n710), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n718), .A2(new_n407), .A3(new_n722), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT103), .B(G146), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G48));
  AOI21_X1  g562(.A(new_n652), .B1(new_n303), .B2(new_n325), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n675), .A2(new_n669), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n314), .B1(new_n403), .B2(new_n405), .ZN(new_n751));
  NAND2_X1  g565(.A1(KEYINPUT104), .A2(G469), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n330), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n314), .B(new_n752), .C1(new_n403), .C2(new_n405), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n750), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(KEYINPUT41), .B(G113), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(G15));
  NOR2_X1   g574(.A1(new_n675), .A2(new_n687), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n749), .A2(new_n761), .A3(new_n757), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G116), .ZN(G18));
  NAND3_X1  g577(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n716), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n718), .A2(new_n765), .A3(new_n592), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G119), .ZN(G21));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n656), .A2(new_n657), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n287), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n286), .B1(new_n308), .B2(new_n260), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n771), .B1(new_n772), .B2(new_n310), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n266), .B1(new_n773), .B2(new_n306), .ZN(new_n774));
  OAI21_X1  g588(.A(KEYINPUT105), .B1(new_n774), .B2(new_n294), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n287), .B1(new_n305), .B2(KEYINPUT71), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n310), .B1(new_n309), .B2(KEYINPUT28), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n289), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT105), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n299), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n775), .A2(new_n780), .A3(new_n282), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT106), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n781), .A2(new_n782), .A3(new_n187), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n782), .B1(new_n781), .B2(new_n187), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n653), .B(new_n770), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n721), .A2(new_n673), .A3(new_n740), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n757), .A2(new_n591), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n768), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n781), .A2(new_n187), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT106), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n781), .A2(new_n782), .A3(new_n187), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n769), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n754), .A2(new_n755), .A3(new_n591), .A4(new_n756), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n672), .A2(new_n674), .A3(new_n739), .A4(new_n737), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n792), .A2(KEYINPUT107), .A3(new_n653), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n788), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G122), .ZN(G24));
  OAI211_X1 g612(.A(new_n770), .B(new_n736), .C1(new_n783), .C2(new_n784), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n757), .A2(new_n722), .A3(new_n745), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT108), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT108), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n764), .A2(new_n716), .A3(new_n744), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n792), .A2(new_n802), .A3(new_n803), .A4(new_n736), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(KEYINPUT109), .B(G125), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(G27));
  AND3_X1   g621(.A1(new_n453), .A2(new_n461), .A3(new_n463), .ZN(new_n808));
  NAND2_X1  g622(.A1(G469), .A2(G902), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n393), .A2(new_n396), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n397), .A2(new_n399), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(G469), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n406), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n808), .A2(new_n813), .A3(new_n755), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n749), .A2(new_n814), .A3(new_n745), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT42), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n749), .A2(new_n814), .A3(KEYINPUT42), .A4(new_n745), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G131), .ZN(G33));
  INV_X1    g634(.A(KEYINPUT110), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n715), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n712), .A2(new_n714), .A3(KEYINPUT110), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n749), .A2(new_n814), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(new_n194), .ZN(G36));
  OR2_X1    g641(.A1(new_n400), .A2(KEYINPUT45), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n400), .A2(KEYINPUT45), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(G469), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n809), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT46), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n406), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n833), .A2(KEYINPUT111), .B1(new_n832), .B2(new_n831), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(KEYINPUT111), .B2(new_n833), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n835), .A2(new_n755), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT43), .B1(new_n584), .B2(KEYINPUT112), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n584), .A2(new_n666), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n736), .A2(new_n839), .A3(new_n658), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT44), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n808), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n840), .B2(new_n841), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n836), .A2(new_n726), .A3(new_n842), .A4(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(G137), .ZN(G39));
  NOR4_X1   g660(.A1(new_n326), .A2(new_n653), .A3(new_n843), .A4(new_n744), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT113), .Z(new_n848));
  AND3_X1   g662(.A1(new_n835), .A2(KEYINPUT47), .A3(new_n755), .ZN(new_n849));
  AOI21_X1  g663(.A(KEYINPUT47), .B1(new_n835), .B2(new_n755), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(KEYINPUT114), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(G140), .ZN(G42));
  NAND2_X1  g670(.A1(new_n754), .A2(new_n756), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT49), .ZN(new_n858));
  OR4_X1    g672(.A1(new_n652), .A2(new_n330), .A3(new_n670), .A4(new_n838), .ZN(new_n859));
  OR4_X1    g673(.A1(new_n733), .A2(new_n858), .A3(new_n859), .A4(new_n735), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n757), .A2(new_n670), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n735), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  INV_X1    g678(.A(new_n586), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n839), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n792), .A2(new_n653), .A3(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT50), .Z(new_n869));
  NOR2_X1   g683(.A1(new_n857), .A2(new_n755), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n849), .A2(new_n850), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n867), .A2(new_n843), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n733), .A2(new_n652), .A3(new_n586), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n843), .A2(new_n764), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n584), .A3(new_n667), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n866), .A2(new_n876), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(new_n799), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT51), .B1(new_n881), .B2(KEYINPUT117), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n882), .B1(KEYINPUT117), .B2(new_n881), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n874), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n877), .A2(new_n668), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(G952), .A3(new_n262), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n866), .A2(new_n749), .A3(new_n876), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT48), .Z(new_n888));
  INV_X1    g702(.A(new_n867), .ZN(new_n889));
  AOI211_X1 g703(.A(new_n886), .B(new_n888), .C1(new_n765), .C2(new_n889), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n890), .A2(KEYINPUT118), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(KEYINPUT118), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n884), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n801), .A2(new_n804), .ZN(new_n895));
  INV_X1    g709(.A(new_n710), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n736), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n407), .A3(new_n733), .A4(new_n786), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n724), .A2(new_n746), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT52), .B1(new_n895), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n724), .A2(new_n746), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT52), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n805), .A3(new_n902), .A4(new_n898), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n758), .A2(new_n766), .A3(new_n762), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n788), .B2(new_n796), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n719), .A2(new_n459), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n443), .A2(new_n409), .A3(new_n452), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n463), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n739), .A2(new_n510), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n591), .B1(new_n910), .B2(new_n668), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(new_n407), .A3(new_n653), .A4(new_n659), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n654), .A2(new_n913), .A3(new_n701), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT115), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n670), .B1(new_n453), .B2(new_n461), .ZN(new_n916));
  AND4_X1   g730(.A1(new_n755), .A2(new_n813), .A3(new_n916), .A4(new_n592), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n749), .B2(new_n700), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT115), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n918), .A2(new_n919), .A3(new_n913), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n915), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n826), .B1(new_n817), .B2(new_n818), .ZN(new_n922));
  NOR4_X1   g736(.A1(new_n683), .A2(new_n737), .A3(new_n565), .A4(new_n896), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n718), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n799), .B2(new_n744), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n814), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n906), .A2(new_n921), .A3(new_n922), .A4(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n894), .B1(new_n904), .B2(new_n927), .ZN(new_n928));
  AND3_X1   g742(.A1(new_n758), .A2(new_n766), .A3(new_n762), .ZN(new_n929));
  AND4_X1   g743(.A1(new_n919), .A2(new_n654), .A3(new_n701), .A4(new_n913), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n919), .B1(new_n918), .B2(new_n913), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n797), .B(new_n929), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n826), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n926), .A2(new_n819), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n900), .A3(new_n903), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n898), .A2(new_n746), .ZN(new_n937));
  AOI21_X1  g751(.A(KEYINPUT53), .B1(new_n937), .B2(KEYINPUT52), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n928), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT54), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n894), .B1(new_n937), .B2(KEYINPUT52), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n935), .A2(new_n900), .A3(new_n903), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n928), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n940), .B1(KEYINPUT54), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n881), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT51), .B1(new_n874), .B2(new_n945), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n893), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(G952), .A2(G953), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n860), .B1(new_n947), .B2(new_n948), .ZN(G75));
  AOI21_X1  g763(.A(new_n314), .B1(new_n928), .B2(new_n942), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT56), .B1(new_n950), .B2(G210), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n456), .B(new_n457), .ZN(new_n952));
  XNOR2_X1  g766(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n262), .A2(G952), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n951), .A2(new_n954), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n959), .A2(KEYINPUT120), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(KEYINPUT120), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G51));
  AND2_X1   g776(.A1(new_n943), .A2(KEYINPUT54), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n943), .A2(KEYINPUT54), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n809), .B(KEYINPUT57), .ZN(new_n966));
  OAI22_X1  g780(.A1(new_n965), .A2(new_n966), .B1(new_n405), .B2(new_n403), .ZN(new_n967));
  INV_X1    g781(.A(new_n830), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n950), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT121), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n956), .B1(new_n967), .B2(new_n970), .ZN(G54));
  NAND3_X1  g785(.A1(new_n950), .A2(KEYINPUT58), .A3(G475), .ZN(new_n972));
  INV_X1    g786(.A(new_n576), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n974), .A2(new_n975), .A3(new_n956), .ZN(G60));
  XOR2_X1   g790(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n977));
  NOR2_X1   g791(.A1(new_n464), .A2(new_n314), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AOI22_X1  g794(.A1(new_n944), .A2(new_n980), .B1(new_n662), .B2(new_n663), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n662), .A2(new_n663), .A3(new_n980), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n957), .B1(new_n965), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n981), .A2(new_n983), .ZN(G63));
  NAND2_X1  g798(.A1(G217), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT123), .Z(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT60), .Z(new_n987));
  NAND2_X1  g801(.A1(new_n943), .A2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n649), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n987), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(new_n928), .B2(new_n942), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n698), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n990), .A2(KEYINPUT61), .A3(new_n957), .A4(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT125), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT61), .ZN(new_n996));
  AOI21_X1  g810(.A(KEYINPUT124), .B1(new_n990), .B2(new_n957), .ZN(new_n997));
  OAI211_X1 g811(.A(KEYINPUT124), .B(new_n957), .C1(new_n992), .C2(new_n649), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n993), .ZN(new_n999));
  OAI211_X1 g813(.A(new_n995), .B(new_n996), .C1(new_n997), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT124), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n649), .B1(new_n943), .B2(new_n987), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1002), .B1(new_n1003), .B2(new_n956), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1004), .A2(new_n998), .A3(new_n993), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n995), .B1(new_n1005), .B2(new_n996), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n994), .B1(new_n1001), .B2(new_n1006), .ZN(G66));
  OAI21_X1  g821(.A(G953), .B1(new_n587), .B2(new_n414), .ZN(new_n1008));
  INV_X1    g822(.A(new_n932), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1008), .B1(new_n1009), .B2(G953), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n439), .B(new_n442), .C1(G898), .C2(new_n262), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(G69));
  AOI21_X1  g826(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n262), .A2(G900), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT127), .Z(new_n1015));
  NAND4_X1  g829(.A1(new_n836), .A2(new_n749), .A3(new_n726), .A4(new_n786), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n901), .A2(new_n805), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n845), .A2(new_n1016), .A3(new_n922), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1018), .B1(new_n853), .B2(new_n854), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1015), .B1(new_n1019), .B2(G953), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n268), .A2(new_n275), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(new_n570), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  AND2_X1   g837(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1017), .A2(new_n742), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n1025), .A2(KEYINPUT62), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(KEYINPUT62), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n910), .A2(new_n668), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1028), .B(KEYINPUT126), .ZN(new_n1029));
  NAND4_X1  g843(.A1(new_n727), .A2(new_n1029), .A3(new_n749), .A4(new_n808), .ZN(new_n1030));
  AND4_X1   g844(.A1(new_n845), .A2(new_n1026), .A3(new_n1027), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(G953), .B1(new_n1031), .B2(new_n855), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n1032), .A2(new_n1023), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1013), .B1(new_n1024), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1013), .ZN(new_n1036));
  OAI211_X1 g850(.A(new_n1035), .B(new_n1036), .C1(new_n1032), .C2(new_n1023), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1034), .A2(new_n1037), .ZN(G72));
  NAND3_X1  g852(.A1(new_n292), .A2(new_n260), .A3(new_n289), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n1019), .A2(new_n1009), .ZN(new_n1040));
  NAND2_X1  g854(.A1(G472), .A2(G902), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT63), .Z(new_n1042));
  AOI21_X1  g856(.A(new_n1039), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1031), .A2(new_n855), .A3(new_n1009), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n729), .B1(new_n1044), .B2(new_n1042), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n322), .A2(new_n298), .ZN(new_n1046));
  AND3_X1   g860(.A1(new_n939), .A2(new_n1042), .A3(new_n1046), .ZN(new_n1047));
  NOR4_X1   g861(.A1(new_n1043), .A2(new_n1045), .A3(new_n956), .A4(new_n1047), .ZN(G57));
endmodule


