//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n749,
    new_n750, new_n751, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT93), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(new_n205), .B2(new_n204), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n208), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT14), .B(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n204), .A2(KEYINPUT15), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n207), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n214), .B1(new_n207), .B2(new_n212), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT94), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G1gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(G1gat), .B2(new_n218), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n215), .B(KEYINPUT94), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(KEYINPUT17), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n215), .A2(KEYINPUT17), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n223), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n202), .B(new_n225), .C1(new_n227), .C2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT18), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(new_n223), .A3(new_n228), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n235), .A2(KEYINPUT18), .A3(new_n202), .A4(new_n225), .ZN(new_n236));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(G197gat), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT11), .B(G169gat), .Z(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n240), .B(KEYINPUT12), .Z(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n223), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n202), .B(KEYINPUT13), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n232), .A2(new_n236), .A3(new_n242), .A4(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n230), .A2(new_n231), .B1(new_n244), .B2(new_n245), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n242), .B1(new_n249), .B2(new_n236), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(G57gat), .A2(G64gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(G57gat), .A2(G64gat), .ZN(new_n253));
  AND2_X1   g052(.A1(G71gat), .A2(G78gat), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n252), .B(new_n253), .C1(new_n254), .C2(KEYINPUT9), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(KEYINPUT95), .B2(new_n254), .ZN(new_n256));
  XNOR2_X1  g055(.A(G71gat), .B(G78gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT21), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G231gat), .A2(G233gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(G127gat), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n223), .B1(new_n258), .B2(new_n259), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT96), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(G155gat), .ZN(new_n268));
  XOR2_X1   g067(.A(G183gat), .B(G211gat), .Z(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n265), .B(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(G232gat), .A2(G233gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(KEYINPUT41), .ZN(new_n273));
  XNOR2_X1  g072(.A(G134gat), .B(G162gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n277));
  NAND2_X1  g076(.A1(G85gat), .A2(G92gat), .ZN(new_n278));
  OR2_X1    g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n278), .ZN(new_n280));
  NAND2_X1  g079(.A1(G99gat), .A2(G106gat), .ZN(new_n281));
  INV_X1    g080(.A(G85gat), .ZN(new_n282));
  INV_X1    g081(.A(G92gat), .ZN(new_n283));
  AOI22_X1  g082(.A1(KEYINPUT8), .A2(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n279), .A2(new_n280), .A3(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(G99gat), .B(G106gat), .Z(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n286), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n234), .A2(new_n228), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n289), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n217), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n272), .A2(KEYINPUT41), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(G190gat), .B(G218gat), .Z(new_n295));
  NOR3_X1   g094(.A1(new_n290), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n295), .ZN(new_n297));
  INV_X1    g096(.A(new_n294), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n234), .A2(new_n228), .A3(new_n289), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n276), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n295), .B1(new_n290), .B2(new_n294), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n298), .A2(new_n297), .A3(new_n299), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n275), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n289), .A2(new_n258), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT10), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n289), .A2(new_n258), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  OR3_X1    g108(.A1(new_n289), .A2(new_n307), .A3(new_n258), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G230gat), .ZN(new_n312));
  INV_X1    g111(.A(G233gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n306), .A2(new_n308), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(new_n314), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G120gat), .B(G148gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(G176gat), .B(G204gat), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n316), .A2(new_n318), .A3(new_n322), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n271), .A2(new_n305), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT85), .ZN(new_n329));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT31), .B(G50gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT81), .ZN(new_n333));
  INV_X1    g132(.A(G228gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n334), .A2(new_n313), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n337));
  AND2_X1   g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(KEYINPUT78), .A3(KEYINPUT2), .ZN(new_n342));
  AND2_X1   g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  OR2_X1    g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(KEYINPUT77), .A3(new_n341), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT77), .ZN(new_n349));
  NOR2_X1   g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n338), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n347), .A2(new_n341), .ZN(new_n354));
  INV_X1    g153(.A(G162gat), .ZN(new_n355));
  OR2_X1    g154(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(KEYINPUT79), .A2(G155gat), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n354), .B(new_n345), .C1(new_n358), .C2(new_n339), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n362));
  XNOR2_X1  g161(.A(G211gat), .B(G218gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(G197gat), .B(G204gat), .ZN(new_n364));
  INV_X1    g163(.A(G211gat), .ZN(new_n365));
  INV_X1    g164(.A(G218gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT73), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT73), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G218gat), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n365), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n363), .B(new_n364), .C1(new_n370), .C2(KEYINPUT22), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT22), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT73), .B(G218gat), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n373), .B1(new_n374), .B2(new_n365), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n363), .B1(new_n375), .B2(new_n364), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n362), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n361), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n363), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n367), .A2(new_n369), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT22), .B1(new_n381), .B2(G211gat), .ZN(new_n382));
  INV_X1    g181(.A(new_n364), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n380), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT74), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n371), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n376), .A2(KEYINPUT74), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n353), .A2(new_n378), .A3(new_n359), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n386), .A2(new_n387), .B1(new_n388), .B2(new_n362), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n336), .B1(new_n379), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n387), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n362), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n335), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n395));
  XNOR2_X1  g194(.A(G141gat), .B(G148gat), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT78), .B1(new_n341), .B2(KEYINPUT2), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g197(.A1(new_n398), .A2(new_n342), .B1(new_n351), .B2(new_n348), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT79), .B(G155gat), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n339), .B1(new_n400), .B2(G162gat), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n354), .A2(new_n345), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n395), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n353), .A2(KEYINPUT80), .A3(new_n359), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n386), .A2(new_n362), .A3(new_n387), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n407), .B2(new_n378), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n390), .B1(new_n394), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(KEYINPUT82), .B(G22gat), .Z(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n409), .A2(KEYINPUT84), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT84), .B1(new_n409), .B2(new_n411), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n390), .B(new_n410), .C1(new_n408), .C2(new_n394), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT83), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n407), .A2(new_n378), .ZN(new_n417));
  INV_X1    g216(.A(new_n406), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n389), .A2(new_n336), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT83), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n421), .A2(new_n422), .A3(new_n390), .A4(new_n410), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n333), .B1(new_n414), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n415), .A2(new_n332), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(G22gat), .B2(new_n409), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n329), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT29), .B1(new_n384), .B2(new_n371), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n360), .B1(new_n430), .B2(KEYINPUT3), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n393), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g231(.A1(new_n419), .A2(new_n420), .B1(new_n432), .B2(new_n336), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n429), .B1(new_n433), .B2(new_n410), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n409), .A2(KEYINPUT84), .A3(new_n411), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n416), .A4(new_n423), .ZN(new_n436));
  INV_X1    g235(.A(new_n333), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n427), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT85), .ZN(new_n439));
  XNOR2_X1  g238(.A(G1gat), .B(G29gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(KEYINPUT0), .ZN(new_n441));
  XNOR2_X1  g240(.A(G57gat), .B(G85gat), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n441), .B(new_n442), .Z(new_n443));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT71), .ZN(new_n445));
  INV_X1    g244(.A(G127gat), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n445), .B1(new_n446), .B2(G134gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT1), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(G113gat), .B2(G120gat), .ZN(new_n449));
  AND2_X1   g248(.A1(G113gat), .A2(G120gat), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G127gat), .B(G134gat), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n452), .B(new_n447), .C1(new_n450), .C2(new_n449), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n456), .A2(new_n353), .A3(new_n359), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT4), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT4), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n456), .A2(new_n353), .A3(new_n459), .A4(new_n359), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n353), .A2(KEYINPUT80), .A3(new_n359), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT80), .B1(new_n353), .B2(new_n359), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n462), .A2(new_n463), .A3(new_n378), .ZN(new_n464));
  INV_X1    g263(.A(new_n456), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n388), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n444), .B(new_n461), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n444), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n462), .A2(new_n463), .A3(new_n456), .ZN(new_n469));
  INV_X1    g268(.A(new_n457), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(KEYINPUT5), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n404), .A2(KEYINPUT3), .A3(new_n405), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n388), .A2(new_n465), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n473), .A2(new_n474), .B1(new_n458), .B2(new_n460), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT5), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(new_n444), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n443), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT6), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n472), .A2(new_n443), .A3(new_n477), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n479), .B1(new_n482), .B2(new_n478), .ZN(new_n483));
  NAND2_X1  g282(.A1(G183gat), .A2(G190gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT24), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT24), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(G183gat), .A3(G190gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n489));
  OR3_X1    g288(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G169gat), .ZN(new_n492));
  INV_X1    g291(.A(G176gat), .ZN(new_n493));
  AND4_X1   g292(.A1(KEYINPUT66), .A2(new_n492), .A3(new_n493), .A4(KEYINPUT23), .ZN(new_n494));
  NOR2_X1   g293(.A1(G169gat), .A2(G176gat), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT66), .B1(new_n495), .B2(KEYINPUT23), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n492), .A2(new_n493), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT67), .ZN(new_n499));
  OAI22_X1  g298(.A1(new_n492), .A2(new_n493), .B1(new_n499), .B2(KEYINPUT23), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(KEYINPUT23), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n491), .A2(new_n497), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT25), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n488), .B1(G183gat), .B2(G190gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT23), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n507), .A2(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n495), .B1(new_n508), .B2(new_n501), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT25), .B1(new_n498), .B2(new_n507), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n504), .A2(new_n505), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n513), .A2(KEYINPUT69), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n513), .A2(KEYINPUT69), .B1(G169gat), .B2(G176gat), .ZN(new_n515));
  NOR3_X1   g314(.A1(new_n498), .A2(KEYINPUT70), .A3(KEYINPUT26), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT70), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT26), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n495), .B2(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n514), .B(new_n515), .C1(new_n516), .C2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G183gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(KEYINPUT27), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT27), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G183gat), .ZN(new_n524));
  INV_X1    g323(.A(G190gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n527));
  OR2_X1    g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n526), .A2(new_n527), .B1(G183gat), .B2(G190gat), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n520), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G226gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(new_n313), .ZN(new_n532));
  OAI22_X1  g331(.A1(new_n512), .A2(new_n530), .B1(KEYINPUT29), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n512), .A2(new_n530), .A3(new_n532), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n391), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n504), .A2(new_n505), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n511), .A2(new_n506), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n528), .A3(new_n529), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n539), .B(new_n540), .C1(new_n531), .C2(new_n313), .ZN(new_n541));
  INV_X1    g340(.A(new_n391), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n542), .A3(new_n533), .ZN(new_n543));
  XNOR2_X1  g342(.A(G8gat), .B(G36gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(G64gat), .B(G92gat), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n544), .B(new_n545), .Z(new_n546));
  NAND3_X1  g345(.A1(new_n536), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT30), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT76), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(KEYINPUT76), .A3(new_n548), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n546), .ZN(new_n554));
  INV_X1    g353(.A(new_n543), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n542), .B1(new_n541), .B2(new_n533), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n536), .A2(new_n543), .A3(KEYINPUT30), .A4(new_n546), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT75), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n558), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT75), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n483), .A2(new_n553), .A3(new_n560), .A4(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n428), .A2(new_n439), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT72), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n539), .A2(new_n566), .A3(new_n540), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT72), .B1(new_n512), .B2(new_n530), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n465), .ZN(new_n569));
  OAI211_X1 g368(.A(KEYINPUT72), .B(new_n456), .C1(new_n512), .C2(new_n530), .ZN(new_n570));
  NAND2_X1  g369(.A1(G227gat), .A2(G233gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(KEYINPUT64), .Z(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT32), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT33), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G15gat), .B(G43gat), .Z(new_n577));
  XNOR2_X1  g376(.A(G71gat), .B(G99gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n574), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n573), .B(KEYINPUT32), .C1(new_n575), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n572), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT34), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(new_n569), .B2(new_n570), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n569), .A2(new_n570), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n571), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n587), .B1(new_n589), .B2(KEYINPUT34), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n580), .A2(new_n590), .A3(new_n582), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n592), .A2(KEYINPUT36), .A3(new_n593), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n461), .B1(new_n464), .B2(new_n466), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT39), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n468), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n601), .A2(new_n443), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT89), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n444), .B(new_n457), .C1(new_n406), .C2(new_n456), .ZN(new_n604));
  OAI211_X1 g403(.A(KEYINPUT39), .B(new_n604), .C1(new_n475), .C2(new_n444), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT40), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n601), .A3(new_n443), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT89), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT88), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n472), .A2(new_n477), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(new_n612), .B2(new_n443), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n478), .A2(KEYINPUT88), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT87), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n605), .A2(new_n601), .A3(KEYINPUT87), .A4(new_n443), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n608), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n610), .A2(new_n613), .A3(new_n614), .A4(new_n618), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n547), .A2(KEYINPUT76), .A3(new_n548), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT76), .B1(new_n547), .B2(new_n548), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n559), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT86), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n553), .A2(KEYINPUT86), .A3(new_n559), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n619), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n436), .A2(new_n437), .ZN(new_n627));
  INV_X1    g426(.A(new_n427), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND2_X1   g428(.A1(new_n480), .A2(new_n481), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n630), .A3(new_n614), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n479), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n536), .A2(new_n543), .A3(KEYINPUT90), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n633), .B(KEYINPUT37), .C1(KEYINPUT90), .C2(new_n543), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT91), .B(KEYINPUT38), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n546), .B1(new_n536), .B2(new_n543), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n554), .A2(KEYINPUT37), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n547), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT37), .B1(new_n555), .B2(new_n556), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n640), .B1(new_n636), .B2(new_n637), .ZN(new_n641));
  INV_X1    g440(.A(new_n635), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n629), .B1(new_n632), .B2(new_n644), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n565), .B(new_n598), .C1(new_n626), .C2(new_n645), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n564), .A2(new_n594), .A3(new_n438), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT35), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n580), .A2(new_n590), .A3(new_n582), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n590), .B1(new_n580), .B2(new_n582), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n629), .A2(new_n651), .A3(new_n624), .A4(new_n625), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n632), .A2(new_n648), .ZN(new_n653));
  OAI22_X1  g452(.A1(new_n647), .A2(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n646), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(KEYINPUT92), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT92), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n646), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  AOI211_X1 g457(.A(new_n251), .B(new_n328), .C1(new_n656), .C2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n483), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT98), .B(G1gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1324gat));
  NAND2_X1  g462(.A1(new_n624), .A2(new_n625), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G8gat), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n659), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n222), .B1(new_n659), .B2(new_n664), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT42), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(KEYINPUT42), .B2(new_n667), .ZN(G1325gat));
  INV_X1    g469(.A(G15gat), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n659), .A2(new_n671), .A3(new_n651), .ZN(new_n672));
  INV_X1    g471(.A(new_n598), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n659), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n672), .B1(new_n675), .B2(new_n671), .ZN(G1326gat));
  NAND2_X1  g475(.A1(new_n428), .A2(new_n439), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n659), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  AND2_X1   g480(.A1(new_n301), .A2(new_n304), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n271), .A2(new_n251), .A3(new_n326), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n646), .A2(new_n657), .A3(new_n654), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n657), .B1(new_n646), .B2(new_n654), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n682), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n686), .A2(G29gat), .A3(new_n483), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT45), .Z(new_n688));
  AOI211_X1 g487(.A(KEYINPUT44), .B(new_n305), .C1(new_n646), .C2(new_n654), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(KEYINPUT44), .ZN(new_n691));
  INV_X1    g490(.A(new_n683), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n691), .A2(new_n483), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n688), .B1(new_n208), .B2(new_n693), .ZN(G1328gat));
  INV_X1    g493(.A(new_n664), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n686), .A2(G36gat), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT46), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n691), .A2(new_n695), .A3(new_n692), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n211), .B2(new_n698), .ZN(G1329gat));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n700));
  INV_X1    g499(.A(G43gat), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n691), .A2(new_n692), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n701), .B1(new_n702), .B2(new_n673), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n686), .A2(G43gat), .A3(new_n594), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n700), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n691), .A2(new_n677), .A3(new_n692), .ZN(new_n708));
  INV_X1    g507(.A(G50gat), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT102), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n677), .A2(G50gat), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n686), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n305), .B1(new_n656), .B2(new_n658), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT101), .B1(new_n715), .B2(new_n683), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n711), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n715), .A2(KEYINPUT101), .A3(new_n683), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n686), .A2(new_n713), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n718), .A2(new_n719), .A3(KEYINPUT102), .A4(new_n712), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n710), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n715), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(new_n438), .B(new_n683), .C1(new_n724), .C2(new_n689), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G50gat), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n714), .A2(new_n716), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n707), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT103), .B1(new_n722), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n709), .B1(new_n702), .B2(new_n438), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT48), .B1(new_n731), .B2(new_n727), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n678), .B(new_n683), .C1(new_n724), .C2(new_n689), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G50gat), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n734), .A2(new_n707), .A3(new_n717), .A4(new_n720), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n732), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n730), .A2(new_n737), .ZN(G1331gat));
  INV_X1    g537(.A(new_n271), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n232), .A2(new_n236), .A3(new_n246), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n241), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n247), .ZN(new_n742));
  NOR4_X1   g541(.A1(new_n739), .A2(new_n742), .A3(new_n682), .A4(new_n327), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n655), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT104), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n660), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT105), .B(G57gat), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1332gat));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n664), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT49), .B(G64gat), .Z(new_n751));
  OAI21_X1  g550(.A(new_n750), .B1(new_n749), .B2(new_n751), .ZN(G1333gat));
  NAND2_X1  g551(.A1(new_n745), .A2(new_n673), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n594), .A2(G71gat), .ZN(new_n754));
  AOI22_X1  g553(.A1(new_n753), .A2(G71gat), .B1(new_n745), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g555(.A1(new_n745), .A2(new_n678), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT106), .B(G78gat), .Z(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1335gat));
  AOI21_X1  g558(.A(new_n305), .B1(new_n646), .B2(new_n654), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n271), .A2(new_n742), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n762), .A2(KEYINPUT51), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(KEYINPUT51), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n326), .A2(new_n660), .A3(new_n282), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT108), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n761), .A2(new_n326), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT107), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n691), .A2(new_n483), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n771), .B2(new_n282), .ZN(G1336gat));
  NOR3_X1   g571(.A1(new_n695), .A2(G92gat), .A3(new_n327), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n762), .A2(KEYINPUT110), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n763), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT110), .B1(new_n762), .B2(new_n775), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n691), .A2(new_n770), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n283), .B1(new_n780), .B2(new_n664), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT52), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n773), .B1(new_n763), .B2(new_n764), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n781), .A2(new_n785), .A3(KEYINPUT111), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n782), .B1(new_n788), .B2(new_n789), .ZN(G1337gat));
  INV_X1    g589(.A(G99gat), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n651), .A2(new_n791), .A3(new_n326), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT112), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n765), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n691), .A2(new_n598), .A3(new_n770), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n791), .ZN(G1338gat));
  NOR3_X1   g595(.A1(new_n327), .A2(new_n629), .A3(G106gat), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n777), .B2(new_n778), .ZN(new_n799));
  INV_X1    g598(.A(G106gat), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n800), .B1(new_n780), .B2(new_n678), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT53), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n780), .A2(new_n438), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G106gat), .ZN(new_n804));
  AOI21_X1  g603(.A(KEYINPUT53), .B1(new_n765), .B2(new_n797), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n804), .A2(new_n805), .A3(KEYINPUT113), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT113), .B1(new_n804), .B2(new_n805), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n802), .B1(new_n806), .B2(new_n807), .ZN(G1339gat));
  NAND3_X1  g607(.A1(new_n309), .A2(new_n310), .A3(new_n314), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n316), .A2(KEYINPUT54), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n314), .B1(new_n309), .B2(new_n310), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n322), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n810), .A2(KEYINPUT55), .A3(new_n813), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n816), .A2(new_n325), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n202), .B1(new_n235), .B2(new_n225), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n244), .A2(new_n245), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n240), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n247), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n682), .A3(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n816), .A2(new_n325), .A3(new_n817), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n305), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(KEYINPUT114), .A3(new_n822), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n326), .A2(new_n247), .A3(new_n821), .ZN(new_n831));
  AOI22_X1  g630(.A1(new_n818), .A2(new_n742), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n822), .A2(KEYINPUT115), .A3(new_n326), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n682), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n739), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n328), .A2(new_n742), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n483), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n652), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n742), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n678), .B1(new_n835), .B2(new_n837), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n695), .A2(new_n660), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(new_n594), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n742), .A2(G113gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(G1340gat));
  OR3_X1    g647(.A1(new_n840), .A2(G120gat), .A3(new_n327), .ZN(new_n849));
  INV_X1    g648(.A(new_n846), .ZN(new_n850));
  OAI21_X1  g649(.A(G120gat), .B1(new_n850), .B2(new_n327), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(KEYINPUT116), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n849), .B1(new_n852), .B2(new_n853), .ZN(G1341gat));
  OAI21_X1  g653(.A(G127gat), .B1(new_n850), .B2(new_n739), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n841), .A2(new_n446), .A3(new_n271), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1342gat));
  OR3_X1    g656(.A1(new_n840), .A2(G134gat), .A3(new_n305), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n859));
  OAI21_X1  g658(.A(G134gat), .B1(new_n850), .B2(new_n305), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(KEYINPUT56), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(G1343gat));
  NOR2_X1   g661(.A1(new_n673), .A2(new_n844), .ZN(new_n863));
  INV_X1    g662(.A(G141gat), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n251), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n677), .A2(new_n867), .ZN(new_n868));
  AND4_X1   g667(.A1(KEYINPUT114), .A2(new_n818), .A3(new_n682), .A4(new_n822), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT114), .B1(new_n827), .B2(new_n822), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n831), .B1(new_n251), .B2(new_n826), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n305), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n271), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n866), .B(new_n868), .C1(new_n874), .C2(new_n836), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n873), .A2(new_n825), .A3(new_n828), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n836), .B1(new_n876), .B2(new_n739), .ZN(new_n877));
  INV_X1    g676(.A(new_n868), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT117), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n835), .A2(new_n837), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n881), .B2(new_n438), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n863), .B(new_n865), .C1(new_n880), .C2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n673), .A2(new_n629), .A3(new_n664), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n838), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n864), .B1(new_n885), .B2(new_n251), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g686(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT119), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n883), .A2(KEYINPUT58), .A3(new_n886), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n887), .A2(new_n892), .A3(new_n888), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(G1344gat));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n863), .B1(new_n880), .B2(new_n882), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n895), .B(G148gat), .C1(new_n896), .C2(new_n327), .ZN(new_n897));
  INV_X1    g696(.A(G148gat), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n873), .A2(new_n823), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n836), .B1(new_n899), .B2(new_n739), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n677), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n900), .A2(new_n901), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n867), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n881), .A2(KEYINPUT57), .A3(new_n438), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n673), .A2(new_n844), .A3(new_n327), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n898), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n897), .B1(new_n909), .B2(new_n895), .ZN(new_n910));
  INV_X1    g709(.A(new_n885), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n898), .A3(new_n326), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1345gat));
  OAI21_X1  g712(.A(new_n400), .B1(new_n896), .B2(new_n739), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n271), .A2(new_n356), .A3(new_n357), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n885), .B2(new_n915), .ZN(G1346gat));
  NOR3_X1   g715(.A1(new_n896), .A2(new_n355), .A3(new_n305), .ZN(new_n917));
  AOI21_X1  g716(.A(G162gat), .B1(new_n911), .B2(new_n682), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n695), .A2(new_n660), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n835), .B2(new_n837), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n594), .A2(new_n438), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n742), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n843), .A2(new_n651), .A3(new_n920), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(new_n492), .A3(new_n251), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n926), .A2(new_n928), .ZN(G1348gat));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n493), .A3(new_n326), .ZN(new_n930));
  OAI21_X1  g729(.A(G176gat), .B1(new_n927), .B2(new_n327), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1349gat));
  AND4_X1   g731(.A1(new_n522), .A2(new_n925), .A3(new_n524), .A4(new_n271), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n934), .A2(KEYINPUT121), .ZN(new_n935));
  INV_X1    g734(.A(new_n927), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n521), .B1(new_n936), .B2(new_n271), .ZN(new_n937));
  OR3_X1    g736(.A1(new_n933), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n933), .B2(new_n937), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1350gat));
  NOR3_X1   g739(.A1(new_n924), .A2(G190gat), .A3(new_n305), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT122), .ZN(new_n942));
  OAI21_X1  g741(.A(G190gat), .B1(new_n927), .B2(new_n305), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n944), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(G1351gat));
  NAND4_X1  g746(.A1(new_n881), .A2(new_n438), .A3(new_n598), .A4(new_n920), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT123), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  XOR2_X1   g749(.A(KEYINPUT124), .B(G197gat), .Z(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(new_n742), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n921), .A2(new_n673), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n907), .A2(new_n742), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n952), .B1(new_n954), .B2(new_n951), .ZN(G1352gat));
  AND2_X1   g754(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n956));
  NOR2_X1   g755(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n948), .A2(G204gat), .A3(new_n327), .ZN(new_n959));
  MUX2_X1   g758(.A(new_n958), .B(new_n956), .S(new_n959), .Z(new_n960));
  INV_X1    g759(.A(new_n904), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT57), .B1(new_n961), .B2(new_n902), .ZN(new_n962));
  INV_X1    g761(.A(new_n906), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n326), .B(new_n953), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT126), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G204gat), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n964), .A2(KEYINPUT126), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n960), .B1(new_n966), .B2(new_n967), .ZN(G1353gat));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n365), .A3(new_n271), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n271), .B(new_n953), .C1(new_n962), .C2(new_n963), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n970), .B2(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  AND4_X1   g772(.A1(new_n381), .A2(new_n907), .A3(new_n682), .A4(new_n953), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n366), .B1(new_n949), .B2(new_n305), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT127), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n977), .B(new_n366), .C1(new_n949), .C2(new_n305), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n974), .B1(new_n976), .B2(new_n978), .ZN(G1355gat));
endmodule


