//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(new_n461), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n467), .A2(KEYINPUT66), .A3(G137), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT66), .B1(new_n467), .B2(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  INV_X1    g046(.A(new_n466), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT65), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n465), .A2(new_n475), .A3(new_n466), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n474), .A2(G125), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n471), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n470), .A2(new_n479), .ZN(G160));
  AOI21_X1  g055(.A(new_n471), .B1(new_n465), .B2(new_n466), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n467), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n472), .C2(new_n473), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G114), .C2(new_n471), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n474), .A2(new_n476), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n492), .B2(new_n495), .ZN(G164));
  AND3_X1   g071(.A1(KEYINPUT67), .A2(KEYINPUT6), .A3(G651), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT6), .B1(KEYINPUT67), .B2(G651), .ZN(new_n498));
  OAI211_X1 g073(.A(G50), .B(G543), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  AND2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT5), .A2(G543), .ZN(new_n501));
  OAI22_X1  g076(.A1(new_n497), .A2(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G88), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n499), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(G62), .B1(new_n500), .B2(new_n501), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT68), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(new_n512), .A3(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n506), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n504), .B1(new_n515), .B2(G651), .ZN(G166));
  NAND2_X1  g091(.A1(KEYINPUT67), .A2(G651), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(KEYINPUT67), .A2(KEYINPUT6), .A3(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n519), .A2(new_n520), .B1(new_n509), .B2(new_n510), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G89), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n524), .A2(new_n525), .B1(new_n511), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n508), .B1(new_n519), .B2(new_n520), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n522), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT69), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT69), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n500), .A2(new_n501), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n537), .A2(G651), .B1(new_n521), .B2(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n528), .A2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G651), .ZN(new_n543));
  OR3_X1    g118(.A1(new_n542), .A2(KEYINPUT70), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(KEYINPUT70), .B1(new_n542), .B2(new_n543), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT71), .B(G43), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n521), .A2(G81), .B1(new_n528), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n535), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n521), .A2(G91), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n528), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT9), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n528), .A2(new_n564), .A3(G53), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n560), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  NAND2_X1  g144(.A1(new_n519), .A2(new_n520), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n570), .A2(G87), .A3(new_n511), .ZN(new_n571));
  OAI211_X1 g146(.A(G49), .B(G543), .C1(new_n497), .C2(new_n498), .ZN(new_n572));
  INV_X1    g147(.A(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n509), .A2(new_n573), .A3(new_n510), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n571), .A2(new_n572), .A3(new_n575), .ZN(G288));
  AOI22_X1  g151(.A1(new_n521), .A2(G86), .B1(new_n528), .B2(G48), .ZN(new_n577));
  OAI21_X1  g152(.A(G61), .B1(new_n500), .B2(new_n501), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n578), .A2(new_n579), .B1(G73), .B2(G543), .ZN(new_n580));
  OAI211_X1 g155(.A(KEYINPUT72), .B(G61), .C1(new_n500), .C2(new_n501), .ZN(new_n581));
  AOI211_X1 g156(.A(KEYINPUT73), .B(new_n543), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT73), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n578), .A2(new_n579), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n584), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n583), .B1(new_n586), .B2(G651), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n577), .B1(new_n582), .B2(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(new_n521), .A2(G85), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n528), .A2(G47), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n589), .B(new_n590), .C1(new_n543), .C2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(G301), .A2(G868), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n521), .A2(G92), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT74), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(G79), .ZN(new_n598));
  OR3_X1    g173(.A1(new_n598), .A2(new_n508), .A3(KEYINPUT75), .ZN(new_n599));
  OAI21_X1  g174(.A(KEYINPUT75), .B1(new_n598), .B2(new_n508), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI211_X1 g176(.A(new_n599), .B(new_n600), .C1(new_n601), .C2(new_n535), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n595), .A2(new_n596), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n593), .B1(new_n606), .B2(G868), .ZN(G284));
  XNOR2_X1  g182(.A(G284), .B(KEYINPUT76), .ZN(G321));
  NOR2_X1   g183(.A1(G299), .A2(G868), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n609), .B1(G168), .B2(G868), .ZN(G297));
  XOR2_X1   g185(.A(G297), .B(KEYINPUT77), .Z(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n606), .B1(new_n612), .B2(G860), .ZN(G148));
  NOR2_X1   g188(.A1(new_n549), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n612), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT78), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g193(.A1(new_n474), .A2(new_n476), .A3(new_n462), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT80), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n481), .A2(G123), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n467), .A2(G135), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n471), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n622), .B2(new_n623), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n625), .A2(new_n632), .ZN(G156));
  XOR2_X1   g208(.A(KEYINPUT15), .B(G2435), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2438), .ZN(new_n635));
  XOR2_X1   g210(.A(G2427), .B(G2430), .Z(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT81), .B(KEYINPUT14), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n635), .A2(new_n636), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT82), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(G14), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n644), .B2(new_n647), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n648), .A2(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT83), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g230(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n653), .A2(new_n654), .ZN(new_n657));
  AOI21_X1  g232(.A(KEYINPUT18), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2100), .ZN(new_n659));
  NOR2_X1   g234(.A1(G2072), .A2(G2078), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n442), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n655), .B2(KEYINPUT18), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(G2096), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n659), .B(new_n663), .ZN(G227));
  XNOR2_X1  g239(.A(G1981), .B(G1986), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n671), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n674), .A2(new_n673), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n674), .A2(KEYINPUT20), .A3(new_n673), .ZN(new_n679));
  OAI221_X1 g254(.A(new_n675), .B1(new_n673), .B2(new_n671), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT85), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT86), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  AND3_X1   g263(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n688), .B1(new_n684), .B2(new_n685), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n666), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n684), .A2(new_n685), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(new_n687), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n684), .A2(new_n685), .A3(new_n688), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(new_n665), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(new_n695), .ZN(G229));
  INV_X1    g271(.A(KEYINPUT102), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT90), .ZN(new_n698));
  INV_X1    g273(.A(G1971), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G22), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n699), .B(new_n701), .C1(G166), .C2(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n505), .A2(KEYINPUT68), .B1(G75), .B2(G543), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n543), .B1(new_n704), .B2(new_n513), .ZN(new_n705));
  OAI21_X1  g280(.A(G16), .B1(new_n705), .B2(new_n504), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n699), .B1(new_n706), .B2(new_n701), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n698), .B1(new_n703), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(G288), .A2(G16), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n700), .A2(G23), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(KEYINPUT33), .ZN(new_n712));
  INV_X1    g287(.A(G1976), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT33), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n709), .A2(new_n714), .A3(new_n710), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n714), .B1(new_n709), .B2(new_n710), .ZN(new_n717));
  INV_X1    g292(.A(new_n710), .ZN(new_n718));
  AOI211_X1 g293(.A(KEYINPUT33), .B(new_n718), .C1(G288), .C2(G16), .ZN(new_n719));
  OAI21_X1  g294(.A(G1976), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n515), .A2(G651), .ZN(new_n722));
  INV_X1    g297(.A(new_n504), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n700), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n701), .ZN(new_n725));
  OAI21_X1  g300(.A(G1971), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n726), .A2(KEYINPUT90), .A3(new_n702), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n708), .A2(new_n721), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT89), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT32), .B(G1981), .ZN(new_n730));
  NAND2_X1  g305(.A1(G305), .A2(G16), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n700), .A2(G6), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n732), .ZN(new_n734));
  INV_X1    g309(.A(new_n730), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n734), .B(new_n735), .C1(G305), .C2(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n729), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n577), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n586), .A2(G651), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(KEYINPUT73), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n586), .A2(new_n583), .A3(G651), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n732), .B1(new_n742), .B2(new_n700), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(new_n735), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n731), .A2(new_n732), .A3(new_n730), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n744), .A2(new_n745), .A3(KEYINPUT89), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n728), .A2(new_n737), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(KEYINPUT91), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT91), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n728), .A2(new_n737), .A3(new_n746), .A4(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n748), .A2(KEYINPUT34), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n748), .A2(KEYINPUT92), .A3(KEYINPUT34), .A4(new_n750), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(KEYINPUT34), .B1(new_n748), .B2(new_n750), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n481), .A2(G119), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT88), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n467), .A2(G131), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n471), .A2(G107), .ZN(new_n760));
  OAI21_X1  g335(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n758), .B(new_n759), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(KEYINPUT87), .B(G29), .Z(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  MUX2_X1   g339(.A(G25), .B(new_n762), .S(new_n764), .Z(new_n765));
  XOR2_X1   g340(.A(KEYINPUT35), .B(G1991), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G24), .B(G290), .S(G16), .Z(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G1986), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n756), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n755), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(KEYINPUT36), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n755), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n606), .A2(G16), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G4), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n777), .B(G1348), .C1(G4), .C2(G16), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n700), .A2(G19), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n549), .B2(new_n700), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(G1341), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n763), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n467), .A2(G140), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n481), .A2(G128), .ZN(new_n788));
  OR2_X1    g363(.A1(G104), .A2(G2105), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n789), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(G29), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n786), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G2067), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n780), .A2(new_n781), .A3(new_n784), .A4(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT93), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(G162), .A2(new_n764), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n764), .A2(G35), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT29), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n804), .A2(G2090), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT101), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(G2090), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT31), .B(G11), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT98), .Z(new_n809));
  INV_X1    g384(.A(G28), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(KEYINPUT30), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT30), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n793), .B1(new_n812), .B2(G28), .ZN(new_n813));
  OAI221_X1 g388(.A(new_n809), .B1(new_n811), .B2(new_n813), .C1(new_n630), .C2(new_n763), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n700), .A2(G5), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G301), .B2(G16), .ZN(new_n816));
  INV_X1    g391(.A(G1961), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(KEYINPUT96), .B1(G29), .B2(G32), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n467), .A2(G141), .B1(G105), .B2(new_n462), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n481), .A2(G129), .ZN(new_n821));
  NAND3_X1  g396(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT26), .Z(new_n823));
  AND3_X1   g398(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G29), .ZN(new_n825));
  MUX2_X1   g400(.A(KEYINPUT96), .B(new_n819), .S(new_n825), .Z(new_n826));
  XOR2_X1   g401(.A(KEYINPUT27), .B(G1996), .Z(new_n827));
  AND2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n807), .B(new_n818), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n700), .A2(G21), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G168), .B2(new_n700), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n764), .A2(G27), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(G164), .B2(new_n764), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G2078), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT100), .ZN(new_n836));
  OAI22_X1  g411(.A1(G1966), .A2(new_n832), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n806), .A2(new_n830), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n793), .A2(G33), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n474), .A2(G127), .A3(new_n476), .ZN(new_n840));
  INV_X1    g415(.A(G115), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n841), .B2(new_n461), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G2105), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n467), .A2(G139), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT94), .B(KEYINPUT25), .Z(new_n845));
  NAND3_X1  g420(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n843), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT95), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n839), .B1(new_n849), .B2(new_n793), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(G2072), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n832), .A2(G1966), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT97), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n700), .A2(G20), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT23), .Z(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G299), .B2(G16), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(G1956), .Z(new_n857));
  NOR2_X1   g432(.A1(new_n816), .A2(new_n817), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT99), .ZN(new_n859));
  NAND2_X1  g434(.A1(G160), .A2(G29), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT24), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(G34), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(G34), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n763), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G2084), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n835), .A2(new_n836), .ZN(new_n868));
  NOR4_X1   g443(.A1(new_n857), .A2(new_n859), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n838), .A2(new_n851), .A3(new_n853), .A4(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n797), .A2(new_n798), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n799), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n697), .B1(new_n776), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n755), .A2(new_n774), .A3(new_n771), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n774), .B1(new_n755), .B2(new_n771), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n697), .B(new_n872), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n873), .A2(new_n877), .ZN(G311));
  NAND2_X1  g453(.A1(new_n776), .A2(new_n872), .ZN(G150));
  NAND2_X1  g454(.A1(new_n606), .A2(G559), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT38), .ZN(new_n881));
  AOI22_X1  g456(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n882));
  INV_X1    g457(.A(G93), .ZN(new_n883));
  OAI22_X1  g458(.A1(new_n882), .A2(new_n543), .B1(new_n883), .B2(new_n502), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n528), .A2(G55), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n548), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n881), .B(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n889), .A2(KEYINPUT39), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n889), .A2(KEYINPUT39), .ZN(new_n891));
  NOR3_X1   g466(.A1(new_n890), .A2(new_n891), .A3(G860), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n886), .A2(G860), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT37), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n892), .A2(new_n894), .ZN(G145));
  XNOR2_X1  g470(.A(new_n762), .B(KEYINPUT104), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n620), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n849), .B(new_n824), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n792), .B(G164), .ZN(new_n900));
  AOI22_X1  g475(.A1(G130), .A2(new_n481), .B1(new_n467), .B2(G142), .ZN(new_n901));
  OAI21_X1  g476(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n903));
  INV_X1    g478(.A(G118), .ZN(new_n904));
  AOI22_X1  g479(.A1(new_n902), .A2(new_n903), .B1(new_n904), .B2(G2105), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n903), .B2(new_n902), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n901), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n900), .B(new_n907), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n899), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n899), .A2(new_n908), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XOR2_X1   g486(.A(G162), .B(new_n630), .Z(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(G160), .Z(new_n913));
  AOI21_X1  g488(.A(G37), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n913), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n909), .A2(new_n915), .A3(new_n910), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n914), .A2(KEYINPUT40), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT40), .B1(new_n914), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(G395));
  NAND2_X1  g494(.A1(new_n604), .A2(new_n605), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(new_n566), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT41), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n920), .B(G299), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT41), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n615), .B(new_n888), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n615), .B(new_n887), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n930), .B1(new_n923), .B2(new_n925), .ZN(new_n931));
  OAI21_X1  g506(.A(KEYINPUT105), .B1(new_n928), .B2(new_n924), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT42), .ZN(new_n934));
  XNOR2_X1  g509(.A(G305), .B(G290), .ZN(new_n935));
  INV_X1    g510(.A(G288), .ZN(new_n936));
  XNOR2_X1  g511(.A(G166), .B(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n935), .B(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n929), .B(new_n940), .C1(new_n931), .C2(new_n932), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n934), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n939), .B1(new_n934), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(G868), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n886), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(G868), .B2(new_n945), .ZN(G295));
  OAI21_X1  g521(.A(new_n944), .B1(G868), .B2(new_n945), .ZN(G331));
  XNOR2_X1  g522(.A(G168), .B(G301), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(new_n888), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n921), .A2(KEYINPUT106), .A3(new_n922), .ZN(new_n950));
  OAI211_X1 g525(.A(new_n949), .B(new_n950), .C1(new_n926), .C2(KEYINPUT106), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n949), .A2(new_n924), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n939), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n948), .B(new_n887), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n957), .B1(new_n923), .B2(new_n925), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(new_n952), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n938), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n955), .A2(new_n956), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n939), .B1(new_n958), .B2(new_n952), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n963), .B2(new_n956), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n955), .A2(KEYINPUT43), .A3(new_n960), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT43), .B1(new_n960), .B2(new_n962), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT44), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n969), .ZN(G397));
  NAND2_X1  g545(.A1(G160), .A2(G40), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(G164), .B2(G1384), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT107), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n791), .B(new_n795), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT108), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(new_n824), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(new_n977), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(G1996), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n982));
  INV_X1    g557(.A(new_n974), .ZN(new_n983));
  OR2_X1    g558(.A1(new_n983), .A2(G1996), .ZN(new_n984));
  OAI22_X1  g559(.A1(new_n979), .A2(new_n981), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(new_n766), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n762), .B(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n985), .B1(new_n987), .B2(new_n975), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n983), .A2(G1986), .A3(G290), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n989), .B(KEYINPUT48), .Z(new_n990));
  AND2_X1   g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n984), .B(KEYINPUT46), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n979), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT47), .Z(new_n994));
  OR2_X1    g569(.A1(new_n762), .A2(new_n986), .ZN(new_n995));
  OAI22_X1  g570(.A1(new_n985), .A2(new_n995), .B1(G2067), .B2(new_n791), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n991), .B(new_n994), .C1(new_n975), .C2(new_n996), .ZN(new_n997));
  OR2_X1    g572(.A1(G305), .A2(G1981), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n739), .A2(new_n577), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(G1981), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(KEYINPUT49), .A3(new_n1000), .ZN(new_n1004));
  INV_X1    g579(.A(G8), .ZN(new_n1005));
  INV_X1    g580(.A(G40), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n470), .A2(new_n479), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G164), .A2(G1384), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1005), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1003), .A2(new_n1004), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1009), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(KEYINPUT112), .A3(new_n1004), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1009), .A2(new_n713), .A3(G288), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n936), .B2(G1976), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1018), .A2(new_n1009), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1009), .A2(new_n1020), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1016), .A2(new_n1017), .A3(new_n1022), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1012), .A2(new_n1015), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G164), .ZN(new_n1025));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(KEYINPUT45), .A3(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n1007), .A3(new_n973), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n699), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1025), .A2(new_n1030), .A3(new_n1026), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n1007), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1029), .B1(G2090), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(G8), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1036));
  NAND3_X1  g611(.A1(G303), .A2(G8), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT110), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1036), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(G166), .B2(new_n1005), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1037), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1038), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1035), .A2(new_n1043), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n1035), .B2(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1031), .A2(new_n1007), .A3(new_n1032), .ZN(new_n1047));
  INV_X1    g622(.A(G1966), .ZN(new_n1048));
  AOI22_X1  g623(.A1(new_n1047), .A2(new_n866), .B1(new_n1028), .B2(new_n1048), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1049), .A2(new_n1005), .A3(G286), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1024), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT63), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1024), .A2(new_n1046), .A3(KEYINPUT63), .A4(new_n1050), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G288), .A2(G1976), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1014), .A2(KEYINPUT112), .A3(new_n1004), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT112), .B1(new_n1014), .B2(new_n1004), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1013), .B1(new_n1059), .B2(new_n998), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1061), .B(new_n1044), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1060), .A2(new_n1063), .A3(KEYINPUT113), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1056), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1066), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1067));
  INV_X1    g642(.A(new_n998), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1009), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1065), .B1(new_n1069), .B2(new_n1062), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1055), .B1(new_n1064), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1028), .A2(new_n1048), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1031), .A2(new_n1007), .A3(new_n1032), .A4(new_n866), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1005), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(G168), .A2(new_n1005), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT51), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT121), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1049), .B2(new_n1005), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1074), .A2(KEYINPUT122), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1075), .A2(KEYINPUT51), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1083), .B(KEYINPUT51), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1077), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n1086));
  OR3_X1    g661(.A1(new_n1049), .A2(new_n1005), .A3(G168), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1028), .A2(G2078), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1091), .A2(KEYINPUT123), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(KEYINPUT123), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n817), .B2(new_n1033), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1086), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1088), .B(new_n1097), .C1(new_n1098), .C2(KEYINPUT126), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1098), .A2(KEYINPUT126), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n560), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n558), .A2(KEYINPUT117), .A3(new_n559), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n563), .A2(new_n1104), .A3(new_n565), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1104), .B1(new_n563), .B2(new_n565), .ZN(new_n1107));
  OAI21_X1  g682(.A(KEYINPUT115), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n566), .A2(new_n1109), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT114), .B(G1956), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n1033), .A2(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT56), .B(G2072), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1027), .A2(new_n1007), .A3(new_n973), .A4(new_n1117), .ZN(new_n1118));
  AND4_X1   g693(.A1(new_n1110), .A2(new_n1114), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1110), .A2(new_n1114), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1123));
  OAI22_X1  g698(.A1(new_n1047), .A2(G1348), .B1(G2067), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n606), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1119), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n1127));
  OR3_X1    g702(.A1(new_n1124), .A2(new_n606), .A3(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n606), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1128), .A2(new_n1129), .B1(new_n1127), .B2(new_n1124), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT119), .B1(new_n1131), .B2(KEYINPUT59), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(KEYINPUT58), .B(G1341), .Z(new_n1134));
  NAND2_X1  g709(.A1(new_n1123), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1135), .B1(new_n1028), .B2(G1996), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1136), .B2(new_n549), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1136), .A2(new_n549), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1132), .B1(KEYINPUT119), .B2(KEYINPUT59), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1110), .A2(new_n1114), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1141), .B1(new_n1119), .B2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1110), .A2(new_n1114), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1122), .A2(KEYINPUT61), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1140), .A2(new_n1143), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1130), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1140), .A2(new_n1143), .A3(KEYINPUT120), .A4(new_n1145), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1126), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1096), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1151));
  XNOR2_X1  g726(.A(G301), .B(KEYINPUT54), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1033), .A2(new_n817), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT124), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1154), .A2(new_n1152), .A3(new_n1095), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1151), .A2(new_n1152), .B1(new_n1094), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n1099), .A2(new_n1100), .B1(new_n1150), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1024), .A2(new_n1046), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n1160), .B(KEYINPUT125), .Z(new_n1161));
  AOI21_X1  g736(.A(new_n1071), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  XOR2_X1   g737(.A(G290), .B(G1986), .Z(new_n1163));
  OAI21_X1  g738(.A(new_n988), .B1(new_n983), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n997), .B1(new_n1162), .B2(new_n1164), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g740(.A(G319), .ZN(new_n1167));
  AOI211_X1 g741(.A(new_n1167), .B(G227), .C1(new_n648), .C2(new_n650), .ZN(new_n1168));
  NAND3_X1  g742(.A1(new_n691), .A2(new_n695), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g743(.A1(new_n1169), .A2(KEYINPUT127), .ZN(new_n1170));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n1171));
  NAND4_X1  g745(.A1(new_n691), .A2(new_n695), .A3(new_n1171), .A4(new_n1168), .ZN(new_n1172));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n914), .A2(new_n916), .ZN(new_n1174));
  AND3_X1   g748(.A1(new_n1173), .A2(new_n964), .A3(new_n1174), .ZN(G308));
  NAND3_X1  g749(.A1(new_n1173), .A2(new_n964), .A3(new_n1174), .ZN(G225));
endmodule


