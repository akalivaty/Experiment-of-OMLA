

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591;

  XNOR2_X1 U324 ( .A(n345), .B(n344), .ZN(n346) );
  NAND2_X1 U325 ( .A1(n539), .A2(n550), .ZN(n292) );
  INV_X1 U326 ( .A(KEYINPUT45), .ZN(n336) );
  XNOR2_X1 U327 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U328 ( .A(n304), .B(n303), .ZN(n307) );
  XNOR2_X1 U329 ( .A(n347), .B(n346), .ZN(n349) );
  XOR2_X1 U330 ( .A(G176GAT), .B(G64GAT), .Z(n389) );
  INV_X1 U331 ( .A(n350), .ZN(n297) );
  XNOR2_X1 U332 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n382) );
  XNOR2_X1 U333 ( .A(n298), .B(n297), .ZN(n311) );
  XNOR2_X1 U334 ( .A(n311), .B(n310), .ZN(n318) );
  OR2_X1 U335 ( .A1(n292), .A2(n461), .ZN(n462) );
  XNOR2_X1 U336 ( .A(n458), .B(G176GAT), .ZN(n459) );
  XNOR2_X1 U337 ( .A(n460), .B(n459), .ZN(G1349GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT81), .B(G92GAT), .Z(n294) );
  XNOR2_X1 U339 ( .A(G190GAT), .B(G218GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U341 ( .A(G36GAT), .B(n295), .Z(n390) );
  XNOR2_X1 U342 ( .A(n390), .B(KEYINPUT66), .ZN(n298) );
  XNOR2_X1 U343 ( .A(G99GAT), .B(G106GAT), .ZN(n296) );
  XNOR2_X1 U344 ( .A(n296), .B(KEYINPUT74), .ZN(n350) );
  XOR2_X1 U345 ( .A(KEYINPUT10), .B(KEYINPUT79), .Z(n300) );
  XNOR2_X1 U346 ( .A(KEYINPUT80), .B(KEYINPUT11), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n304) );
  NAND2_X1 U348 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  INV_X1 U349 ( .A(KEYINPUT78), .ZN(n301) );
  INV_X1 U350 ( .A(n307), .ZN(n305) );
  NAND2_X1 U351 ( .A1(n305), .A2(KEYINPUT9), .ZN(n309) );
  INV_X1 U352 ( .A(KEYINPUT9), .ZN(n306) );
  NAND2_X1 U353 ( .A1(n307), .A2(n306), .ZN(n308) );
  NAND2_X1 U354 ( .A1(n309), .A2(n308), .ZN(n310) );
  XOR2_X1 U355 ( .A(KEYINPUT72), .B(KEYINPUT7), .Z(n313) );
  XNOR2_X1 U356 ( .A(G50GAT), .B(G43GAT), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U358 ( .A(KEYINPUT8), .B(n314), .Z(n368) );
  XOR2_X1 U359 ( .A(G85GAT), .B(G162GAT), .Z(n316) );
  XNOR2_X1 U360 ( .A(G29GAT), .B(G134GAT), .ZN(n315) );
  XNOR2_X1 U361 ( .A(n316), .B(n315), .ZN(n411) );
  XNOR2_X1 U362 ( .A(n368), .B(n411), .ZN(n317) );
  XNOR2_X1 U363 ( .A(n318), .B(n317), .ZN(n566) );
  XOR2_X1 U364 ( .A(KEYINPUT82), .B(n566), .Z(n550) );
  XOR2_X1 U365 ( .A(KEYINPUT36), .B(n550), .Z(n587) );
  XOR2_X1 U366 ( .A(KEYINPUT83), .B(KEYINPUT12), .Z(n320) );
  XNOR2_X1 U367 ( .A(G8GAT), .B(KEYINPUT14), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n335) );
  XOR2_X1 U369 ( .A(G183GAT), .B(G211GAT), .Z(n384) );
  XOR2_X1 U370 ( .A(G64GAT), .B(KEYINPUT13), .Z(n322) );
  XNOR2_X1 U371 ( .A(G1GAT), .B(G57GAT), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U373 ( .A(n384), .B(n323), .Z(n325) );
  NAND2_X1 U374 ( .A1(G231GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U375 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U376 ( .A(KEYINPUT15), .B(KEYINPUT85), .Z(n327) );
  XNOR2_X1 U377 ( .A(KEYINPUT84), .B(KEYINPUT86), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U379 ( .A(n329), .B(n328), .Z(n333) );
  XNOR2_X1 U380 ( .A(G15GAT), .B(G127GAT), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n330), .B(G71GAT), .ZN(n453) );
  XNOR2_X1 U382 ( .A(G22GAT), .B(G155GAT), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n331), .B(G78GAT), .ZN(n421) );
  XNOR2_X1 U384 ( .A(n453), .B(n421), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n584) );
  OR2_X1 U387 ( .A1(n587), .A2(n584), .ZN(n337) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n373) );
  XOR2_X1 U389 ( .A(G204GAT), .B(G78GAT), .Z(n339) );
  XNOR2_X1 U390 ( .A(G71GAT), .B(G120GAT), .ZN(n338) );
  XOR2_X1 U391 ( .A(n339), .B(n338), .Z(n354) );
  XOR2_X1 U392 ( .A(G92GAT), .B(n389), .Z(n341) );
  XOR2_X1 U393 ( .A(G148GAT), .B(G57GAT), .Z(n403) );
  XNOR2_X1 U394 ( .A(G85GAT), .B(n403), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n347) );
  XOR2_X1 U396 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n343) );
  XNOR2_X1 U397 ( .A(KEYINPUT33), .B(KEYINPUT13), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n345) );
  AND2_X1 U399 ( .A1(G230GAT), .A2(G233GAT), .ZN(n344) );
  INV_X1 U400 ( .A(KEYINPUT32), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n349), .B(n348), .ZN(n352) );
  XNOR2_X1 U402 ( .A(n350), .B(KEYINPUT76), .ZN(n351) );
  XNOR2_X1 U403 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n580) );
  XOR2_X1 U405 ( .A(KEYINPUT70), .B(G15GAT), .Z(n356) );
  XNOR2_X1 U406 ( .A(G22GAT), .B(G197GAT), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U408 ( .A(n357), .B(G36GAT), .Z(n359) );
  XOR2_X1 U409 ( .A(G169GAT), .B(G8GAT), .Z(n385) );
  XNOR2_X1 U410 ( .A(n385), .B(G29GAT), .ZN(n358) );
  XNOR2_X1 U411 ( .A(n359), .B(n358), .ZN(n364) );
  XNOR2_X1 U412 ( .A(G141GAT), .B(G113GAT), .ZN(n360) );
  XNOR2_X1 U413 ( .A(n360), .B(G1GAT), .ZN(n400) );
  XOR2_X1 U414 ( .A(n400), .B(KEYINPUT68), .Z(n362) );
  NAND2_X1 U415 ( .A1(G229GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U417 ( .A(n364), .B(n363), .Z(n370) );
  XOR2_X1 U418 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n366) );
  XNOR2_X1 U419 ( .A(KEYINPUT30), .B(KEYINPUT71), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U421 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U422 ( .A(n370), .B(n369), .ZN(n576) );
  XNOR2_X1 U423 ( .A(n576), .B(KEYINPUT73), .ZN(n568) );
  INV_X1 U424 ( .A(n568), .ZN(n371) );
  AND2_X1 U425 ( .A1(n580), .A2(n371), .ZN(n372) );
  AND2_X1 U426 ( .A1(n373), .A2(n372), .ZN(n381) );
  XOR2_X1 U427 ( .A(n584), .B(KEYINPUT114), .Z(n572) );
  XOR2_X1 U428 ( .A(KEYINPUT46), .B(KEYINPUT115), .Z(n375) );
  XOR2_X1 U429 ( .A(KEYINPUT41), .B(n580), .Z(n559) );
  NOR2_X1 U430 ( .A1(n559), .A2(n576), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n376) );
  NOR2_X1 U432 ( .A1(n572), .A2(n376), .ZN(n377) );
  AND2_X1 U433 ( .A1(n377), .A2(n566), .ZN(n379) );
  INV_X1 U434 ( .A(KEYINPUT47), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n380) );
  NOR2_X1 U436 ( .A1(n381), .A2(n380), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n383), .B(n382), .ZN(n538) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n396) );
  XNOR2_X1 U439 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n386), .B(KEYINPUT18), .ZN(n451) );
  XOR2_X1 U441 ( .A(G204GAT), .B(KEYINPUT93), .Z(n388) );
  XNOR2_X1 U442 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n420) );
  XNOR2_X1 U444 ( .A(n451), .B(n420), .ZN(n394) );
  XOR2_X1 U445 ( .A(n390), .B(n389), .Z(n392) );
  NAND2_X1 U446 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U447 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n396), .B(n395), .ZN(n526) );
  XNOR2_X1 U450 ( .A(n526), .B(KEYINPUT122), .ZN(n397) );
  NOR2_X1 U451 ( .A1(n538), .A2(n397), .ZN(n398) );
  XNOR2_X1 U452 ( .A(n398), .B(KEYINPUT54), .ZN(n416) );
  XNOR2_X1 U453 ( .A(KEYINPUT94), .B(KEYINPUT3), .ZN(n399) );
  XNOR2_X1 U454 ( .A(n399), .B(KEYINPUT2), .ZN(n428) );
  XNOR2_X1 U455 ( .A(n400), .B(n428), .ZN(n415) );
  XOR2_X1 U456 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n402) );
  XNOR2_X1 U457 ( .A(KEYINPUT6), .B(KEYINPUT4), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n407) );
  XOR2_X1 U459 ( .A(n403), .B(G155GAT), .Z(n405) );
  XOR2_X1 U460 ( .A(KEYINPUT0), .B(G120GAT), .Z(n444) );
  XNOR2_X1 U461 ( .A(G127GAT), .B(n444), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U463 ( .A(n407), .B(n406), .Z(n409) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U466 ( .A(n410), .B(KEYINPUT97), .Z(n413) );
  XNOR2_X1 U467 ( .A(n411), .B(KEYINPUT98), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n476) );
  XNOR2_X1 U470 ( .A(KEYINPUT99), .B(n476), .ZN(n523) );
  NAND2_X1 U471 ( .A1(n416), .A2(n523), .ZN(n417) );
  XNOR2_X1 U472 ( .A(n417), .B(KEYINPUT64), .ZN(n575) );
  XOR2_X1 U473 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n419) );
  XNOR2_X1 U474 ( .A(G148GAT), .B(KEYINPUT92), .ZN(n418) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(n437) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n435) );
  XOR2_X1 U477 ( .A(KEYINPUT95), .B(G106GAT), .Z(n423) );
  XNOR2_X1 U478 ( .A(G162GAT), .B(KEYINPUT78), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U480 ( .A(G211GAT), .B(KEYINPUT96), .Z(n425) );
  XNOR2_X1 U481 ( .A(G141GAT), .B(KEYINPUT24), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U483 ( .A(n427), .B(n426), .Z(n433) );
  XOR2_X1 U484 ( .A(n428), .B(G218GAT), .Z(n430) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U487 ( .A(G50GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n479) );
  NOR2_X1 U491 ( .A1(n575), .A2(n479), .ZN(n438) );
  XNOR2_X1 U492 ( .A(n438), .B(KEYINPUT55), .ZN(n461) );
  XOR2_X1 U493 ( .A(KEYINPUT65), .B(KEYINPUT20), .Z(n440) );
  XNOR2_X1 U494 ( .A(KEYINPUT88), .B(G183GAT), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n448) );
  XOR2_X1 U496 ( .A(KEYINPUT89), .B(KEYINPUT90), .Z(n442) );
  XNOR2_X1 U497 ( .A(G190GAT), .B(G99GAT), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U499 ( .A(n443), .B(G134GAT), .Z(n446) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U502 ( .A(n448), .B(n447), .ZN(n457) );
  XOR2_X1 U503 ( .A(G176GAT), .B(G113GAT), .Z(n450) );
  NAND2_X1 U504 ( .A1(G227GAT), .A2(G233GAT), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n452) );
  XOR2_X1 U506 ( .A(n452), .B(n451), .Z(n455) );
  XNOR2_X1 U507 ( .A(G169GAT), .B(n453), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U509 ( .A(n457), .B(n456), .Z(n539) );
  INV_X1 U510 ( .A(n539), .ZN(n529) );
  NOR2_X1 U511 ( .A1(n461), .A2(n529), .ZN(n571) );
  INV_X1 U512 ( .A(n559), .ZN(n544) );
  NAND2_X1 U513 ( .A1(n571), .A2(n544), .ZN(n460) );
  XOR2_X1 U514 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n458) );
  INV_X1 U515 ( .A(G190GAT), .ZN(n465) );
  XOR2_X1 U516 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n463) );
  XNOR2_X1 U517 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U518 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  NAND2_X1 U519 ( .A1(n568), .A2(n580), .ZN(n466) );
  XOR2_X1 U520 ( .A(KEYINPUT77), .B(n466), .Z(n500) );
  OR2_X1 U521 ( .A1(n550), .A2(n584), .ZN(n467) );
  XNOR2_X1 U522 ( .A(n467), .B(KEYINPUT87), .ZN(n468) );
  XNOR2_X1 U523 ( .A(n468), .B(KEYINPUT16), .ZN(n486) );
  NOR2_X1 U524 ( .A1(n529), .A2(n526), .ZN(n469) );
  NOR2_X1 U525 ( .A1(n479), .A2(n469), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT25), .B(n470), .Z(n474) );
  XNOR2_X1 U527 ( .A(n526), .B(KEYINPUT27), .ZN(n480) );
  XOR2_X1 U528 ( .A(KEYINPUT101), .B(KEYINPUT26), .Z(n472) );
  NAND2_X1 U529 ( .A1(n529), .A2(n479), .ZN(n471) );
  XOR2_X1 U530 ( .A(n472), .B(n471), .Z(n556) );
  INV_X1 U531 ( .A(n556), .ZN(n574) );
  NOR2_X1 U532 ( .A1(n480), .A2(n574), .ZN(n473) );
  NOR2_X1 U533 ( .A1(n474), .A2(n473), .ZN(n475) );
  NOR2_X1 U534 ( .A1(n476), .A2(n475), .ZN(n477) );
  XOR2_X1 U535 ( .A(KEYINPUT102), .B(n477), .Z(n485) );
  XOR2_X1 U536 ( .A(KEYINPUT91), .B(n529), .Z(n483) );
  XOR2_X1 U537 ( .A(KEYINPUT67), .B(KEYINPUT28), .Z(n478) );
  XOR2_X1 U538 ( .A(n479), .B(n478), .Z(n534) );
  INV_X1 U539 ( .A(n534), .ZN(n542) );
  NOR2_X1 U540 ( .A1(n523), .A2(n480), .ZN(n481) );
  XOR2_X1 U541 ( .A(KEYINPUT100), .B(n481), .Z(n537) );
  NOR2_X1 U542 ( .A1(n542), .A2(n537), .ZN(n482) );
  NAND2_X1 U543 ( .A1(n483), .A2(n482), .ZN(n484) );
  NAND2_X1 U544 ( .A1(n485), .A2(n484), .ZN(n497) );
  NAND2_X1 U545 ( .A1(n486), .A2(n497), .ZN(n512) );
  OR2_X1 U546 ( .A1(n500), .A2(n512), .ZN(n494) );
  NOR2_X1 U547 ( .A1(n523), .A2(n494), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT34), .B(KEYINPUT103), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(n489), .ZN(G1324GAT) );
  NOR2_X1 U551 ( .A1(n526), .A2(n494), .ZN(n490) );
  XOR2_X1 U552 ( .A(G8GAT), .B(n490), .Z(G1325GAT) );
  NOR2_X1 U553 ( .A1(n529), .A2(n494), .ZN(n492) );
  XNOR2_X1 U554 ( .A(KEYINPUT35), .B(KEYINPUT104), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U556 ( .A(G15GAT), .B(n493), .ZN(G1326GAT) );
  NOR2_X1 U557 ( .A1(n534), .A2(n494), .ZN(n496) );
  XNOR2_X1 U558 ( .A(G22GAT), .B(KEYINPUT105), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(G1327GAT) );
  NAND2_X1 U560 ( .A1(n584), .A2(n497), .ZN(n498) );
  NOR2_X1 U561 ( .A1(n587), .A2(n498), .ZN(n499) );
  XNOR2_X1 U562 ( .A(KEYINPUT37), .B(n499), .ZN(n522) );
  NOR2_X1 U563 ( .A1(n522), .A2(n500), .ZN(n502) );
  XOR2_X1 U564 ( .A(KEYINPUT38), .B(KEYINPUT106), .Z(n501) );
  XNOR2_X1 U565 ( .A(n502), .B(n501), .ZN(n509) );
  NOR2_X1 U566 ( .A1(n523), .A2(n509), .ZN(n504) );
  XNOR2_X1 U567 ( .A(KEYINPUT107), .B(KEYINPUT39), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U569 ( .A(G29GAT), .B(n505), .Z(G1328GAT) );
  NOR2_X1 U570 ( .A1(n526), .A2(n509), .ZN(n506) );
  XOR2_X1 U571 ( .A(G36GAT), .B(n506), .Z(G1329GAT) );
  NOR2_X1 U572 ( .A1(n529), .A2(n509), .ZN(n507) );
  XOR2_X1 U573 ( .A(KEYINPUT40), .B(n507), .Z(n508) );
  XNOR2_X1 U574 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NOR2_X1 U575 ( .A1(n534), .A2(n509), .ZN(n510) );
  XOR2_X1 U576 ( .A(G50GAT), .B(n510), .Z(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT108), .B(n511), .ZN(G1331GAT) );
  NAND2_X1 U578 ( .A1(n576), .A2(n544), .ZN(n521) );
  OR2_X1 U579 ( .A1(n521), .A2(n512), .ZN(n517) );
  NOR2_X1 U580 ( .A1(n523), .A2(n517), .ZN(n513) );
  XOR2_X1 U581 ( .A(n513), .B(KEYINPUT42), .Z(n514) );
  XNOR2_X1 U582 ( .A(G57GAT), .B(n514), .ZN(G1332GAT) );
  NOR2_X1 U583 ( .A1(n526), .A2(n517), .ZN(n515) );
  XOR2_X1 U584 ( .A(G64GAT), .B(n515), .Z(G1333GAT) );
  NOR2_X1 U585 ( .A1(n529), .A2(n517), .ZN(n516) );
  XOR2_X1 U586 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U587 ( .A1(n534), .A2(n517), .ZN(n519) );
  XNOR2_X1 U588 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U589 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U590 ( .A(G78GAT), .B(n520), .Z(G1335GAT) );
  OR2_X1 U591 ( .A1(n522), .A2(n521), .ZN(n533) );
  NOR2_X1 U592 ( .A1(n523), .A2(n533), .ZN(n524) );
  XOR2_X1 U593 ( .A(G85GAT), .B(n524), .Z(n525) );
  XNOR2_X1 U594 ( .A(KEYINPUT110), .B(n525), .ZN(G1336GAT) );
  NOR2_X1 U595 ( .A1(n526), .A2(n533), .ZN(n528) );
  XNOR2_X1 U596 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n527) );
  XNOR2_X1 U597 ( .A(n528), .B(n527), .ZN(G1337GAT) );
  NOR2_X1 U598 ( .A1(n529), .A2(n533), .ZN(n530) );
  XOR2_X1 U599 ( .A(G99GAT), .B(n530), .Z(G1338GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n532) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(KEYINPUT112), .ZN(n531) );
  XNOR2_X1 U602 ( .A(n532), .B(n531), .ZN(n536) );
  NOR2_X1 U603 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U604 ( .A(n536), .B(n535), .Z(G1339GAT) );
  NOR2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n557) );
  NAND2_X1 U606 ( .A1(n557), .A2(n539), .ZN(n540) );
  XOR2_X1 U607 ( .A(KEYINPUT117), .B(n540), .Z(n541) );
  NOR2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n568), .A2(n551), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n543), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U612 ( .A1(n551), .A2(n544), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n548) );
  NAND2_X1 U615 ( .A1(n551), .A2(n572), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U617 ( .A(G127GAT), .B(n549), .Z(G1342GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n555) );
  XOR2_X1 U621 ( .A(G134GAT), .B(KEYINPUT119), .Z(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n565) );
  NOR2_X1 U624 ( .A1(n576), .A2(n565), .ZN(n558) );
  XOR2_X1 U625 ( .A(G141GAT), .B(n558), .Z(G1344GAT) );
  NOR2_X1 U626 ( .A1(n565), .A2(n559), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n561) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT121), .ZN(n560) );
  XNOR2_X1 U629 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U631 ( .A1(n584), .A2(n565), .ZN(n564) );
  XOR2_X1 U632 ( .A(G155GAT), .B(n564), .Z(G1346GAT) );
  NOR2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U634 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  XOR2_X1 U635 ( .A(G169GAT), .B(KEYINPUT123), .Z(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n568), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1348GAT) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  OR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n588) );
  NOR2_X1 U641 ( .A1(n576), .A2(n588), .ZN(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n579), .ZN(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n588), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(G204GAT), .B(n583), .Z(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n588), .ZN(n585) );
  XOR2_X1 U650 ( .A(KEYINPUT126), .B(n585), .Z(n586) );
  XNOR2_X1 U651 ( .A(G211GAT), .B(n586), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U653 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

