//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1190, new_n1191, new_n1192, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n214), .A2(G20), .A3(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI22_X1  g0020(.A1(new_n218), .A2(new_n219), .B1(new_n203), .B2(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n221), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G77), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT64), .B(G244), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n222), .B(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT65), .Z(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XOR2_X1   g0041(.A(G107), .B(G116), .Z(new_n242));
  XOR2_X1   g0042(.A(new_n241), .B(new_n242), .Z(new_n243));
  XOR2_X1   g0043(.A(new_n243), .B(KEYINPUT68), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G68), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n215), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT84), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT6), .ZN(new_n255));
  NOR3_X1   g0055(.A1(new_n255), .A2(new_n202), .A3(G107), .ZN(new_n256));
  XNOR2_X1  g0056(.A(G97), .B(G107), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n256), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n254), .B1(new_n207), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT7), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT3), .B(G33), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(new_n261), .B2(G20), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n267), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n203), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n251), .B1(new_n259), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G97), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(new_n215), .A3(new_n250), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n206), .B2(G33), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n272), .B1(new_n274), .B2(G97), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT5), .B(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  OAI211_X1 g0078(.A(G1), .B(G13), .C1(new_n263), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n206), .A2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n277), .A2(new_n279), .A3(G274), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n277), .A2(new_n281), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n279), .ZN(new_n284));
  INV_X1    g0084(.A(G257), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G1698), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n261), .A2(G244), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT4), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n261), .A2(KEYINPUT4), .A3(G244), .A4(new_n287), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G283), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n290), .A2(new_n291), .A3(new_n292), .A4(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n286), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n276), .B1(G169), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n295), .ZN(new_n298));
  INV_X1    g0098(.A(new_n286), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT72), .B(G179), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n300), .A2(KEYINPUT85), .A3(G200), .ZN(new_n305));
  INV_X1    g0105(.A(new_n276), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT85), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n296), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n296), .A2(G190), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n305), .A2(new_n306), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT86), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n276), .B1(G190), .B2(new_n296), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT86), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n313), .A2(new_n314), .A3(new_n305), .A4(new_n309), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n304), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n261), .A2(G222), .A3(new_n287), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT70), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n317), .B(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n267), .A2(new_n287), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(G223), .B1(G77), .B2(new_n267), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n279), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n324), .A2(new_n279), .A3(G274), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT69), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n206), .B(KEYINPUT69), .C1(G41), .C2(G45), .ZN(new_n328));
  AND3_X1   g0128(.A1(new_n327), .A2(new_n279), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n325), .B1(new_n329), .B2(G226), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n322), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT10), .B1(new_n332), .B2(G190), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT8), .B(G58), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n207), .A2(G33), .ZN(new_n335));
  INV_X1    g0135(.A(G150), .ZN(new_n336));
  INV_X1    g0136(.A(new_n252), .ZN(new_n337));
  OAI22_X1  g0137(.A1(new_n334), .A2(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(G50), .A2(G58), .ZN(new_n339));
  INV_X1    g0139(.A(G68), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n207), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n251), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n273), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n218), .B1(new_n206), .B2(G20), .ZN(new_n344));
  INV_X1    g0144(.A(new_n271), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n343), .A2(new_n344), .B1(new_n218), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n347), .A2(KEYINPUT9), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(KEYINPUT9), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT76), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(G200), .B1(new_n322), .B2(new_n331), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n348), .A2(KEYINPUT76), .A3(new_n349), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n333), .A2(new_n352), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G190), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n317), .B(KEYINPUT70), .ZN(new_n357));
  INV_X1    g0157(.A(new_n321), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n295), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n330), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n350), .B(new_n353), .C1(new_n356), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT10), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n347), .ZN(new_n364));
  INV_X1    g0164(.A(G169), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(KEYINPUT71), .B1(new_n301), .B2(new_n332), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n347), .B1(new_n332), .B2(G169), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT71), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n334), .B1(KEYINPUT75), .B2(new_n337), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(KEYINPUT75), .B2(new_n337), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT15), .B(G87), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n373), .B1(new_n207), .B2(new_n224), .C1(new_n335), .C2(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n375), .A2(new_n251), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n206), .A2(G20), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G77), .ZN(new_n378));
  OAI22_X1  g0178(.A1(new_n273), .A2(new_n378), .B1(G77), .B2(new_n271), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n324), .A2(new_n279), .A3(G274), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n327), .A2(new_n279), .A3(new_n328), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(new_n225), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT73), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G232), .A2(G1698), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n287), .A2(G238), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n261), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n389), .B(new_n295), .C1(G107), .C2(new_n261), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n384), .A2(new_n385), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n386), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT74), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n386), .A2(KEYINPUT74), .A3(new_n390), .A4(new_n391), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n365), .A3(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(new_n394), .A2(new_n395), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n381), .B(new_n396), .C1(new_n397), .C2(new_n302), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n394), .A2(G200), .A3(new_n395), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n380), .B(new_n399), .C1(new_n397), .C2(new_n356), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n363), .A2(new_n371), .A3(new_n398), .A4(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT77), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n345), .A2(new_n340), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT12), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n340), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n224), .B2(new_n335), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(KEYINPUT11), .A3(new_n251), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n343), .A2(G68), .A3(new_n377), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n405), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT11), .B1(new_n407), .B2(new_n251), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT78), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n261), .A2(G232), .A3(G1698), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n261), .A2(G226), .A3(new_n287), .ZN(new_n416));
  NAND2_X1  g0216(.A1(G33), .A2(G97), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n295), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n325), .B1(new_n329), .B2(G238), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT13), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(new_n419), .B2(new_n420), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n414), .B(G169), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n419), .A2(new_n420), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT13), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(G179), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n427), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n414), .B1(new_n430), .B2(G169), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n413), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n422), .A2(new_n423), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT14), .B1(new_n433), .B2(new_n365), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n434), .A2(KEYINPUT78), .A3(new_n428), .A4(new_n424), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n412), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(G190), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n430), .A2(G200), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(new_n438), .A3(new_n412), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n362), .A2(new_n355), .B1(new_n367), .B2(new_n370), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n442), .A2(KEYINPUT77), .A3(new_n400), .A4(new_n398), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n403), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT17), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n327), .A2(G232), .A3(new_n279), .A4(new_n328), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n382), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT80), .ZN(new_n448));
  INV_X1    g0248(.A(G87), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n263), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(G223), .A2(G1698), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n451), .B1(new_n219), .B2(G1698), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n450), .B1(new_n452), .B2(new_n261), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n448), .B1(new_n453), .B2(new_n279), .ZN(new_n454));
  INV_X1    g0254(.A(G223), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n287), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n219), .A2(G1698), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n264), .A2(new_n456), .A3(new_n266), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n450), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(KEYINPUT80), .A3(new_n295), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n447), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n356), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n453), .A2(new_n279), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n308), .B1(new_n464), .B2(new_n447), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT7), .B1(new_n267), .B2(new_n207), .ZN(new_n468));
  AOI211_X1 g0268(.A(new_n260), .B(G20), .C1(new_n264), .C2(new_n266), .ZN(new_n469));
  OAI21_X1  g0269(.A(G68), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G58), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n340), .ZN(new_n472));
  NOR2_X1   g0272(.A1(G58), .A2(G68), .ZN(new_n473));
  OAI21_X1  g0273(.A(G20), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n252), .A2(G159), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n470), .A2(KEYINPUT16), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT16), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n340), .B1(new_n262), .B2(new_n268), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(new_n476), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n481), .A3(new_n251), .ZN(new_n482));
  XOR2_X1   g0282(.A(KEYINPUT8), .B(G58), .Z(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n377), .ZN(new_n484));
  OAI22_X1  g0284(.A1(new_n484), .A2(new_n273), .B1(new_n271), .B2(new_n483), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT79), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI221_X1 g0287(.A(KEYINPUT79), .B1(new_n271), .B2(new_n483), .C1(new_n484), .C2(new_n273), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n445), .B1(new_n467), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n487), .A2(new_n488), .ZN(new_n492));
  INV_X1    g0292(.A(new_n251), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n470), .A2(new_n477), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(new_n494), .B2(new_n479), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n492), .B1(new_n495), .B2(new_n478), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(new_n466), .A3(KEYINPUT17), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT18), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n446), .A2(new_n382), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT80), .B1(new_n460), .B2(new_n295), .ZN(new_n501));
  AOI211_X1 g0301(.A(new_n448), .B(new_n279), .C1(new_n458), .C2(new_n459), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n301), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT81), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT81), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n462), .A2(new_n505), .A3(new_n301), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n365), .B1(new_n464), .B2(new_n447), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT82), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n496), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n504), .A2(new_n506), .A3(KEYINPUT82), .A4(new_n507), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n499), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n507), .B1(new_n503), .B2(KEYINPUT81), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n505), .B1(new_n462), .B2(new_n301), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND4_X1   g0315(.A1(new_n499), .A2(new_n515), .A3(new_n490), .A4(new_n511), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT83), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n490), .A3(new_n511), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT18), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n510), .A2(new_n499), .A3(new_n511), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT83), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n498), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n444), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n261), .A2(G238), .A3(new_n287), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G116), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n261), .A2(G1698), .ZN(new_n528));
  INV_X1    g0328(.A(G244), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n295), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n280), .A2(G250), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n279), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n279), .A2(G274), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n280), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n365), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n261), .A2(new_n207), .A3(G68), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT19), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n207), .B1(new_n417), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(G87), .B2(new_n204), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n335), .B2(new_n202), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(new_n251), .B1(new_n345), .B2(new_n374), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n343), .B1(G1), .B2(new_n263), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n374), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n538), .B(new_n547), .C1(new_n302), .C2(new_n537), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n274), .A2(G87), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n535), .B1(new_n530), .B2(new_n295), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G190), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n550), .B(new_n552), .C1(new_n308), .C2(new_n551), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n261), .A2(new_n207), .A3(G87), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT22), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT22), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n261), .A2(new_n557), .A3(new_n207), .A4(G87), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT24), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n527), .A2(G20), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT23), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n207), .B2(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n561), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n559), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n560), .B1(new_n559), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n251), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT25), .B1(new_n345), .B2(new_n203), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n345), .A2(KEYINPUT25), .A3(new_n203), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n274), .A2(G107), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G250), .A2(G1698), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n285), .B2(G1698), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(new_n261), .B1(G33), .B2(G294), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n295), .B1(new_n281), .B2(new_n277), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n576), .A2(new_n295), .B1(G264), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n578), .A2(G190), .A3(new_n282), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(G264), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n580), .B(new_n282), .C1(new_n279), .C2(new_n575), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G200), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n568), .A2(new_n572), .A3(new_n579), .A4(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n293), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n584));
  INV_X1    g0384(.A(G116), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G20), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n251), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT20), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n271), .A2(G116), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n274), .B2(G116), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n261), .A2(G257), .A3(new_n287), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n261), .A2(KEYINPUT87), .A3(G257), .A4(new_n287), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n320), .A2(G264), .B1(G303), .B2(new_n267), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n279), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(G270), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n282), .B1(new_n284), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(G200), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n602), .ZN(new_n604));
  INV_X1    g0404(.A(G303), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n528), .A2(new_n220), .B1(new_n605), .B2(new_n261), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n596), .B2(new_n597), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n604), .B1(new_n607), .B2(new_n279), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n593), .B(new_n603), .C1(new_n356), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n583), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT21), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n600), .A2(new_n602), .ZN(new_n612));
  INV_X1    g0412(.A(new_n590), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n546), .B2(new_n585), .ZN(new_n614));
  OAI21_X1  g0414(.A(G169), .B1(new_n614), .B2(new_n588), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n611), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n608), .A2(new_n592), .A3(KEYINPUT21), .A4(G169), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n612), .A2(G179), .A3(new_n592), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n581), .A2(new_n365), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n620), .B1(G179), .B2(new_n581), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n568), .B2(new_n572), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n610), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n316), .A2(new_n525), .A3(new_n554), .A4(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n583), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n568), .A2(new_n572), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n627), .B(new_n620), .C1(G179), .C2(new_n581), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n625), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n316), .A2(new_n629), .A3(new_n554), .ZN(new_n630));
  INV_X1    g0430(.A(new_n548), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n297), .A2(new_n303), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n548), .A2(new_n553), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n554), .A2(KEYINPUT26), .A3(new_n304), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n631), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n525), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n498), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n398), .A2(new_n440), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n436), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n512), .A2(new_n516), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI22_X1  g0444(.A1(new_n644), .A2(new_n363), .B1(new_n370), .B2(new_n367), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n639), .A2(new_n645), .ZN(G369));
  NAND3_X1  g0446(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n593), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n619), .B(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n655), .A2(new_n609), .ZN(new_n656));
  XOR2_X1   g0456(.A(KEYINPUT88), .B(G330), .Z(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n628), .A2(new_n652), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n627), .A2(new_n652), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n622), .B1(new_n583), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT89), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n626), .A2(new_n652), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n628), .B2(new_n652), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n665), .A2(new_n668), .ZN(G399));
  INV_X1    g0469(.A(new_n210), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G41), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n672), .A2(G1), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n213), .B2(new_n672), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  INV_X1    g0476(.A(G179), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n600), .A2(new_n677), .A3(new_n602), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n551), .A2(new_n578), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(KEYINPUT30), .A4(new_n296), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n298), .A2(new_n551), .A3(new_n299), .A4(new_n578), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n604), .B(G179), .C1(new_n607), .C2(new_n279), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n302), .B1(new_n578), .B2(new_n282), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n685), .A2(new_n608), .A3(new_n300), .A4(new_n537), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n680), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(KEYINPUT31), .B1(new_n687), .B2(new_n652), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n684), .A2(new_n686), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT90), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n684), .A2(KEYINPUT90), .A3(new_n686), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(new_n680), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n652), .A2(KEYINPUT31), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n688), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n316), .A2(new_n623), .A3(new_n554), .A4(new_n653), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n657), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n652), .B1(new_n630), .B2(new_n637), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT29), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n697), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n676), .B1(new_n702), .B2(G1), .ZN(G364));
  AND2_X1   g0503(.A1(new_n207), .A2(G13), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n206), .B1(new_n704), .B2(G45), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n671), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n659), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n656), .A2(new_n658), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(G13), .A2(G33), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(G20), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n656), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT91), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n210), .B(new_n261), .C1(new_n716), .C2(G355), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT91), .B1(new_n204), .B2(G87), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n717), .A2(new_n718), .B1(G116), .B2(new_n210), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n670), .A2(new_n261), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(G45), .B2(new_n213), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT92), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n248), .A2(G45), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n719), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n215), .B1(G20), .B2(new_n365), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n713), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g0526(.A(new_n726), .B(KEYINPUT93), .Z(new_n727));
  OAI21_X1  g0527(.A(new_n707), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n207), .A2(new_n356), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n308), .A2(G179), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G87), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n207), .A2(G190), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n730), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n733), .B(new_n261), .C1(new_n203), .C2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n302), .A2(G20), .A3(G200), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G190), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n736), .B1(G68), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G179), .A2(G200), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G159), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n207), .B1(new_n740), .B2(G190), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n743), .A2(KEYINPUT32), .B1(G97), .B2(new_n745), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n739), .B(new_n746), .C1(KEYINPUT32), .C2(new_n743), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n302), .A2(new_n308), .A3(new_n729), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n302), .A2(new_n308), .A3(new_n734), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI22_X1  g0551(.A1(G58), .A2(new_n749), .B1(new_n751), .B2(G77), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n737), .A2(new_n356), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n752), .B1(new_n218), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n267), .B1(new_n731), .B2(new_n605), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT94), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  INV_X1    g0558(.A(G329), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n735), .A2(new_n758), .B1(new_n741), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n760), .B1(G294), .B2(new_n745), .ZN(new_n761));
  INV_X1    g0561(.A(G322), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n757), .B(new_n761), .C1(new_n762), .C2(new_n748), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n753), .A2(G326), .ZN(new_n764));
  INV_X1    g0564(.A(G311), .ZN(new_n765));
  INV_X1    g0565(.A(new_n738), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT33), .B(G317), .Z(new_n767));
  OAI221_X1 g0567(.A(new_n764), .B1(new_n765), .B2(new_n750), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  OAI22_X1  g0568(.A1(new_n747), .A2(new_n755), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n769), .A2(KEYINPUT95), .ZN(new_n770));
  INV_X1    g0570(.A(new_n725), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n769), .B2(KEYINPUT95), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n728), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n708), .A2(new_n710), .B1(new_n715), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(G396));
  NOR2_X1   g0575(.A1(new_n398), .A2(new_n652), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n400), .B1(new_n380), .B2(new_n653), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(new_n777), .B2(new_n398), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n698), .B(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n697), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n707), .B1(new_n779), .B2(new_n780), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n707), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n725), .A2(new_n711), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(new_n224), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n778), .A2(new_n712), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G283), .A2(new_n738), .B1(new_n753), .B2(G303), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n585), .B2(new_n750), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT96), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n267), .B1(new_n731), .B2(new_n203), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT97), .Z(new_n793));
  NOR2_X1   g0593(.A1(new_n735), .A2(new_n449), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G311), .B2(new_n742), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n202), .B2(new_n744), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(G294), .B2(new_n749), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n791), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G137), .A2(new_n753), .B1(new_n738), .B2(G150), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT98), .ZN(new_n800));
  INV_X1    g0600(.A(G143), .ZN(new_n801));
  INV_X1    g0601(.A(G159), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n800), .B1(new_n801), .B2(new_n748), .C1(new_n802), .C2(new_n750), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT34), .Z(new_n804));
  INV_X1    g0604(.A(new_n735), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G68), .A2(new_n805), .B1(new_n742), .B2(G132), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n267), .B1(new_n732), .B2(G50), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(new_n471), .C2(new_n744), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n798), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n787), .B(new_n788), .C1(new_n725), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n783), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(G384));
  INV_X1    g0612(.A(KEYINPUT35), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n258), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n814), .A2(G20), .A3(G116), .A4(new_n216), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT99), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n815), .A2(new_n816), .B1(new_n813), .B2(new_n258), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(new_n816), .B2(new_n815), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT36), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n214), .B(G77), .C1(new_n471), .C2(new_n340), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n218), .A2(G68), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n206), .B(G13), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT37), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n650), .B1(new_n482), .B2(new_n489), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n466), .B2(new_n496), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n518), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT100), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n518), .A2(new_n826), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(KEYINPUT37), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n829), .A2(KEYINPUT100), .A3(KEYINPUT37), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n825), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n523), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT38), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n833), .B(KEYINPUT38), .C1(new_n523), .C2(new_n834), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n837), .A2(KEYINPUT39), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT101), .B1(new_n467), .B2(new_n490), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT101), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n496), .A2(new_n466), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n840), .A2(new_n842), .A3(new_n834), .ZN(new_n843));
  INV_X1    g0643(.A(new_n518), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT37), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n845), .A2(new_n827), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n834), .B1(new_n643), .B2(new_n640), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n836), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n838), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT39), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n432), .A2(new_n435), .ZN(new_n852));
  INV_X1    g0652(.A(new_n412), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(new_n652), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n839), .A2(new_n851), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n650), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n643), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n837), .A2(new_n838), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n776), .B1(new_n698), .B2(new_n778), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n412), .A2(new_n653), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n854), .A2(new_n439), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n861), .B1(new_n436), .B2(new_n440), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n858), .B1(new_n859), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n856), .A2(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n523), .B(new_n444), .C1(new_n700), .C2(new_n701), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n645), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n869), .B(new_n871), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n521), .B1(new_n519), .B2(new_n520), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n640), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n825), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT38), .B1(new_n876), .B2(new_n833), .ZN(new_n877));
  INV_X1    g0677(.A(new_n838), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT40), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n687), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(new_n688), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n696), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n865), .A2(new_n880), .A3(new_n778), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n862), .B1(new_n854), .B2(new_n439), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n436), .A2(new_n440), .A3(new_n861), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n778), .B(new_n883), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n838), .B2(new_n848), .ZN(new_n888));
  OAI22_X1  g0688(.A1(new_n879), .A2(new_n884), .B1(new_n880), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n525), .A2(new_n883), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n889), .B(new_n890), .Z(new_n891));
  OAI21_X1  g0691(.A(new_n872), .B1(new_n891), .B2(new_n657), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n206), .B2(new_n704), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n872), .A2(new_n891), .A3(new_n657), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n823), .B1(new_n893), .B2(new_n894), .ZN(G367));
  NOR2_X1   g0695(.A1(new_n550), .A2(new_n653), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n634), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n631), .A2(new_n896), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT43), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n316), .B1(new_n306), .B2(new_n653), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n304), .A2(new_n652), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n906), .A2(new_n667), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT102), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n633), .B1(new_n903), .B2(new_n628), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n908), .A2(KEYINPUT42), .B1(new_n653), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n902), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(KEYINPUT43), .B2(new_n899), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n665), .A2(new_n905), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n910), .A2(new_n901), .A3(new_n900), .A4(new_n912), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n914), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n899), .A2(KEYINPUT43), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n919), .B(new_n902), .C1(new_n910), .C2(new_n912), .ZN(new_n920));
  INV_X1    g0720(.A(new_n917), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n915), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n671), .B(KEYINPUT41), .Z(new_n923));
  NAND2_X1  g0723(.A1(new_n668), .A2(new_n906), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT44), .Z(new_n925));
  NOR2_X1   g0725(.A1(new_n668), .A2(new_n906), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT45), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n665), .ZN(new_n929));
  INV_X1    g0729(.A(new_n665), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(new_n927), .A3(new_n925), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT103), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n659), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n663), .B(new_n666), .Z(new_n934));
  XNOR2_X1  g0734(.A(new_n933), .B(new_n934), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n929), .A2(new_n702), .A3(new_n931), .A4(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n923), .B1(new_n936), .B2(new_n702), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n918), .B(new_n922), .C1(new_n937), .C2(new_n706), .ZN(new_n938));
  INV_X1    g0738(.A(new_n374), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n727), .B1(new_n670), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n720), .A2(new_n239), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n784), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n754), .A2(new_n765), .B1(new_n758), .B2(new_n750), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(G303), .B2(new_n749), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n731), .A2(new_n585), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n945), .A2(KEYINPUT46), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n945), .A2(KEYINPUT46), .B1(G107), .B2(new_n745), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n735), .A2(new_n202), .ZN(new_n948));
  INV_X1    g0748(.A(G317), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n267), .B1(new_n741), .B2(new_n949), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n948), .B(new_n950), .C1(new_n738), .C2(G294), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n944), .A2(new_n946), .A3(new_n947), .A4(new_n951), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n738), .A2(G159), .B1(new_n751), .B2(G50), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT104), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n261), .B1(new_n744), .B2(new_n340), .C1(new_n224), .C2(new_n735), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G150), .B2(new_n749), .ZN(new_n956));
  INV_X1    g0756(.A(G137), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n731), .A2(new_n471), .B1(new_n741), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT105), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n956), .B(new_n959), .C1(new_n801), .C2(new_n754), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n952), .B1(new_n954), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT47), .Z(new_n962));
  OAI221_X1 g0762(.A(new_n942), .B1(new_n714), .B2(new_n899), .C1(new_n962), .C2(new_n771), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n938), .A2(new_n963), .ZN(G387));
  NAND2_X1  g0764(.A1(new_n935), .A2(new_n706), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n935), .A2(new_n702), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n935), .A2(new_n702), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n671), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n738), .A2(new_n483), .B1(new_n751), .B2(G68), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n753), .A2(G159), .B1(new_n749), .B2(G50), .ZN(new_n970));
  XNOR2_X1  g0770(.A(KEYINPUT106), .B(G150), .ZN(new_n971));
  OAI22_X1  g0771(.A1(new_n731), .A2(new_n224), .B1(new_n741), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n744), .A2(new_n374), .ZN(new_n973));
  NOR4_X1   g0773(.A1(new_n972), .A2(new_n948), .A3(new_n973), .A4(new_n267), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n969), .A2(new_n970), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n261), .B1(new_n742), .B2(G326), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n732), .A2(G294), .B1(new_n745), .B2(G283), .ZN(new_n977));
  AOI22_X1  g0777(.A1(G303), .A2(new_n751), .B1(new_n749), .B2(G317), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n754), .B2(new_n762), .C1(new_n765), .C2(new_n766), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT107), .Z(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n977), .B1(new_n981), .B2(KEYINPUT48), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n982), .B1(KEYINPUT48), .B2(new_n981), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT108), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT49), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n976), .B1(new_n585), .B2(new_n735), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n984), .A2(new_n985), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n975), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n988), .A2(new_n725), .ZN(new_n989));
  INV_X1    g0789(.A(new_n673), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n990), .A2(new_n210), .A3(new_n261), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(G107), .B2(new_n210), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n236), .A2(G45), .ZN(new_n993));
  INV_X1    g0793(.A(new_n720), .ZN(new_n994));
  AOI211_X1 g0794(.A(G45), .B(new_n990), .C1(G68), .C2(G77), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n334), .A2(G50), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT50), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n994), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n992), .B1(new_n993), .B2(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n707), .B1(new_n727), .B2(new_n999), .C1(new_n663), .C2(new_n714), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n965), .B1(new_n966), .B2(new_n968), .C1(new_n989), .C2(new_n1000), .ZN(G393));
  INV_X1    g0801(.A(new_n929), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n931), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n967), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1004), .A2(new_n671), .A3(new_n936), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n753), .A2(G150), .B1(new_n749), .B2(G159), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT51), .Z(new_n1007));
  OAI22_X1  g0807(.A1(new_n731), .A2(new_n340), .B1(new_n741), .B2(new_n801), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n744), .A2(new_n224), .ZN(new_n1009));
  NOR4_X1   g0809(.A1(new_n1008), .A2(new_n794), .A3(new_n1009), .A4(new_n267), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n738), .A2(G50), .B1(new_n751), .B2(new_n483), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n753), .A2(G317), .B1(new_n749), .B2(G311), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT52), .Z(new_n1014));
  OAI21_X1  g0814(.A(new_n267), .B1(new_n735), .B2(new_n203), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n731), .A2(new_n758), .B1(new_n741), .B2(new_n762), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(G116), .C2(new_n745), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n738), .A2(G303), .B1(new_n751), .B2(G294), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1014), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1012), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n771), .B1(new_n1020), .B2(KEYINPUT110), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(KEYINPUT110), .B2(new_n1020), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n727), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n202), .B2(new_n210), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n994), .A2(new_n243), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n707), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT109), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1022), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n906), .B2(new_n713), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1029), .B1(new_n1030), .B2(new_n706), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1005), .A2(new_n1031), .ZN(G390));
  NAND2_X1  g0832(.A1(new_n839), .A2(new_n851), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n698), .A2(new_n778), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n776), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n855), .B1(new_n1036), .B2(new_n865), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n849), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n697), .A2(new_n778), .A3(new_n865), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n887), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1043), .A2(G330), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1037), .B1(new_n851), .B2(new_n839), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1037), .A2(new_n849), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1048), .A2(new_n705), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1033), .A2(new_n711), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n785), .ZN(new_n1051));
  INV_X1    g0851(.A(G132), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(KEYINPUT54), .B(G143), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n1052), .A2(new_n748), .B1(new_n750), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G137), .B2(new_n738), .ZN(new_n1055));
  INV_X1    g0855(.A(G125), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n261), .B1(new_n741), .B2(new_n1056), .C1(new_n218), .C2(new_n735), .ZN(new_n1057));
  OR3_X1    g0857(.A1(new_n731), .A2(new_n971), .A3(KEYINPUT53), .ZN(new_n1058));
  OAI21_X1  g0858(.A(KEYINPUT53), .B1(new_n731), .B2(new_n971), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(new_n802), .C2(new_n744), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1057), .B(new_n1060), .C1(G128), .C2(new_n753), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n766), .A2(new_n203), .B1(new_n585), .B2(new_n748), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n754), .A2(new_n758), .B1(new_n202), .B2(new_n750), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n805), .A2(G68), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n742), .A2(G294), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n733), .A2(new_n1065), .A3(new_n1066), .A4(new_n267), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1067), .A2(new_n1009), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1055), .A2(new_n1061), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n707), .B1(new_n483), .B2(new_n1051), .C1(new_n1069), .C2(new_n771), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT111), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1049), .B1(new_n1050), .B2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n883), .A2(G330), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1073), .A2(new_n778), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n860), .A2(new_n866), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n867), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1036), .A2(new_n865), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n697), .A2(new_n778), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n860), .A2(new_n866), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n444), .A2(new_n1073), .A3(new_n523), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n698), .B(KEYINPUT29), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1082), .B(new_n645), .C1(new_n1083), .C2(new_n524), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1048), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1084), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1042), .A2(new_n1047), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1087), .A2(new_n671), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1072), .A2(new_n1090), .ZN(G378));
  XOR2_X1   g0891(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT114), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n364), .A2(new_n650), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n442), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n442), .A2(new_n1096), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1094), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1099), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n1101), .A2(new_n1097), .A3(KEYINPUT114), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1093), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(KEYINPUT114), .B1(new_n1101), .B2(new_n1097), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1098), .A2(new_n1099), .A3(new_n1094), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n1105), .A3(new_n1092), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n889), .B2(G330), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n880), .B1(new_n849), .B2(new_n1043), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n884), .B1(new_n837), .B2(new_n838), .ZN(new_n1110));
  OAI211_X1 g0910(.A(G330), .B(new_n1107), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n869), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(G330), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1107), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n856), .A2(new_n868), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1117), .A3(new_n1111), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1113), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n706), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n784), .B1(new_n218), .B2(new_n785), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n731), .A2(new_n1053), .B1(new_n744), .B2(new_n336), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n753), .A2(G125), .B1(new_n749), .B2(G128), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n957), .B2(new_n750), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1122), .B(new_n1124), .C1(G132), .C2(new_n738), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT59), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n263), .B(new_n278), .C1(new_n735), .C2(new_n802), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G124), .B2(new_n742), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1127), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n766), .A2(new_n202), .B1(new_n374), .B2(new_n750), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G116), .B2(new_n753), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n748), .A2(new_n203), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT112), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n735), .A2(new_n471), .B1(new_n741), .B2(new_n758), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n278), .B(new_n267), .C1(new_n731), .C2(new_n224), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1136), .B(new_n1137), .C1(G68), .C2(new_n745), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1133), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT113), .B(KEYINPUT58), .ZN(new_n1140));
  OR2_X1    g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1142));
  AOI21_X1  g0942(.A(G50), .B1(new_n263), .B2(new_n278), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n261), .B2(G41), .ZN(new_n1144));
  AND4_X1   g0944(.A1(new_n1131), .A2(new_n1141), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n1121), .B1(new_n771), .B2(new_n1145), .C1(new_n1107), .C2(new_n712), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1120), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1089), .A2(new_n1085), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1119), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n671), .B1(new_n1149), .B2(KEYINPUT57), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1148), .A2(KEYINPUT57), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT115), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1113), .A2(new_n1152), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1116), .A2(new_n1117), .A3(new_n1111), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1116), .A2(new_n1111), .B1(new_n856), .B2(new_n868), .ZN(new_n1155));
  OAI21_X1  g0955(.A(KEYINPUT115), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1151), .B1(new_n1153), .B2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1147), .B1(new_n1150), .B2(new_n1157), .ZN(G375));
  NAND2_X1  g0958(.A1(new_n1081), .A2(new_n706), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n784), .B1(new_n340), .B2(new_n785), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n731), .A2(new_n202), .B1(new_n741), .B2(new_n605), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n261), .B1(new_n805), .B2(G77), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT116), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n973), .B(new_n1161), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n1163), .B2(new_n1162), .C1(new_n203), .C2(new_n750), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n753), .A2(G294), .B1(new_n749), .B2(G283), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n585), .B2(new_n766), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1168), .A2(KEYINPUT117), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(KEYINPUT117), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n744), .A2(new_n218), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n754), .A2(new_n1052), .B1(new_n957), .B2(new_n748), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n766), .A2(new_n1053), .B1(new_n336), .B2(new_n750), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G159), .A2(new_n732), .B1(new_n742), .B2(G128), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1174), .B(new_n261), .C1(new_n471), .C2(new_n735), .ZN(new_n1175));
  OR4_X1    g0975(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .A4(new_n1175), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1169), .A2(new_n1170), .A3(new_n1176), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1160), .B1(new_n771), .B2(new_n1177), .C1(new_n865), .C2(new_n712), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1159), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n923), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1076), .A2(new_n1084), .A3(new_n1080), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1086), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1183), .ZN(G381));
  OR4_X1    g0984(.A1(G396), .A2(G390), .A3(G393), .A4(G384), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1185), .A2(G387), .A3(G381), .ZN(new_n1186));
  INV_X1    g0986(.A(G378), .ZN(new_n1187));
  INV_X1    g0987(.A(G375), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(G407));
  NAND2_X1  g0989(.A1(new_n651), .A2(G213), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n1187), .A3(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(G407), .A2(G213), .A3(new_n1192), .ZN(G409));
  XNOR2_X1  g0993(.A(G393), .B(new_n774), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n938), .A2(new_n963), .A3(G390), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G390), .B1(new_n938), .B2(new_n963), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1195), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1198), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT61), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1152), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1155), .A2(KEYINPUT115), .ZN(new_n1205));
  OAI21_X1  g1005(.A(KEYINPUT119), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT119), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1156), .A2(new_n1207), .A3(new_n1153), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1206), .A2(new_n1208), .A3(new_n706), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1119), .A2(new_n1148), .A3(new_n1181), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT118), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1119), .A2(new_n1148), .A3(KEYINPUT118), .A4(new_n1181), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n1146), .A3(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1187), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(G378), .B(new_n1147), .C1(new_n1150), .C2(new_n1157), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1191), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT120), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT60), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1182), .B1(new_n1088), .B2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1076), .A2(new_n1084), .A3(new_n1080), .A4(KEYINPUT60), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1221), .A2(new_n671), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n811), .B(new_n1179), .C1(new_n1220), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1220), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G384), .B1(new_n1225), .B2(new_n1180), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1218), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1086), .A2(KEYINPUT60), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1222), .B1(new_n1228), .B2(new_n1182), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n811), .B1(new_n1229), .B2(new_n1179), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1225), .A2(G384), .A3(new_n1180), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(KEYINPUT120), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1191), .A2(G2897), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1227), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT121), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1233), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1227), .A2(new_n1232), .A3(new_n1235), .A4(new_n1233), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1203), .B1(new_n1217), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT123), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT123), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n1203), .C1(new_n1217), .C2(new_n1241), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1227), .A2(new_n1232), .ZN(new_n1248));
  OR2_X1    g1048(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1247), .A2(new_n1190), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1249), .B1(new_n1217), .B2(new_n1248), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1202), .B1(new_n1246), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT122), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1241), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1217), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1241), .A2(new_n1256), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1217), .A2(KEYINPUT63), .A3(new_n1248), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT63), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1248), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1258), .B2(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1202), .A2(KEYINPUT61), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1260), .A2(new_n1261), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1255), .A2(new_n1266), .ZN(G405));
  XNOR2_X1  g1067(.A(G375), .B(G378), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1236), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1188), .A2(G378), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1216), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1248), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1272), .A3(KEYINPUT125), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT125), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1268), .A2(new_n1274), .A3(new_n1236), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1202), .A2(KEYINPUT126), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1273), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1199), .A2(new_n1201), .A3(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(KEYINPUT127), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT127), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1279), .B(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1283), .A2(new_n1273), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(G402));
endmodule


