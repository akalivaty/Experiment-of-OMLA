//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n812, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT14), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT14), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n209), .A2(KEYINPUT88), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n209), .B2(KEYINPUT88), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n204), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT89), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n202), .A2(new_n203), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n204), .A2(new_n209), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n213), .A2(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT17), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(G1gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(G1gat), .B2(new_n221), .ZN(new_n224));
  XOR2_X1   g023(.A(new_n224), .B(G8gat), .Z(new_n225));
  NAND2_X1  g024(.A1(new_n215), .A2(new_n218), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT17), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n220), .A2(new_n225), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n225), .A2(KEYINPUT90), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n225), .A2(KEYINPUT90), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(new_n226), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT18), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n232), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n219), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(new_n233), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n230), .B(KEYINPUT13), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n229), .A2(KEYINPUT18), .A3(new_n230), .A4(new_n233), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G197gat), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT11), .B(G169gat), .Z(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g046(.A(new_n247), .B(KEYINPUT12), .Z(new_n248));
  NAND2_X1  g047(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n248), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n236), .A2(new_n241), .A3(new_n250), .A4(new_n242), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G78gat), .B(G106gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT31), .B(G50gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G228gat), .A2(G233gat), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n258), .B(KEYINPUT81), .Z(new_n259));
  NAND2_X1  g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260));
  INV_X1    g059(.A(G155gat), .ZN(new_n261));
  INV_X1    g060(.A(G162gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n260), .B1(new_n263), .B2(KEYINPUT2), .ZN(new_n264));
  INV_X1    g063(.A(G141gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G148gat), .ZN(new_n266));
  INV_X1    g065(.A(G148gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G141gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT74), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n265), .A2(KEYINPUT74), .A3(G148gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n264), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G141gat), .B(G148gat), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n260), .B(new_n263), .C1(new_n273), .C2(KEYINPUT2), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT29), .ZN(new_n276));
  XNOR2_X1  g075(.A(G211gat), .B(G218gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(G197gat), .B(G204gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(G211gat), .A2(G218gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT22), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n277), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n277), .B1(new_n281), .B2(new_n278), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n276), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n275), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n278), .A2(new_n281), .ZN(new_n288));
  INV_X1    g087(.A(new_n277), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n282), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n272), .A2(new_n274), .A3(new_n286), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(new_n276), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n259), .B1(new_n287), .B2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT82), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT3), .B1(new_n285), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT29), .B1(new_n290), .B2(new_n282), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT82), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n275), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n293), .ZN(new_n300));
  INV_X1    g099(.A(new_n258), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n294), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G22gat), .ZN(new_n304));
  INV_X1    g103(.A(G22gat), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n294), .B(new_n305), .C1(new_n299), .C2(new_n302), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n257), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n256), .B1(new_n303), .B2(G22gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n272), .A2(new_n274), .ZN(new_n309));
  INV_X1    g108(.A(new_n298), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n286), .B1(new_n297), .B2(KEYINPUT82), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n312), .A2(new_n300), .A3(new_n301), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT83), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n313), .A2(new_n314), .A3(new_n305), .A4(new_n294), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n306), .A2(KEYINPUT83), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n308), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT84), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n308), .A2(new_n316), .A3(new_n315), .A4(KEYINPUT84), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n307), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(KEYINPUT24), .ZN(new_n326));
  INV_X1    g125(.A(G183gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G190gat), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(G183gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n326), .B1(new_n331), .B2(KEYINPUT24), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT25), .ZN(new_n333));
  INV_X1    g132(.A(G169gat), .ZN(new_n334));
  INV_X1    g133(.A(G176gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n333), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n337), .A2(G169gat), .A3(G176gat), .ZN(new_n339));
  AND2_X1   g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT64), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT23), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT64), .ZN(new_n344));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n332), .A2(new_n338), .A3(new_n341), .A4(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT24), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(G183gat), .A3(G190gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(G183gat), .B(G190gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n348), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n337), .B1(G169gat), .B2(G176gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n343), .A2(new_n352), .A3(new_n345), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n333), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT72), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT26), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n336), .A2(new_n357), .A3(new_n345), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n342), .A2(KEYINPUT26), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n325), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n361), .A2(KEYINPUT65), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT27), .B(G183gat), .ZN(new_n363));
  AOI21_X1  g162(.A(G190gat), .B1(new_n361), .B2(KEYINPUT65), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n362), .A3(new_n364), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n355), .A2(new_n356), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n356), .B1(new_n355), .B2(new_n368), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n324), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT71), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT29), .B1(new_n355), .B2(new_n368), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(new_n324), .ZN(new_n374));
  INV_X1    g173(.A(new_n367), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n375), .A2(new_n360), .A3(new_n365), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(new_n354), .B2(new_n347), .ZN(new_n377));
  OAI211_X1 g176(.A(KEYINPUT71), .B(new_n323), .C1(new_n377), .C2(KEYINPUT29), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n371), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT73), .ZN(new_n380));
  INV_X1    g179(.A(new_n291), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n323), .A2(new_n276), .ZN(new_n383));
  INV_X1    g182(.A(new_n369), .ZN(new_n384));
  INV_X1    g183(.A(new_n370), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n329), .A2(G183gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n327), .A2(G190gat), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT24), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n389), .A2(new_n349), .A3(new_n338), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n339), .A2(KEYINPUT64), .A3(new_n340), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n344), .B1(new_n343), .B2(new_n345), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n340), .B1(KEYINPUT23), .B2(new_n342), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n389), .A2(new_n349), .A3(new_n394), .A4(new_n352), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n390), .A2(new_n393), .B1(new_n395), .B2(new_n333), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n396), .A2(new_n323), .A3(new_n376), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n291), .B1(new_n386), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n380), .B1(new_n379), .B2(new_n381), .ZN(new_n400));
  XNOR2_X1  g199(.A(G8gat), .B(G36gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n401), .B(new_n402), .Z(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n399), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT30), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n404), .B1(new_n399), .B2(new_n400), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n379), .A2(new_n381), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT73), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n409), .A2(new_n398), .A3(new_n382), .A4(new_n403), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n407), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT39), .ZN(new_n414));
  INV_X1    g213(.A(G120gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G113gat), .ZN(new_n416));
  INV_X1    g215(.A(G113gat), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(G120gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n418), .A3(KEYINPUT66), .ZN(new_n419));
  OR3_X1    g218(.A1(new_n415), .A2(KEYINPUT66), .A3(G113gat), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT1), .ZN(new_n421));
  XNOR2_X1  g220(.A(G127gat), .B(G134gat), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(G127gat), .B(G134gat), .Z(new_n424));
  XNOR2_X1  g223(.A(G113gat), .B(G120gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n424), .B1(KEYINPUT1), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n427), .A2(new_n309), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n426), .A2(new_n423), .B1(new_n272), .B2(new_n274), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(G225gat), .A2(G233gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n431), .B(KEYINPUT75), .Z(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n414), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n309), .A2(KEYINPUT3), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(new_n427), .A3(new_n292), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n423), .A2(new_n426), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(new_n275), .A3(KEYINPUT4), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n439), .B1(new_n427), .B2(new_n309), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n438), .A2(KEYINPUT79), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT79), .B1(new_n438), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n436), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n434), .B1(new_n444), .B2(new_n433), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n414), .A3(new_n432), .ZN(new_n446));
  XNOR2_X1  g245(.A(G57gat), .B(G85gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT78), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G1gat), .B(G29gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n450), .B(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n446), .A2(KEYINPUT85), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT85), .B1(new_n446), .B2(new_n452), .ZN(new_n454));
  OAI211_X1 g253(.A(KEYINPUT40), .B(new_n445), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT76), .B1(new_n430), .B2(new_n433), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n436), .A2(new_n440), .A3(new_n438), .A4(new_n433), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT76), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n458), .B(new_n432), .C1(new_n428), .C2(new_n429), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT5), .A4(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT5), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n436), .A2(new_n461), .A3(new_n433), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(new_n441), .B2(new_n442), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n452), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n445), .B1(new_n453), .B2(new_n454), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT40), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n413), .A2(new_n455), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT37), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n409), .A2(new_n469), .A3(new_n398), .A4(new_n382), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT86), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n382), .A2(new_n398), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT86), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n469), .A4(new_n409), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n386), .A2(new_n397), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n469), .B1(new_n476), .B2(new_n381), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n379), .A2(new_n291), .ZN(new_n478));
  AOI211_X1 g277(.A(KEYINPUT38), .B(new_n403), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n460), .A2(new_n463), .ZN(new_n481));
  INV_X1    g280(.A(new_n452), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT6), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n460), .A2(new_n452), .A3(new_n463), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n464), .A2(KEYINPUT6), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT87), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n487), .A2(KEYINPUT87), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n488), .A2(new_n405), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n480), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT38), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n472), .A2(new_n409), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n403), .B1(new_n493), .B2(KEYINPUT37), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n475), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n322), .B(new_n468), .C1(new_n491), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n486), .A2(new_n487), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n497), .B1(new_n405), .B2(KEYINPUT30), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n407), .B1(new_n410), .B2(new_n411), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT80), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n410), .A2(new_n411), .B1(new_n486), .B2(new_n487), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT80), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n501), .A2(new_n406), .A3(new_n502), .A4(new_n407), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(new_n321), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n437), .B1(new_n396), .B2(new_n376), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n355), .A2(new_n368), .A3(new_n427), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(G227gat), .A2(G233gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT34), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n511), .B1(new_n509), .B2(KEYINPUT70), .ZN(new_n512));
  XOR2_X1   g311(.A(new_n510), .B(new_n512), .Z(new_n513));
  XNOR2_X1  g312(.A(G15gat), .B(G43gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT69), .ZN(new_n515));
  XOR2_X1   g314(.A(G71gat), .B(G99gat), .Z(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n509), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n506), .A2(new_n518), .A3(new_n507), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT67), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT67), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n506), .A2(new_n521), .A3(new_n518), .A4(new_n507), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n517), .B1(new_n523), .B2(KEYINPUT32), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT33), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT68), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT68), .ZN(new_n527));
  AOI211_X1 g326(.A(new_n527), .B(KEYINPUT33), .C1(new_n520), .C2(new_n522), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n524), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n523), .B(KEYINPUT32), .C1(new_n525), .C2(new_n517), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n513), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n513), .A3(new_n530), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(KEYINPUT36), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n529), .A2(new_n513), .A3(new_n530), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(new_n531), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n496), .A2(new_n505), .A3(new_n538), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n536), .A2(new_n531), .A3(new_n321), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n500), .A3(new_n503), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n488), .A2(new_n489), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n413), .A2(new_n543), .A3(KEYINPUT35), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n540), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n253), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT92), .B(G57gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G64gat), .ZN(new_n549));
  INV_X1    g348(.A(G64gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G57gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552));
  NAND2_X1  g351(.A1(G71gat), .A2(G78gat), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n549), .A2(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G71gat), .B(G78gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT93), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(G71gat), .A2(G78gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n553), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n559), .B2(new_n558), .ZN(new_n561));
  INV_X1    g360(.A(new_n551), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n550), .A2(G57gat), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT9), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT21), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G127gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n237), .B1(new_n567), .B2(new_n566), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(G155gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n574), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT94), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(KEYINPUT94), .A2(G85gat), .A3(G92gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(KEYINPUT7), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT7), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n583), .B(new_n589), .C1(new_n584), .C2(new_n585), .ZN(new_n590));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  AOI22_X1  g390(.A1(KEYINPUT8), .A2(new_n591), .B1(new_n584), .B2(new_n585), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  OR2_X1    g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n591), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n588), .A2(new_n596), .A3(new_n590), .A4(new_n592), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n566), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n566), .A2(new_n598), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n598), .B(KEYINPUT95), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT10), .ZN(new_n606));
  NOR3_X1   g405(.A1(new_n605), .A2(new_n606), .A3(new_n566), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n606), .A3(new_n600), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT96), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(KEYINPUT96), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n602), .B(KEYINPUT97), .Z(new_n612));
  OAI21_X1  g411(.A(new_n604), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n604), .B(new_n616), .C1(new_n611), .C2(new_n603), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n605), .ZN(new_n621));
  AND2_X1   g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  AOI22_X1  g421(.A1(new_n621), .A2(new_n226), .B1(KEYINPUT41), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n220), .A2(new_n228), .A3(new_n605), .ZN(new_n624));
  XOR2_X1   g423(.A(G190gat), .B(G218gat), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(new_n624), .B2(new_n623), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OR3_X1    g431(.A1(new_n627), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n632), .B1(new_n627), .B2(new_n628), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n582), .A2(new_n620), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n547), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n497), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n413), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n643), .A2(G8gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT16), .B(G8gat), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT42), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(KEYINPUT42), .B2(new_n646), .ZN(G1325gat));
  AND3_X1   g447(.A1(new_n534), .A2(KEYINPUT98), .A3(new_n537), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT98), .B1(new_n534), .B2(new_n537), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(G15gat), .B1(new_n638), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n536), .A2(new_n531), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(G15gat), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n652), .B1(new_n638), .B2(new_n655), .ZN(G1326gat));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n321), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT99), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT43), .B(G22gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(G1327gat));
  INV_X1    g459(.A(new_n620), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n547), .A2(new_n661), .A3(new_n582), .A4(new_n636), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n662), .A2(G29gat), .A3(new_n497), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT45), .Z(new_n664));
  NAND2_X1  g463(.A1(new_n582), .A2(new_n661), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n253), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT100), .Z(new_n667));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n541), .A2(KEYINPUT35), .B1(new_n544), .B2(new_n540), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n475), .A2(new_n494), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n480), .B(new_n490), .C1(new_n670), .C2(new_n492), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n467), .A2(new_n455), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n321), .B1(new_n672), .B2(new_n413), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n671), .A2(new_n673), .B1(new_n504), .B2(new_n321), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n669), .B1(new_n674), .B2(new_n651), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n668), .B1(new_n675), .B2(new_n635), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n539), .A2(new_n546), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n635), .A2(new_n668), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n667), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G29gat), .B1(new_n680), .B2(new_n497), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n664), .A2(new_n681), .ZN(G1328gat));
  INV_X1    g481(.A(new_n413), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n662), .A2(G36gat), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT46), .ZN(new_n685));
  OAI21_X1  g484(.A(G36gat), .B1(new_n680), .B2(new_n683), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(G1329gat));
  OAI21_X1  g486(.A(G43gat), .B1(new_n680), .B2(new_n651), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n654), .A2(G43gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n662), .B2(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT47), .Z(G1330gat));
  NAND2_X1  g490(.A1(new_n321), .A2(G50gat), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n662), .A2(new_n322), .ZN(new_n693));
  OAI22_X1  g492(.A1(new_n680), .A2(new_n692), .B1(new_n693), .B2(G50gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g494(.A1(new_n582), .A2(new_n636), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n253), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n661), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT101), .Z(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n675), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n640), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(new_n548), .Z(G1332gat));
  AOI21_X1  g501(.A(new_n683), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n704), .B(KEYINPUT102), .Z(new_n705));
  NOR2_X1   g504(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1333gat));
  INV_X1    g506(.A(G71gat), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n700), .A2(new_n708), .A3(new_n653), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n699), .A2(new_n651), .A3(new_n675), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n709), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g511(.A1(new_n700), .A2(new_n321), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G78gat), .ZN(G1335gat));
  OR3_X1    g513(.A1(new_n581), .A2(KEYINPUT103), .A3(new_n252), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT103), .B1(new_n581), .B2(new_n252), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n661), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT98), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n538), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n534), .A2(new_n537), .A3(KEYINPUT98), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n496), .A2(new_n719), .A3(new_n505), .A4(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n635), .B1(new_n721), .B2(new_n546), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n679), .B(new_n717), .C1(new_n722), .C2(KEYINPUT44), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n676), .A2(KEYINPUT104), .A3(new_n679), .A4(new_n717), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G85gat), .B1(new_n727), .B2(new_n497), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n715), .A2(new_n716), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n722), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n722), .A2(KEYINPUT51), .A3(new_n729), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n661), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(new_n584), .A3(new_n640), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n728), .A2(new_n735), .ZN(G1336gat));
  NOR2_X1   g535(.A1(new_n683), .A2(G92gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n723), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n741), .A2(KEYINPUT105), .A3(new_n413), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT105), .B1(new_n741), .B2(new_n413), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n585), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n740), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(G92gat), .B1(new_n727), .B2(new_n683), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n739), .B1(new_n746), .B2(new_n738), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n748));
  OR3_X1    g547(.A1(new_n745), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n745), .B2(new_n747), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(G1337gat));
  OAI21_X1  g550(.A(G99gat), .B1(new_n727), .B2(new_n651), .ZN(new_n752));
  INV_X1    g551(.A(G99gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n734), .A2(new_n753), .A3(new_n653), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1338gat));
  NOR2_X1   g554(.A1(new_n322), .A2(G106gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n734), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758));
  OAI21_X1  g557(.A(G106gat), .B1(new_n723), .B2(new_n322), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n725), .A2(new_n321), .A3(new_n726), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G106gat), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n763), .A2(KEYINPUT107), .B1(new_n734), .B2(new_n756), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n762), .A2(new_n765), .A3(G106gat), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n761), .B(new_n758), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(KEYINPUT107), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n766), .A3(new_n757), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT108), .B1(new_n769), .B2(KEYINPUT53), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n760), .B1(new_n767), .B2(new_n770), .ZN(G1339gat));
  INV_X1    g570(.A(new_n612), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n609), .A2(new_n610), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n772), .B(new_n773), .C1(new_n774), .C2(new_n607), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n611), .A2(new_n612), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT54), .B1(new_n611), .B2(new_n603), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n775), .B(new_n617), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n611), .A2(new_n612), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n616), .B1(new_n782), .B2(new_n773), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n776), .B(KEYINPUT54), .C1(new_n603), .C2(new_n611), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n784), .A3(KEYINPUT55), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n781), .A2(new_n252), .A3(new_n619), .A4(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n239), .A2(new_n240), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n230), .B1(new_n229), .B2(new_n233), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n247), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n620), .A2(new_n251), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n636), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n619), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT55), .B1(new_n783), .B2(new_n784), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n789), .A2(new_n251), .ZN(new_n794));
  NOR4_X1   g593(.A1(new_n792), .A2(new_n793), .A3(new_n635), .A4(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n582), .B1(new_n791), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n696), .A2(new_n253), .A3(new_n661), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n796), .A2(KEYINPUT110), .A3(new_n797), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n540), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n413), .A2(new_n497), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n253), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(new_n417), .ZN(G1340gat));
  NOR2_X1   g607(.A1(new_n806), .A2(new_n661), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n810), .B2(new_n415), .ZN(new_n811));
  XOR2_X1   g610(.A(KEYINPUT111), .B(G120gat), .Z(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n809), .B2(new_n812), .ZN(G1341gat));
  NOR2_X1   g612(.A1(new_n806), .A2(new_n582), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(new_n571), .ZN(G1342gat));
  NOR4_X1   g614(.A1(new_n413), .A2(new_n635), .A3(G134gat), .A4(new_n497), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n804), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g616(.A(new_n817), .B(KEYINPUT112), .Z(new_n818));
  OR2_X1    g617(.A1(new_n818), .A2(KEYINPUT56), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(KEYINPUT56), .ZN(new_n820));
  OAI21_X1  g619(.A(G134gat), .B1(new_n806), .B2(new_n635), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(G1343gat));
  OR3_X1    g621(.A1(new_n802), .A2(KEYINPUT116), .A3(new_n497), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT116), .B1(new_n802), .B2(new_n497), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n649), .A2(new_n650), .A3(new_n322), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n413), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n253), .A2(G141gat), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT58), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n785), .A2(new_n252), .A3(new_n619), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT113), .ZN(new_n832));
  AOI211_X1 g631(.A(new_n832), .B(KEYINPUT55), .C1(new_n783), .C2(new_n784), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT113), .B1(new_n779), .B2(new_n780), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n790), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n830), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n781), .A2(new_n832), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n793), .A2(KEYINPUT113), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g639(.A(KEYINPUT114), .B(new_n790), .C1(new_n840), .C2(new_n831), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n837), .A2(new_n635), .A3(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n795), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n581), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n797), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n321), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT57), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n800), .A2(new_n848), .A3(new_n321), .A4(new_n801), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n651), .A2(new_n805), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n847), .A2(new_n849), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT117), .B1(new_n852), .B2(new_n253), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n850), .B1(new_n846), .B2(KEYINPUT57), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n854), .A2(new_n855), .A3(new_n252), .A4(new_n849), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n853), .A2(G141gat), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n829), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n828), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n826), .A2(new_n413), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n852), .A2(KEYINPUT115), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n854), .A2(new_n862), .A3(new_n849), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n252), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n860), .B1(new_n864), .B2(G141gat), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n858), .B1(new_n865), .B2(new_n866), .ZN(G1344gat));
  NAND3_X1  g666(.A1(new_n827), .A2(new_n267), .A3(new_n620), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(G148gat), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n854), .A2(new_n862), .A3(new_n849), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n862), .B1(new_n854), .B2(new_n849), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n870), .B1(new_n873), .B2(new_n620), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT118), .B1(new_n844), .B2(new_n845), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n790), .B1(new_n840), .B2(new_n831), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n636), .B1(new_n877), .B2(new_n830), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n795), .B1(new_n878), .B2(new_n841), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n876), .B(new_n797), .C1(new_n879), .C2(new_n581), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n322), .A2(KEYINPUT57), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n875), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT57), .B1(new_n802), .B2(new_n322), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n850), .A2(new_n661), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n882), .A2(new_n883), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n886), .A2(G148gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT119), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n869), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n868), .B1(new_n874), .B2(new_n890), .ZN(G1345gat));
  NAND2_X1  g690(.A1(new_n861), .A2(new_n863), .ZN(new_n892));
  OAI21_X1  g691(.A(G155gat), .B1(new_n892), .B2(new_n582), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n827), .A2(new_n261), .A3(new_n581), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1346gat));
  OAI21_X1  g694(.A(G162gat), .B1(new_n892), .B2(new_n635), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n683), .A2(new_n262), .A3(new_n636), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n826), .B2(new_n897), .ZN(G1347gat));
  INV_X1    g697(.A(KEYINPUT121), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n800), .A2(new_n497), .A3(new_n801), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n800), .A2(KEYINPUT120), .A3(new_n497), .A4(new_n801), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n803), .A2(new_n683), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n899), .A3(new_n905), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n907), .A2(new_n334), .A3(new_n252), .A4(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT122), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n683), .A2(new_n640), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n804), .A2(new_n252), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n910), .B1(new_n912), .B2(G169gat), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n910), .A3(G169gat), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n909), .B(KEYINPUT123), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n915), .A2(new_n913), .ZN(new_n918));
  INV_X1    g717(.A(new_n905), .ZN(new_n919));
  AOI211_X1 g718(.A(KEYINPUT121), .B(new_n919), .C1(new_n902), .C2(new_n903), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n252), .A2(new_n334), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n906), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n917), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n916), .A2(new_n923), .ZN(G1348gat));
  AND2_X1   g723(.A1(new_n804), .A2(new_n911), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n925), .A2(G176gat), .A3(new_n620), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n906), .A2(new_n920), .A3(new_n661), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(G176gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n907), .A2(new_n620), .A3(new_n908), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(KEYINPUT124), .A3(new_n335), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n926), .B1(new_n929), .B2(new_n931), .ZN(G1349gat));
  AND4_X1   g731(.A1(new_n363), .A2(new_n904), .A3(new_n581), .A4(new_n905), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n327), .B1(new_n925), .B2(new_n581), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n935), .B(new_n936), .ZN(G1350gat));
  NAND4_X1  g736(.A1(new_n907), .A2(new_n329), .A3(new_n636), .A4(new_n908), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n329), .B1(new_n925), .B2(new_n636), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n939), .A2(new_n940), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n938), .B1(new_n942), .B2(new_n943), .ZN(G1351gat));
  AND2_X1   g743(.A1(new_n882), .A2(new_n884), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n651), .A2(new_n911), .ZN(new_n946));
  XOR2_X1   g745(.A(new_n946), .B(KEYINPUT126), .Z(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(G197gat), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n948), .A2(new_n949), .A3(new_n253), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n825), .A2(new_n413), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT125), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n904), .A2(new_n252), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n950), .B1(new_n949), .B2(new_n953), .ZN(G1352gat));
  NAND2_X1  g753(.A1(new_n904), .A2(new_n952), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n955), .A2(G204gat), .A3(new_n661), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n948), .B2(new_n661), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n956), .A2(new_n957), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(G1353gat));
  OR3_X1    g760(.A1(new_n955), .A2(G211gat), .A3(new_n582), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n945), .A2(new_n581), .A3(new_n947), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n963), .B2(G211gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1354gat));
  OAI21_X1  g765(.A(G218gat), .B1(new_n948), .B2(new_n635), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n635), .A2(G218gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n955), .B2(new_n968), .ZN(G1355gat));
endmodule


