//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n567, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166,
    new_n1167, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT67), .B(G96), .Z(G221));
  XOR2_X1   g012(.A(KEYINPUT68), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT69), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G567), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n451), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(G2106), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT71), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT71), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G137), .A4(new_n459), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n463), .A2(new_n466), .B1(G101), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT70), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n460), .B2(new_n461), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n470), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  AOI211_X1 g049(.A(KEYINPUT70), .B(new_n459), .C1(new_n471), .C2(new_n472), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n469), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n460), .A2(new_n461), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n459), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT73), .ZN(new_n481));
  OR2_X1    g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT72), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT72), .B1(new_n478), .B2(G2105), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G136), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n459), .A2(G112), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n481), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT74), .ZN(G162));
  INV_X1    g068(.A(KEYINPUT75), .ZN(new_n494));
  NAND2_X1  g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n482), .B2(new_n483), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n459), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n494), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n501), .A2(new_n504), .A3(KEYINPUT75), .ZN(new_n505));
  OAI211_X1 g080(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n464), .A2(new_n508), .A3(G138), .A4(new_n459), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n500), .A2(new_n505), .B1(new_n507), .B2(new_n509), .ZN(G164));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT76), .ZN(new_n512));
  AND3_X1   g087(.A1(new_n512), .A2(KEYINPUT6), .A3(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(KEYINPUT6), .B1(new_n512), .B2(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT77), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(KEYINPUT77), .A2(KEYINPUT5), .A3(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n511), .A2(new_n516), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n522), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G651), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G166));
  AND2_X1   g104(.A1(new_n520), .A2(new_n521), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n513), .A2(new_n514), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n531), .A2(new_n519), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  AND2_X1   g110(.A1(G63), .A2(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n522), .A2(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n533), .A2(new_n535), .A3(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  INV_X1    g117(.A(G52), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n543), .A2(new_n516), .B1(new_n523), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT79), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n534), .A2(G52), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT79), .ZN(new_n548));
  OAI211_X1 g123(.A(new_n547), .B(new_n548), .C1(new_n544), .C2(new_n523), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n530), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n527), .B1(new_n553), .B2(KEYINPUT78), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n554), .B1(KEYINPUT78), .B2(new_n553), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n550), .A2(new_n555), .ZN(G171));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n530), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(KEYINPUT80), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT80), .ZN(new_n561));
  OAI211_X1 g136(.A(new_n561), .B(new_n557), .C1(new_n530), .C2(new_n558), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(G651), .A3(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n532), .A2(G81), .B1(new_n534), .B2(G43), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(G860), .A3(new_n564), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT81), .Z(G188));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n530), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(new_n532), .B2(G91), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT82), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n516), .C2(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n577), .B1(KEYINPUT82), .B2(KEYINPUT9), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n534), .B(new_n579), .C1(KEYINPUT82), .C2(KEYINPUT9), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n574), .A2(new_n578), .A3(new_n580), .ZN(G299));
  NAND2_X1  g156(.A1(new_n550), .A2(new_n555), .ZN(G301));
  INV_X1    g157(.A(G166), .ZN(G303));
  NAND2_X1  g158(.A1(new_n532), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n522), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n534), .A2(G49), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(new_n534), .A2(G48), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n520), .B2(new_n521), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT83), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n515), .A2(G86), .A3(new_n522), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n588), .A2(new_n593), .A3(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n522), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n527), .ZN(new_n597));
  INV_X1    g172(.A(G47), .ZN(new_n598));
  INV_X1    g173(.A(G85), .ZN(new_n599));
  OAI221_X1 g174(.A(new_n597), .B1(new_n598), .B2(new_n516), .C1(new_n599), .C2(new_n523), .ZN(G290));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n523), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n532), .A2(KEYINPUT10), .A3(G92), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n530), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(new_n534), .B2(G54), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT84), .B1(new_n611), .B2(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  MUX2_X1   g188(.A(KEYINPUT84), .B(new_n612), .S(new_n613), .Z(G284));
  MUX2_X1   g189(.A(KEYINPUT84), .B(new_n612), .S(new_n613), .Z(G321));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(G299), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n616), .B2(G168), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(new_n616), .B2(G168), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n611), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n563), .A2(new_n564), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n611), .A2(new_n620), .ZN(new_n623));
  MUX2_X1   g198(.A(new_n622), .B(new_n623), .S(G868), .Z(G323));
  XOR2_X1   g199(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n625));
  XNOR2_X1  g200(.A(G323), .B(new_n625), .ZN(G282));
  NAND2_X1  g201(.A1(new_n464), .A2(new_n468), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT13), .Z(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(G2100), .ZN(new_n631));
  OAI21_X1  g206(.A(KEYINPUT87), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G111), .B2(new_n459), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n459), .A2(G111), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n467), .B1(new_n634), .B2(KEYINPUT87), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n479), .A2(G123), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n486), .A2(new_n487), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n630), .A2(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(G2096), .ZN(new_n642));
  NAND4_X1  g217(.A1(new_n631), .A2(new_n640), .A3(new_n641), .A4(new_n642), .ZN(G156));
  XOR2_X1   g218(.A(G2443), .B(G2446), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT89), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2451), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT92), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n646), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT14), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT91), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2427), .B(G2430), .Z(new_n654));
  AOI21_X1  g229(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n655), .B1(new_n654), .B2(new_n653), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n649), .B(new_n656), .Z(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT88), .B(KEYINPUT16), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT90), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2454), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(G14), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n657), .A2(new_n660), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(G401));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT17), .Z(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  INV_X1    g245(.A(new_n667), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(new_n665), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n669), .B(new_n670), .C1(new_n668), .C2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n665), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT18), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2096), .B(G2100), .Z(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G227));
  XOR2_X1   g256(.A(G1971), .B(G1976), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1956), .B(G2474), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(new_n686), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT20), .Z(new_n690));
  AOI211_X1 g265(.A(new_n688), .B(new_n690), .C1(new_n683), .C2(new_n687), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1991), .B(G1996), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  XNOR2_X1  g272(.A(KEYINPUT97), .B(G16), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n699), .A2(G22), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(G1971), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(G23), .B(G288), .S(G16), .Z(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  MUX2_X1   g281(.A(G6), .B(G305), .S(G16), .Z(new_n707));
  XOR2_X1   g282(.A(KEYINPUT32), .B(G1981), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n703), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n710), .A2(KEYINPUT34), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G25), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n479), .A2(G119), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n459), .A2(G107), .ZN(new_n715));
  OAI21_X1  g290(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n716));
  INV_X1    g291(.A(G131), .ZN(new_n717));
  OAI221_X1 g292(.A(new_n714), .B1(new_n715), .B2(new_n716), .C1(new_n637), .C2(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT95), .Z(new_n719));
  OAI21_X1  g294(.A(new_n713), .B1(new_n719), .B2(new_n712), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT35), .B(G1991), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT96), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n720), .B(new_n722), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n710), .A2(KEYINPUT34), .ZN(new_n724));
  MUX2_X1   g299(.A(G24), .B(G290), .S(new_n699), .Z(new_n725));
  XOR2_X1   g300(.A(KEYINPUT98), .B(G1986), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n711), .A2(new_n723), .A3(new_n724), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(KEYINPUT99), .A2(KEYINPUT36), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n728), .B(new_n729), .Z(new_n730));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G5), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G171), .B2(new_n731), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1961), .ZN(new_n734));
  MUX2_X1   g309(.A(G19), .B(new_n622), .S(new_n699), .Z(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(G1341), .B2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT102), .B(KEYINPUT24), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G34), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(new_n712), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n476), .B2(new_n712), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G2084), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT30), .B(G28), .ZN(new_n742));
  OR2_X1    g317(.A1(KEYINPUT31), .A2(G11), .ZN(new_n743));
  NAND2_X1  g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n742), .A2(new_n712), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n639), .B2(new_n712), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT103), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n731), .A2(G4), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n611), .B2(new_n731), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n741), .B(new_n747), .C1(G1348), .C2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n698), .A2(G20), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT23), .Z(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G299), .B2(G16), .ZN(new_n753));
  INV_X1    g328(.A(G1956), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n735), .A2(G1341), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n750), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n731), .A2(G21), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G168), .B2(new_n731), .ZN(new_n759));
  INV_X1    g334(.A(G1966), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n712), .A2(G27), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G164), .B2(new_n712), .ZN(new_n763));
  INV_X1    g338(.A(G2078), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n749), .A2(G1348), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n712), .A2(G26), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT28), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n479), .A2(G128), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n459), .A2(G116), .ZN(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n771));
  INV_X1    g346(.A(G140), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n769), .B1(new_n770), .B2(new_n771), .C1(new_n637), .C2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(G29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2067), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n761), .A2(new_n765), .A3(new_n766), .A4(new_n775), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n712), .A2(G33), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT25), .Z(new_n779));
  INV_X1    g354(.A(G139), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n637), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT100), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n464), .A2(G127), .ZN(new_n783));
  AND2_X1   g358(.A1(G115), .A2(G2104), .ZN(new_n784));
  OAI21_X1  g359(.A(G2105), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n777), .B1(new_n786), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT101), .B(G2072), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n776), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n736), .A2(new_n757), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n712), .A2(G32), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n488), .A2(G141), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n468), .A2(G105), .ZN(new_n793));
  NAND3_X1  g368(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT26), .ZN(new_n795));
  AOI211_X1 g370(.A(new_n793), .B(new_n795), .C1(G129), .C2(new_n479), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n791), .B1(new_n798), .B2(new_n712), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT27), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1996), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n787), .B2(new_n788), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n712), .A2(G35), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G162), .B2(new_n712), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT29), .B(G2090), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n790), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n730), .A2(new_n807), .ZN(G150));
  INV_X1    g383(.A(G150), .ZN(G311));
  NAND2_X1  g384(.A1(new_n611), .A2(G559), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT38), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n532), .A2(G93), .B1(new_n534), .B2(G55), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n522), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(new_n527), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n815), .A2(new_n563), .A3(new_n564), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n814), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n622), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n811), .B(new_n819), .Z(new_n820));
  OR2_X1    g395(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  INV_X1    g396(.A(G860), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n817), .A2(G860), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(G145));
  NAND2_X1  g402(.A1(new_n479), .A2(G130), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT104), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n488), .A2(G142), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n459), .A2(G118), .ZN(new_n831));
  OAI21_X1  g406(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n829), .B(new_n830), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n719), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(new_n629), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n797), .B(new_n773), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n786), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n501), .A2(new_n504), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n507), .B2(new_n509), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n837), .B(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT105), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n835), .A2(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n835), .A2(new_n840), .A3(KEYINPUT105), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(G162), .B(new_n639), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n476), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n843), .A2(new_n848), .ZN(new_n851));
  AOI21_X1  g426(.A(G37), .B1(new_n851), .B2(new_n841), .ZN(new_n852));
  AOI21_X1  g427(.A(KEYINPUT40), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n848), .B1(new_n844), .B2(new_n845), .ZN(new_n854));
  INV_X1    g429(.A(new_n852), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT40), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n853), .A2(new_n857), .ZN(G395));
  INV_X1    g433(.A(KEYINPUT42), .ZN(new_n859));
  XOR2_X1   g434(.A(G290), .B(G305), .Z(new_n860));
  XNOR2_X1  g435(.A(G166), .B(G288), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n862), .A2(KEYINPUT107), .ZN(new_n863));
  OAI21_X1  g438(.A(KEYINPUT107), .B1(new_n862), .B2(KEYINPUT108), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n859), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n819), .B(new_n623), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n610), .A2(G299), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n610), .A2(G299), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(KEYINPUT41), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n610), .B(G299), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n878), .A2(new_n867), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n872), .B2(new_n871), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n864), .A2(new_n859), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n866), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n881), .B1(new_n866), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g459(.A(G868), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT109), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n885), .B(new_n886), .C1(G868), .C2(new_n815), .ZN(new_n887));
  INV_X1    g462(.A(new_n882), .ZN(new_n888));
  OAI221_X1 g463(.A(new_n880), .B1(new_n872), .B2(new_n871), .C1(new_n888), .C2(new_n865), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n866), .A2(new_n881), .A3(new_n882), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n616), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n815), .A2(G868), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT109), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n893), .ZN(G295));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n885), .B(new_n895), .C1(G868), .C2(new_n815), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT110), .B1(new_n891), .B2(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n899));
  INV_X1    g474(.A(new_n862), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n819), .A2(G171), .ZN(new_n901));
  NAND3_X1  g476(.A1(G301), .A2(new_n818), .A3(new_n816), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n901), .A2(G168), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(G168), .B1(new_n901), .B2(new_n902), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n903), .A2(new_n878), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n902), .ZN(new_n906));
  AOI21_X1  g481(.A(G301), .B1(new_n818), .B2(new_n816), .ZN(new_n907));
  OAI21_X1  g482(.A(G286), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(G168), .A3(new_n902), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n875), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n900), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n870), .B1(new_n903), .B2(new_n904), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n908), .A2(new_n877), .A3(new_n874), .A4(new_n909), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n862), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT111), .B1(new_n917), .B2(G37), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n915), .A2(new_n916), .A3(new_n862), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n914), .A2(new_n918), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n911), .A2(new_n913), .A3(new_n920), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n899), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n914), .A2(new_n918), .A3(new_n920), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT112), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT43), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n926), .B1(new_n925), .B2(KEYINPUT43), .ZN(new_n928));
  AND4_X1   g503(.A1(new_n919), .A2(new_n911), .A3(new_n913), .A4(new_n920), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n924), .B1(new_n930), .B2(new_n899), .ZN(G397));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n507), .A2(new_n509), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n496), .A2(new_n499), .ZN(new_n934));
  AOI21_X1  g509(.A(G1384), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT113), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n932), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n937), .B1(new_n936), .B2(new_n935), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n469), .B(G40), .C1(new_n474), .C2(new_n475), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n719), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n943), .A2(new_n722), .ZN(new_n944));
  XOR2_X1   g519(.A(new_n773), .B(G2067), .Z(new_n945));
  INV_X1    g520(.A(G1996), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n797), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n722), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n944), .A2(new_n945), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(G290), .B(G1986), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n942), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n508), .B1(new_n484), .B2(G138), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n506), .A2(KEYINPUT4), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n934), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n939), .A2(new_n956), .A3(G2067), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n954), .A2(new_n958), .A3(new_n955), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT114), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT114), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n935), .A2(new_n961), .A3(new_n958), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n939), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT115), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n500), .A2(new_n505), .ZN(new_n965));
  AOI21_X1  g540(.A(G1384), .B1(new_n965), .B2(new_n933), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n964), .B1(new_n966), .B2(new_n958), .ZN(new_n967));
  OAI211_X1 g542(.A(KEYINPUT115), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n963), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G1348), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n957), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT124), .B1(new_n972), .B2(KEYINPUT60), .ZN(new_n973));
  AOI21_X1  g548(.A(G1348), .B1(new_n963), .B2(new_n969), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT124), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT60), .ZN(new_n976));
  NOR4_X1   g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .A4(new_n957), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n973), .A2(new_n977), .A3(new_n610), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n967), .A2(new_n968), .ZN(new_n979));
  NOR4_X1   g554(.A1(new_n839), .A2(KEYINPUT114), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n961), .B1(new_n935), .B2(new_n958), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n940), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n971), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n957), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(KEYINPUT60), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(new_n975), .A3(new_n610), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n976), .B1(new_n974), .B2(new_n957), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT125), .B1(new_n978), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n985), .A2(new_n975), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n972), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n611), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT125), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(new_n993), .A3(new_n987), .A4(new_n986), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n966), .A2(new_n958), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n956), .A2(KEYINPUT50), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n940), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n754), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n935), .A2(KEYINPUT45), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n932), .B1(G164), .B2(G1384), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT56), .B(G2072), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n940), .A2(new_n1000), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G299), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n574), .A2(new_n578), .A3(KEYINPUT57), .A4(new_n580), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n995), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT122), .ZN(new_n1011));
  AND3_X1   g586(.A1(new_n940), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1012), .A2(new_n1002), .B1(new_n998), .B2(new_n754), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1011), .B1(new_n1013), .B2(new_n1008), .ZN(new_n1014));
  AND4_X1   g589(.A1(new_n1011), .A2(new_n999), .A3(new_n1008), .A4(new_n1003), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1010), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT123), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT123), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1018), .B(new_n1010), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n940), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n939), .A2(new_n956), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT58), .B(G1341), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n1021), .A2(G1996), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n563), .A2(KEYINPUT119), .A3(new_n564), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1025), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT59), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT120), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n1027), .ZN(new_n1034));
  NOR3_X1   g609(.A1(new_n1013), .A2(KEYINPUT121), .A3(new_n1008), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(KEYINPUT61), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1013), .A2(new_n1008), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(KEYINPUT121), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1030), .A2(new_n1034), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n989), .A2(new_n994), .A3(new_n1020), .A4(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1038), .B1(new_n972), .B2(new_n610), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1037), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1041), .A2(KEYINPUT126), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT126), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1045));
  NAND3_X1  g620(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1048));
  OR2_X1    g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1021), .A2(new_n702), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(G2090), .B2(new_n998), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1049), .B1(G8), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n970), .A2(G2090), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1054), .B2(new_n1050), .ZN(new_n1055));
  INV_X1    g630(.A(G8), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1022), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1976), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(G288), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT52), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(G288), .B2(new_n1058), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1057), .B(new_n1061), .C1(new_n1058), .C2(G288), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n588), .A2(new_n594), .ZN(new_n1063));
  INV_X1    g638(.A(G1981), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1063), .A2(KEYINPUT116), .A3(new_n1064), .A4(new_n593), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(G305), .B2(G1981), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1065), .A2(new_n1067), .B1(G305), .B2(G1981), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1068), .A2(KEYINPUT49), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1057), .B1(new_n1068), .B2(KEYINPUT49), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1060), .B(new_n1062), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1052), .A2(new_n1055), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1961), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n970), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n965), .A2(new_n933), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1075), .A2(KEYINPUT45), .A3(new_n955), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n932), .B1(new_n839), .B2(G1384), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n940), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n1079));
  OR3_X1    g654(.A1(new_n1078), .A2(new_n1079), .A3(G2078), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1079), .B1(new_n1021), .B2(G2078), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1074), .A2(new_n1080), .A3(G301), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n938), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n764), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n473), .B2(G2105), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1083), .A2(new_n469), .A3(new_n1000), .A4(new_n1085), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1086), .A2(new_n1074), .A3(new_n1081), .ZN(new_n1087));
  OAI211_X1 g662(.A(KEYINPUT54), .B(new_n1082), .C1(new_n1087), .C2(G301), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1072), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(G301), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1074), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G171), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT54), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT127), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1078), .A2(KEYINPUT117), .A3(new_n760), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT117), .B1(new_n1078), .B2(new_n760), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G2084), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n963), .A2(new_n969), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(G286), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1078), .A2(new_n760), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1078), .A2(KEYINPUT117), .A3(new_n760), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1104), .A2(G286), .A3(new_n1100), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(G8), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT51), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT51), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1104), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1110), .B(G8), .C1(new_n1111), .C2(G286), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1095), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(G168), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1056), .B1(new_n1114), .B2(new_n1106), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1095), .B(new_n1112), .C1(new_n1115), .C2(new_n1110), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1094), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1044), .A2(new_n1045), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT62), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1112), .B1(new_n1115), .B2(new_n1110), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT127), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(new_n1123), .A3(new_n1116), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1072), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(new_n1092), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1120), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1128), .A2(G1976), .A3(G288), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1057), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1055), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1132), .B1(new_n1071), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1055), .A2(new_n1071), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1054), .A2(new_n1050), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1135), .B(KEYINPUT63), .C1(new_n1049), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1101), .A2(G8), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1125), .B2(new_n1138), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1134), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1127), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n951), .B1(new_n1119), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n949), .A2(new_n942), .ZN(new_n1145));
  NOR2_X1   g720(.A1(G290), .A2(G1986), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n942), .A2(KEYINPUT48), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT48), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1146), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1148), .B1(new_n941), .B2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1145), .A2(new_n1147), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n945), .A2(new_n947), .ZN(new_n1152));
  OAI22_X1  g727(.A1(new_n944), .A2(new_n1152), .B1(G2067), .B2(new_n773), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n942), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n941), .B1(new_n798), .B2(new_n945), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT46), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n942), .A2(new_n946), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1155), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT47), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1151), .B(new_n1154), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1160), .B2(new_n1159), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1144), .A2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g738(.A(G319), .B(new_n680), .C1(new_n662), .C2(new_n663), .ZN(new_n1165));
  NOR2_X1   g739(.A1(G229), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g740(.A(new_n1166), .B1(new_n854), .B2(new_n855), .ZN(new_n1167));
  NOR2_X1   g741(.A1(new_n930), .A2(new_n1167), .ZN(G308));
  NAND2_X1  g742(.A1(new_n850), .A2(new_n852), .ZN(new_n1169));
  OR2_X1    g743(.A1(new_n928), .A2(new_n929), .ZN(new_n1170));
  OAI211_X1 g744(.A(new_n1169), .B(new_n1166), .C1(new_n1170), .C2(new_n927), .ZN(G225));
endmodule


