//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n535, new_n536, new_n537, new_n538, new_n539, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1126, new_n1127;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G235), .A2(G238), .A3(G237), .A4(G236), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT68), .Z(new_n454));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n468), .B1(new_n465), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n465), .A2(new_n467), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G137), .ZN(new_n475));
  NAND2_X1  g050(.A1(G101), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n473), .A2(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n465), .A2(new_n467), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n463), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n463), .B2(G112), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n481), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT70), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n489), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(new_n469), .B2(new_n470), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n474), .A2(new_n463), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n494), .B2(new_n489), .ZN(new_n495));
  OAI211_X1 g070(.A(KEYINPUT71), .B(new_n490), .C1(new_n469), .C2(new_n470), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n493), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(G114), .A2(G2104), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n479), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n464), .A2(G2105), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n500), .A2(G2105), .B1(G102), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT72), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n497), .A2(new_n505), .A3(new_n502), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n508), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n519), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n516), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT73), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n520), .A2(G51), .ZN(new_n529));
  XNOR2_X1  g104(.A(KEYINPUT74), .B(G89), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n528), .B(new_n529), .C1(new_n523), .C2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XOR2_X1   g107(.A(new_n532), .B(KEYINPUT7), .Z(new_n533));
  NOR2_X1   g108(.A1(new_n531), .A2(new_n533), .ZN(G168));
  NAND2_X1  g109(.A1(new_n520), .A2(G52), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n523), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n515), .B2(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n515), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n520), .A2(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n523), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n549), .A2(new_n552), .ZN(G188));
  NAND3_X1  g128(.A1(new_n509), .A2(new_n511), .A3(G65), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT75), .B1(new_n556), .B2(G651), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  AOI211_X1 g133(.A(new_n558), .B(new_n515), .C1(new_n554), .C2(new_n555), .ZN(new_n559));
  INV_X1    g134(.A(G91), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n557), .A2(new_n559), .B1(new_n560), .B2(new_n523), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(KEYINPUT9), .B1(new_n520), .B2(G53), .ZN(new_n563));
  INV_X1    g138(.A(new_n519), .ZN(new_n564));
  OAI211_X1 g139(.A(G53), .B(G543), .C1(new_n564), .C2(new_n517), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n562), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G168), .ZN(G286));
  INV_X1    g145(.A(G166), .ZN(G303));
  INV_X1    g146(.A(new_n523), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n520), .A2(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  AOI22_X1  g151(.A1(new_n513), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n515), .ZN(new_n578));
  NAND2_X1  g153(.A1(G48), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G86), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n512), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(new_n522), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(G72), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G60), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n512), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT76), .Z(new_n588));
  AOI21_X1  g163(.A(new_n588), .B1(G47), .B2(new_n520), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n572), .A2(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  AND3_X1   g167(.A1(new_n513), .A2(G92), .A3(new_n522), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n520), .A2(G54), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n513), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n515), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n592), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n592), .B1(new_n599), .B2(G868), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G299), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G168), .B2(new_n602), .ZN(G297));
  OAI21_X1  g179(.A(new_n603), .B1(G168), .B2(new_n602), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n599), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n609), .A2(KEYINPUT77), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(KEYINPUT77), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n610), .B(new_n611), .C1(G868), .C2(new_n547), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g188(.A1(new_n469), .A2(new_n470), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n501), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT78), .B(KEYINPUT12), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT13), .B(G2100), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n480), .A2(G123), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n482), .A2(G135), .ZN(new_n621));
  NOR2_X1   g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND2_X1  g200(.A1(new_n619), .A2(new_n625), .ZN(G156));
  INV_X1    g201(.A(G14), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT79), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n634), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  NOR2_X1   g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT80), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(KEYINPUT80), .ZN(new_n643));
  AOI211_X1 g218(.A(new_n627), .B(new_n640), .C1(new_n642), .C2(new_n643), .ZN(G401));
  XOR2_X1   g219(.A(KEYINPUT81), .B(KEYINPUT18), .Z(new_n645));
  XOR2_X1   g220(.A(G2067), .B(G2678), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  OAI21_X1  g223(.A(KEYINPUT17), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n648), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n650), .A2(new_n646), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n645), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n652), .B(new_n653), .C1(new_n651), .C2(new_n645), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2096), .B(G2100), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  AND2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n660), .A2(KEYINPUT82), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(KEYINPUT82), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n661), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n658), .A2(new_n659), .ZN(new_n669));
  OR3_X1    g244(.A1(new_n664), .A2(new_n660), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n666), .A2(new_n667), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n664), .A2(new_n669), .ZN(new_n672));
  NAND4_X1  g247(.A1(new_n668), .A2(new_n670), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1986), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1981), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1991), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G229));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G25), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n480), .A2(G119), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n482), .A2(G131), .ZN(new_n683));
  OR2_X1    g258(.A1(G95), .A2(G2105), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n684), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n681), .B1(new_n687), .B2(new_n680), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT35), .B(G1991), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n691), .A2(G24), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G290), .B2(G16), .ZN(new_n693));
  INV_X1    g268(.A(G1986), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n690), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(G23), .ZN(new_n696));
  INV_X1    g271(.A(G288), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(new_n691), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT33), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1976), .ZN(new_n700));
  MUX2_X1   g275(.A(G6), .B(G305), .S(G16), .Z(new_n701));
  XOR2_X1   g276(.A(KEYINPUT32), .B(G1981), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n691), .A2(G22), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n691), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT83), .B(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n700), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n695), .B1(new_n708), .B2(KEYINPUT34), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(KEYINPUT34), .B2(new_n708), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n694), .B2(new_n693), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT84), .B(KEYINPUT36), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(G168), .A2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G16), .B2(G21), .ZN(new_n715));
  INV_X1    g290(.A(G1966), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n547), .A2(new_n691), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n691), .B2(G19), .ZN(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n715), .A2(new_n716), .B1(new_n719), .B2(G1341), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n691), .A2(G4), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n599), .B2(new_n691), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G1348), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n720), .B(new_n723), .C1(new_n716), .C2(new_n715), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n719), .A2(G1341), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G5), .B2(G16), .ZN(new_n727));
  OR3_X1    g302(.A1(new_n726), .A2(G5), .A3(G16), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n727), .B(new_n728), .C1(G301), .C2(new_n691), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT93), .ZN(new_n730));
  INV_X1    g305(.A(G1961), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n680), .B1(new_n733), .B2(G28), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(KEYINPUT91), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(G28), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n734), .A2(KEYINPUT91), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n738), .B1(new_n680), .B2(new_n624), .C1(new_n722), .C2(G1348), .ZN(new_n739));
  NOR4_X1   g314(.A1(new_n724), .A2(new_n725), .A3(new_n732), .A4(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(KEYINPUT24), .A2(G34), .ZN(new_n741));
  NOR2_X1   g316(.A1(KEYINPUT24), .A2(G34), .ZN(new_n742));
  NOR3_X1   g317(.A1(new_n741), .A2(new_n742), .A3(G29), .ZN(new_n743));
  INV_X1    g318(.A(G160), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G29), .ZN(new_n745));
  INV_X1    g320(.A(G2084), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT85), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n730), .A2(new_n731), .ZN(new_n749));
  OR2_X1    g324(.A1(G29), .A2(G33), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n482), .A2(G139), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n501), .A2(G103), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT25), .Z(new_n753));
  AOI22_X1  g328(.A1(new_n614), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n751), .B(new_n753), .C1(new_n754), .C2(new_n463), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n750), .B1(new_n755), .B2(new_n680), .ZN(new_n756));
  INV_X1    g331(.A(G2072), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n745), .A2(new_n746), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n680), .A2(G26), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n480), .A2(G128), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n482), .A2(G140), .ZN(new_n762));
  NOR2_X1   g337(.A1(G104), .A2(G2105), .ZN(new_n763));
  OAI21_X1  g338(.A(G2104), .B1(new_n463), .B2(G116), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n761), .B(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n760), .B1(new_n765), .B2(G29), .ZN(new_n766));
  MUX2_X1   g341(.A(new_n760), .B(new_n766), .S(KEYINPUT28), .Z(new_n767));
  INV_X1    g342(.A(G2067), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n749), .A2(new_n758), .A3(new_n759), .A4(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n768), .B2(new_n767), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT31), .B(G11), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n740), .A2(new_n748), .A3(new_n771), .A4(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G27), .A2(G29), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G164), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2078), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT94), .B(KEYINPUT23), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n691), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G299), .B2(G16), .ZN(new_n780));
  INV_X1    g355(.A(G1956), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(G29), .A2(G35), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G162), .B2(G29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT29), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2090), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n773), .A2(new_n776), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n756), .A2(new_n757), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT86), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n480), .A2(G129), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT88), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n482), .A2(G141), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT87), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT26), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n501), .A2(G105), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n791), .A2(new_n794), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT89), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G29), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(KEYINPUT90), .C1(G29), .C2(G32), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(KEYINPUT90), .B2(new_n800), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT27), .B(G1996), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n713), .A2(new_n787), .A3(new_n789), .A4(new_n804), .ZN(G150));
  INV_X1    g380(.A(G150), .ZN(G311));
  AOI22_X1  g381(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n515), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n520), .A2(G55), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT95), .B(G93), .Z(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n523), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G860), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT96), .B(KEYINPUT97), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT37), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n599), .A2(G559), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n547), .B(new_n812), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT39), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n817), .B1(new_n822), .B2(G860), .ZN(G145));
  MUX2_X1   g398(.A(new_n799), .B(new_n798), .S(new_n755), .Z(new_n824));
  XOR2_X1   g399(.A(new_n503), .B(new_n765), .Z(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(G130), .A2(new_n480), .B1(new_n482), .B2(G142), .ZN(new_n827));
  OAI21_X1  g402(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(KEYINPUT98), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(KEYINPUT98), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n829), .B(new_n830), .C1(G118), .C2(new_n463), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n687), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(new_n617), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n826), .B(new_n834), .Z(new_n835));
  XNOR2_X1  g410(.A(G160), .B(new_n624), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n487), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT99), .ZN(new_n839));
  INV_X1    g414(.A(G37), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n841));
  OR3_X1    g416(.A1(new_n826), .A2(new_n841), .A3(new_n834), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n826), .B1(new_n841), .B2(new_n834), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n842), .A2(new_n837), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n839), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT40), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n839), .A2(new_n847), .A3(new_n840), .A4(new_n844), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G395));
  NOR2_X1   g424(.A1(new_n813), .A2(G868), .ZN(new_n850));
  XNOR2_X1  g425(.A(G290), .B(G288), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n851), .A2(KEYINPUT103), .ZN(new_n852));
  XNOR2_X1  g427(.A(G303), .B(G305), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(KEYINPUT103), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OR3_X1    g431(.A1(new_n851), .A2(KEYINPUT103), .A3(new_n854), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT42), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n820), .B(KEYINPUT101), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n608), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n598), .B(G299), .Z(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n865));
  NOR3_X1   g440(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT41), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n863), .B(KEYINPUT41), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n866), .B1(new_n867), .B2(new_n865), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n864), .B2(new_n862), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n860), .A2(KEYINPUT104), .A3(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n870), .A2(KEYINPUT104), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n870), .A2(KEYINPUT104), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n859), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n850), .B1(new_n875), .B2(G868), .ZN(G331));
  XNOR2_X1  g451(.A(G331), .B(KEYINPUT105), .ZN(G295));
  XNOR2_X1  g452(.A(G168), .B(G301), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(KEYINPUT106), .A3(new_n820), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n878), .B(new_n820), .Z(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n879), .B1(new_n881), .B2(KEYINPUT106), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(new_n863), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n868), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n886), .A3(new_n858), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n858), .A2(new_n886), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(new_n884), .A3(new_n883), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(new_n840), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT43), .ZN(new_n891));
  OAI22_X1  g466(.A1(new_n882), .A2(new_n867), .B1(new_n864), .B2(new_n881), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n858), .ZN(new_n893));
  OAI211_X1 g468(.A(new_n893), .B(new_n840), .C1(new_n858), .C2(new_n885), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n894), .B2(KEYINPUT43), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n894), .B2(new_n896), .ZN(new_n898));
  MUX2_X1   g473(.A(new_n895), .B(new_n898), .S(KEYINPUT44), .Z(G397));
  INV_X1    g474(.A(KEYINPUT46), .ZN(new_n900));
  INV_X1    g475(.A(G1384), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n503), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g480(.A(KEYINPUT109), .B(G40), .Z(new_n906));
  NOR3_X1   g481(.A1(new_n473), .A2(new_n477), .A3(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n900), .B1(new_n910), .B2(G1996), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n765), .B(new_n768), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n909), .B1(new_n798), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G1996), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n909), .A2(KEYINPUT46), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n911), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n917), .B(KEYINPUT47), .Z(new_n918));
  AND2_X1   g493(.A1(new_n798), .A2(G1996), .ZN(new_n919));
  AOI211_X1 g494(.A(new_n913), .B(new_n919), .C1(new_n799), .C2(new_n915), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n920), .A2(new_n689), .A3(new_n687), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n765), .A2(G2067), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n909), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n923), .B(KEYINPUT127), .Z(new_n924));
  XNOR2_X1  g499(.A(new_n686), .B(new_n689), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n909), .ZN(new_n927));
  NOR2_X1   g502(.A1(G290), .A2(G1986), .ZN(new_n928));
  XOR2_X1   g503(.A(new_n928), .B(KEYINPUT110), .Z(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n909), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT48), .ZN(new_n931));
  AOI211_X1 g506(.A(new_n918), .B(new_n924), .C1(new_n927), .C2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT57), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT114), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n934), .B1(new_n563), .B2(new_n567), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n520), .A2(KEYINPUT9), .A3(G53), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n565), .A2(new_n566), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT114), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n933), .B1(new_n939), .B2(new_n561), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT115), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n562), .A2(KEYINPUT57), .A3(new_n568), .ZN(new_n943));
  OAI211_X1 g518(.A(KEYINPUT115), .B(new_n933), .C1(new_n939), .C2(new_n561), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT116), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT116), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n942), .A2(new_n943), .A3(new_n947), .A4(new_n944), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n504), .A2(new_n950), .A3(new_n901), .A4(new_n506), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n902), .A2(KEYINPUT50), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n907), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n781), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n504), .A2(new_n901), .A3(new_n506), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n904), .ZN(new_n956));
  AOI21_X1  g531(.A(G1384), .B1(new_n497), .B2(new_n502), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(KEYINPUT45), .ZN(new_n958));
  XNOR2_X1  g533(.A(KEYINPUT56), .B(G2072), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n956), .A2(new_n907), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n949), .A2(new_n954), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT117), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n949), .A2(new_n954), .A3(new_n960), .A4(KEYINPUT117), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n954), .A2(new_n960), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT119), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n949), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n954), .A2(new_n960), .A3(KEYINPUT119), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n955), .A2(KEYINPUT50), .ZN(new_n972));
  AOI211_X1 g547(.A(KEYINPUT50), .B(G1384), .C1(new_n497), .C2(new_n502), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n907), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT118), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G1348), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n972), .A2(KEYINPUT118), .A3(new_n907), .A4(new_n974), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n902), .A2(new_n908), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n768), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n598), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n963), .B(new_n964), .C1(new_n971), .C2(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n980), .A2(new_n598), .A3(new_n982), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT60), .B1(new_n985), .B2(new_n983), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT60), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n980), .A2(new_n987), .A3(new_n599), .A4(new_n982), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n956), .A2(new_n907), .A3(new_n958), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n990), .B(G1341), .ZN(new_n991));
  OAI22_X1  g566(.A1(new_n989), .A2(G1996), .B1(new_n981), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n547), .ZN(new_n993));
  NOR2_X1   g568(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(new_n994), .ZN(new_n996));
  NAND2_X1  g571(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n992), .A2(new_n547), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n988), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n986), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT61), .B1(new_n965), .B2(new_n968), .ZN(new_n1001));
  AND3_X1   g576(.A1(new_n1001), .A2(new_n963), .A3(new_n964), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n961), .A2(KEYINPUT122), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n961), .A2(KEYINPUT122), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n970), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1002), .B1(new_n1005), .B2(KEYINPUT61), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n984), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT123), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  AOI211_X1 g584(.A(new_n908), .B(new_n973), .C1(new_n955), .C2(KEYINPUT50), .ZN(new_n1010));
  INV_X1    g585(.A(G2090), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1971), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n989), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1009), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(G303), .A2(G8), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT55), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT111), .B(G8), .Z(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  NOR2_X1   g597(.A1(G288), .A2(new_n1022), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n981), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1024), .B(new_n1025), .C1(G1976), .C2(new_n697), .ZN(new_n1026));
  XNOR2_X1  g601(.A(G305), .B(G1981), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT49), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n981), .A2(new_n1021), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1029), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1026), .B(new_n1032), .C1(new_n1025), .C2(new_n1024), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n908), .B1(new_n955), .B2(new_n904), .ZN(new_n1035));
  AOI21_X1  g610(.A(G1971), .B1(new_n1035), .B2(new_n958), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n953), .A2(G2090), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1020), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1017), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1019), .A2(new_n1034), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n989), .B2(G2078), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n977), .A2(new_n731), .A3(new_n979), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n907), .B1(new_n957), .B2(KEYINPUT45), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT112), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1041), .A2(G2078), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n504), .A2(new_n901), .A3(new_n506), .A4(new_n903), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1049), .B(new_n907), .C1(new_n957), .C2(KEYINPUT45), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1044), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT125), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1044), .A2(KEYINPUT125), .A3(new_n1051), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1043), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(G301), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n744), .B1(new_n957), .B2(KEYINPUT45), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n905), .A2(new_n1059), .A3(G40), .A4(new_n1047), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1044), .A2(new_n1042), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1058), .B1(new_n1061), .B2(G171), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1040), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n1061), .A2(G171), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n1056), .B2(G301), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT124), .ZN(new_n1066));
  NOR2_X1   g641(.A1(G168), .A2(new_n1021), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1046), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1010), .A2(new_n746), .B1(new_n1069), .B2(new_n716), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1068), .B1(new_n1070), .B2(new_n1009), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n716), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n972), .A2(new_n746), .A3(new_n907), .A4(new_n974), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1020), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1067), .A2(KEYINPUT51), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1071), .A2(KEYINPUT51), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1070), .A2(new_n1068), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1066), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1009), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT51), .B1(new_n1080), .B2(new_n1067), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1076), .B1(new_n1070), .B2(new_n1021), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1078), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(KEYINPUT124), .A3(new_n1084), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1065), .A2(new_n1058), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1087), .B(new_n984), .C1(new_n1000), .C2(new_n1006), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1008), .A2(new_n1063), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT63), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1075), .A2(G286), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1090), .B1(new_n1040), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1017), .A2(KEYINPUT113), .ZN(new_n1094));
  OR2_X1    g669(.A1(new_n1015), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1090), .B1(new_n1015), .B2(new_n1094), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1034), .A4(new_n1091), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1093), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1034), .A2(new_n1018), .A3(new_n1015), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1032), .A2(new_n1022), .A3(new_n697), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(G1981), .B2(G305), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1030), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1098), .A2(new_n1099), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT124), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1104));
  AOI211_X1 g679(.A(new_n1066), .B(new_n1078), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1040), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1055), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT125), .B1(new_n1044), .B2(new_n1051), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1042), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(G171), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1079), .A2(new_n1085), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(KEYINPUT62), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1103), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1089), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n929), .B1(G1986), .B2(G290), .ZN(new_n1117));
  INV_X1    g692(.A(new_n926), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n910), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT126), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT126), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1122), .B(new_n1119), .C1(new_n1089), .C2(new_n1115), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n932), .B1(new_n1121), .B2(new_n1123), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g699(.A1(G229), .A2(new_n461), .ZN(new_n1126));
  NOR2_X1   g700(.A1(G401), .A2(G227), .ZN(new_n1127));
  AND4_X1   g701(.A1(new_n845), .A2(new_n895), .A3(new_n1126), .A4(new_n1127), .ZN(G308));
  NAND4_X1  g702(.A1(new_n845), .A2(new_n895), .A3(new_n1126), .A4(new_n1127), .ZN(G225));
endmodule


