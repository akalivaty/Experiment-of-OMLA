//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G116), .A2(G270), .ZN(new_n210));
  XNOR2_X1  g0010(.A(KEYINPUT65), .B(G238), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(new_n212), .A2(G68), .B1(G77), .B2(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G97), .A2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G50), .A2(G226), .ZN(new_n219));
  AND4_X1   g0019(.A1(new_n210), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G87), .A2(G250), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n209), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  INV_X1    g0023(.A(G13), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n209), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  INV_X1    g0028(.A(new_n201), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n230), .A2(new_n208), .A3(new_n231), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n223), .A2(new_n228), .A3(new_n232), .ZN(G361));
  XOR2_X1   g0033(.A(G226), .B(G232), .Z(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT67), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n231), .ZN(new_n252));
  XOR2_X1   g0052(.A(KEYINPUT8), .B(G58), .Z(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n254), .A2(new_n257), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n208), .B1(new_n201), .B2(new_n202), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n262), .B(KEYINPUT68), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n252), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n252), .B1(new_n207), .B2(G20), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G50), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT9), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G222), .A2(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G223), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G1), .A3(G13), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n275), .B(new_n278), .C1(G77), .C2(new_n271), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n280));
  INV_X1    g0080(.A(G274), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G226), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n277), .A2(new_n280), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n279), .B(new_n283), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G200), .ZN(new_n287));
  INV_X1    g0087(.A(G190), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n270), .B(new_n287), .C1(new_n288), .C2(new_n286), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT10), .ZN(new_n290));
  OR2_X1    g0090(.A1(new_n286), .A2(G179), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n286), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n269), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT13), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n284), .A2(new_n273), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n215), .A2(G1698), .ZN(new_n299));
  AND2_X1   g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  NOR2_X1   g0100(.A1(KEYINPUT3), .A2(G33), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n298), .B(new_n299), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G97), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n282), .B1(new_n304), .B2(new_n278), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n277), .A2(G238), .A3(new_n280), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n297), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n277), .B1(new_n302), .B2(new_n303), .ZN(new_n309));
  NOR4_X1   g0109(.A1(new_n309), .A2(KEYINPUT13), .A3(new_n306), .A4(new_n282), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT14), .B1(new_n311), .B2(new_n292), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT14), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n313), .B(G169), .C1(new_n308), .C2(new_n310), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT74), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n311), .B2(G179), .ZN(new_n316));
  INV_X1    g0116(.A(G179), .ZN(new_n317));
  NOR4_X1   g0117(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT74), .A4(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n312), .B(new_n314), .C1(new_n316), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n265), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT12), .ZN(new_n321));
  INV_X1    g0121(.A(G68), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT73), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT70), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n265), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n207), .A2(KEYINPUT70), .A3(G13), .A4(G20), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n321), .B1(new_n328), .B2(new_n322), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n328), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(G68), .A3(new_n267), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n208), .A2(G33), .A3(G77), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n322), .A2(G20), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n333), .B(new_n334), .C1(new_n260), .C2(new_n202), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT72), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n335), .A2(new_n336), .A3(new_n252), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n335), .B2(new_n252), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT11), .ZN(new_n339));
  OR3_X1    g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n337), .B2(new_n338), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n330), .A2(new_n332), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n319), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n342), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n311), .A2(G190), .ZN(new_n345));
  INV_X1    g0145(.A(G200), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n344), .B(new_n345), .C1(new_n346), .C2(new_n311), .ZN(new_n347));
  INV_X1    g0147(.A(new_n252), .ZN(new_n348));
  XNOR2_X1  g0148(.A(KEYINPUT15), .B(G87), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT69), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n350), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(new_n256), .A3(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n253), .A2(new_n259), .B1(G20), .B2(G77), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n348), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND4_X1   g0155(.A1(G77), .A2(new_n267), .A3(new_n326), .A4(new_n327), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n331), .A2(G77), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n271), .A2(G232), .A3(new_n273), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n300), .A2(new_n301), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G107), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n271), .A2(G1698), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n359), .B(new_n361), .C1(new_n362), .C2(new_n211), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n278), .ZN(new_n364));
  INV_X1    g0164(.A(new_n285), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G244), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n364), .A2(new_n317), .A3(new_n283), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT71), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n282), .B1(new_n363), .B2(new_n278), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT71), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n369), .A2(new_n370), .A3(new_n317), .A4(new_n366), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n358), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n369), .A2(new_n366), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n292), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(G200), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n376), .B(new_n358), .C1(new_n288), .C2(new_n373), .ZN(new_n377));
  AND4_X1   g0177(.A1(new_n343), .A2(new_n347), .A3(new_n375), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT75), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT17), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT16), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G58), .A2(G68), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n208), .B1(new_n229), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT3), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n255), .ZN(new_n385));
  NAND2_X1  g0185(.A1(KEYINPUT3), .A2(G33), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n208), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n385), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n386), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n383), .B1(new_n391), .B2(G68), .ZN(new_n392));
  INV_X1    g0192(.A(G159), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n260), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n381), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n322), .B1(new_n389), .B2(new_n390), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n397), .A2(KEYINPUT16), .A3(new_n394), .A4(new_n383), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n252), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n254), .A2(new_n320), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n267), .A2(new_n253), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n284), .A2(G1698), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n271), .B(new_n402), .C1(G223), .C2(G1698), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n277), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n282), .B1(new_n365), .B2(G232), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n288), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n407), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n346), .B1(new_n409), .B2(new_n405), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n399), .A2(new_n400), .A3(new_n401), .A4(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n379), .A2(KEYINPUT17), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n380), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n379), .A3(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n292), .B1(new_n409), .B2(new_n405), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n406), .A2(new_n317), .A3(new_n407), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n418), .A2(KEYINPUT18), .A3(new_n419), .A4(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n296), .A2(new_n378), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n360), .A2(G20), .ZN(new_n430));
  NOR2_X1   g0230(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n431), .B(KEYINPUT80), .ZN(new_n432));
  NAND2_X1  g0232(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n430), .A2(new_n432), .A3(G87), .A4(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT80), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n431), .B(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n271), .A2(new_n208), .A3(G87), .ZN(new_n437));
  INV_X1    g0237(.A(new_n433), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G116), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n208), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n208), .A2(G107), .ZN(new_n444));
  XNOR2_X1  g0244(.A(new_n444), .B(KEYINPUT23), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n440), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT24), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n434), .A2(new_n439), .B1(new_n208), .B2(new_n442), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT24), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n449), .A3(new_n445), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n348), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(G257), .B(G1698), .C1(new_n300), .C2(new_n301), .ZN(new_n452));
  OAI211_X1 g0252(.A(G250), .B(new_n273), .C1(new_n300), .C2(new_n301), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G294), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n278), .ZN(new_n456));
  INV_X1    g0256(.A(G45), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G1), .ZN(new_n458));
  INV_X1    g0258(.A(G41), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT5), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G41), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n458), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(new_n281), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT5), .B(G41), .ZN(new_n466));
  INV_X1    g0266(.A(new_n231), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n466), .A2(new_n458), .B1(new_n467), .B2(new_n276), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G264), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n456), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G200), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n470), .A2(G190), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n252), .B1(new_n207), .B2(G33), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n265), .ZN(new_n476));
  INV_X1    g0276(.A(G107), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n320), .A2(KEYINPUT25), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT25), .B1(new_n320), .B2(new_n477), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n476), .A2(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n451), .A2(new_n474), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n471), .A2(new_n317), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n470), .A2(new_n292), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND4_X1   g0285(.A1(new_n449), .A2(new_n440), .A3(new_n443), .A4(new_n445), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n449), .B1(new_n448), .B2(new_n445), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n252), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n481), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT81), .B1(new_n482), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n488), .B(new_n489), .C1(new_n473), .C2(new_n472), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n483), .B(new_n484), .C1(new_n451), .C2(new_n481), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT81), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(G244), .B(new_n273), .C1(new_n300), .C2(new_n301), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n271), .A2(KEYINPUT4), .A3(G244), .A4(new_n273), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G283), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n499), .A2(new_n500), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n278), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n463), .A2(G257), .A3(new_n277), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n504), .A2(G179), .A3(new_n465), .A4(new_n506), .ZN(new_n507));
  AOI211_X1 g0307(.A(new_n464), .B(new_n505), .C1(new_n503), .C2(new_n278), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n292), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n265), .A2(G97), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT7), .B1(new_n360), .B2(new_n208), .ZN(new_n511));
  INV_X1    g0311(.A(new_n390), .ZN(new_n512));
  OAI21_X1  g0312(.A(G107), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n260), .A2(new_n203), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT6), .ZN(new_n515));
  AND2_X1   g0315(.A1(G97), .A2(G107), .ZN(new_n516));
  NOR2_X1   g0316(.A1(G97), .A2(G107), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n477), .A2(KEYINPUT6), .A3(G97), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n514), .B1(new_n520), .B2(G20), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n513), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n510), .B1(new_n522), .B2(new_n252), .ZN(new_n523));
  INV_X1    g0323(.A(G97), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n476), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT76), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n348), .B1(new_n513), .B2(new_n521), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT76), .ZN(new_n529));
  NOR4_X1   g0329(.A1(new_n528), .A2(new_n529), .A3(new_n525), .A4(new_n510), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n509), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n430), .A2(G68), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n257), .B2(new_n524), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n208), .B1(new_n303), .B2(new_n533), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT78), .ZN(new_n536));
  XNOR2_X1  g0336(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NOR3_X1   g0337(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n532), .B(new_n534), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n351), .A2(new_n352), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n539), .A2(new_n252), .B1(new_n328), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g0341(.A1(G238), .A2(G1698), .ZN(new_n542));
  INV_X1    g0342(.A(G244), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G1698), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n542), .B(new_n544), .C1(new_n300), .C2(new_n301), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n277), .B1(new_n545), .B2(new_n441), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n207), .A2(G45), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(new_n281), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n277), .A2(G250), .A3(new_n547), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n546), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G190), .ZN(new_n552));
  INV_X1    g0352(.A(new_n548), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n545), .A2(new_n441), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n553), .B(new_n549), .C1(new_n554), .C2(new_n277), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G200), .ZN(new_n556));
  INV_X1    g0356(.A(new_n476), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G87), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n541), .A2(new_n552), .A3(new_n556), .A4(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n504), .A2(new_n465), .A3(new_n506), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G200), .ZN(new_n561));
  NOR3_X1   g0361(.A1(new_n528), .A2(new_n525), .A3(new_n510), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n561), .B(new_n562), .C1(new_n288), .C2(new_n560), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT77), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n551), .A2(G169), .ZN(new_n565));
  NOR4_X1   g0365(.A1(new_n546), .A2(new_n550), .A3(G179), .A4(new_n548), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n566), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n555), .A2(new_n292), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT77), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n539), .A2(new_n252), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n540), .A2(new_n328), .ZN(new_n572));
  INV_X1    g0372(.A(new_n540), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n557), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n571), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n567), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n531), .A2(new_n559), .A3(new_n563), .A4(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(G116), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n328), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n331), .A2(G116), .A3(new_n475), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n501), .B(new_n208), .C1(G33), .C2(new_n524), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n581), .B(new_n252), .C1(new_n208), .C2(G116), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT20), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n579), .B(new_n580), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(G257), .B(new_n273), .C1(new_n300), .C2(new_n301), .ZN(new_n587));
  OAI211_X1 g0387(.A(G264), .B(G1698), .C1(new_n300), .C2(new_n301), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n385), .A2(G303), .A3(new_n386), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(new_n278), .B1(new_n468), .B2(G270), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n465), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n586), .A2(G169), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT21), .ZN(new_n594));
  OR2_X1    g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  INV_X1    g0396(.A(new_n586), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n590), .A2(new_n278), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n468), .A2(G270), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n598), .A2(G179), .A3(new_n465), .A4(new_n599), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n592), .A2(G200), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n597), .B(new_n602), .C1(new_n288), .C2(new_n592), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n595), .A2(new_n596), .A3(new_n601), .A4(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n577), .A2(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n429), .A2(new_n496), .A3(new_n605), .ZN(G372));
  NAND3_X1  g0406(.A1(new_n347), .A2(new_n374), .A3(new_n372), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n343), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(new_n417), .B1(new_n423), .B2(new_n424), .ZN(new_n609));
  INV_X1    g0409(.A(new_n290), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n294), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n611), .B(KEYINPUT83), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n595), .A2(new_n596), .A3(new_n601), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n492), .B1(new_n490), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n531), .A2(new_n559), .A3(new_n563), .ZN(new_n615));
  OR2_X1    g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT82), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n575), .B1(new_n617), .B2(new_n569), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n568), .B1(new_n565), .B2(KEYINPUT82), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n559), .B1(new_n618), .B2(new_n619), .ZN(new_n621));
  INV_X1    g0421(.A(new_n562), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n509), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g0423(.A1(new_n621), .A2(KEYINPUT26), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n559), .B(new_n509), .C1(new_n527), .C2(new_n530), .ZN(new_n626));
  INV_X1    g0426(.A(new_n576), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT26), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n616), .A2(new_n620), .A3(new_n625), .A4(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n612), .B1(new_n428), .B2(new_n630), .ZN(G369));
  NOR2_X1   g0431(.A1(new_n224), .A2(G20), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n207), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G213), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n451), .B2(new_n481), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n496), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n638), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n493), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n597), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n613), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n604), .B2(new_n643), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n645), .A2(G330), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n490), .A2(new_n641), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n613), .A2(new_n641), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n496), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(G399));
  NOR2_X1   g0451(.A1(new_n225), .A2(G41), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n538), .A2(new_n578), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n653), .A2(G1), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n230), .B2(new_n653), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n657), .B(KEYINPUT28), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n620), .B1(new_n614), .B2(new_n615), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT26), .B1(new_n621), .B2(new_n623), .ZN(new_n660));
  INV_X1    g0460(.A(new_n531), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(new_n559), .A3(new_n576), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n660), .B1(new_n662), .B2(KEYINPUT26), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n641), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT29), .ZN(new_n665));
  OAI211_X1 g0465(.A(new_n620), .B(new_n628), .C1(new_n614), .C2(new_n615), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n641), .B1(new_n666), .B2(new_n624), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n665), .B1(KEYINPUT29), .B2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n605), .A2(new_n491), .A3(new_n495), .A4(new_n641), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n600), .A2(new_n555), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n505), .B1(new_n503), .B2(new_n278), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n670), .A2(KEYINPUT30), .A3(new_n471), .A4(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT30), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n455), .A2(new_n278), .B1(new_n468), .B2(G264), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n504), .A2(new_n465), .A3(new_n674), .A4(new_n506), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n551), .A2(new_n591), .A3(G179), .A4(new_n465), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n673), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n465), .B1(new_n674), .B2(new_n591), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n678), .A2(new_n560), .A3(new_n317), .A4(new_n555), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n672), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n638), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT31), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n680), .A2(KEYINPUT31), .A3(new_n638), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n669), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n668), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n658), .B1(new_n688), .B2(G1), .ZN(G364));
  NAND2_X1  g0489(.A1(new_n632), .A2(G45), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n653), .A2(G1), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n646), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(G330), .B2(new_n645), .ZN(new_n694));
  NOR2_X1   g0494(.A1(G13), .A2(G33), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(G20), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n645), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n208), .A2(new_n288), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n317), .A2(G200), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT86), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n702), .A2(new_n703), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G322), .ZN(new_n709));
  XOR2_X1   g0509(.A(KEYINPUT33), .B(G317), .Z(new_n710));
  NOR2_X1   g0510(.A1(new_n317), .A2(new_n346), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n208), .A2(G190), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n346), .A2(G179), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n700), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G303), .ZN(new_n717));
  NOR2_X1   g0517(.A1(G179), .A2(G200), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G329), .ZN(new_n720));
  OAI22_X1  g0520(.A1(new_n716), .A2(new_n717), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n700), .A2(new_n711), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI211_X1 g0523(.A(new_n714), .B(new_n721), .C1(G326), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n712), .A2(new_n701), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G311), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n712), .A2(new_n715), .ZN(new_n728));
  INV_X1    g0528(.A(G283), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n208), .B1(new_n718), .B2(G190), .ZN(new_n730));
  INV_X1    g0530(.A(G294), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n728), .A2(new_n729), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n271), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n709), .A2(new_n724), .A3(new_n727), .A4(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n716), .ZN(new_n735));
  AOI22_X1  g0535(.A1(G87), .A2(new_n735), .B1(new_n726), .B2(G77), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n322), .B2(new_n713), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n728), .A2(new_n477), .ZN(new_n738));
  NOR3_X1   g0538(.A1(new_n737), .A2(new_n360), .A3(new_n738), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n708), .A2(G58), .B1(G50), .B2(new_n723), .ZN(new_n740));
  INV_X1    g0540(.A(new_n730), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G97), .ZN(new_n742));
  INV_X1    g0542(.A(new_n719), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G159), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(KEYINPUT32), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n739), .A2(new_n740), .A3(new_n742), .A4(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n744), .A2(KEYINPUT32), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n734), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AND2_X1   g0548(.A1(KEYINPUT85), .A2(G169), .ZN(new_n749));
  NOR2_X1   g0549(.A1(KEYINPUT85), .A2(G169), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n749), .A2(new_n750), .A3(new_n208), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n231), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n225), .A2(new_n271), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n246), .B2(G45), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(G45), .B2(new_n230), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n225), .A2(new_n360), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT84), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G355), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n757), .B(new_n760), .C1(G116), .C2(new_n226), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n752), .A2(new_n697), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n699), .A2(new_n753), .A3(new_n763), .A4(new_n692), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n694), .A2(new_n764), .ZN(G396));
  INV_X1    g0565(.A(new_n358), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n638), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n375), .A2(new_n377), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n368), .A2(new_n371), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n769), .A2(new_n374), .A3(new_n766), .A4(new_n638), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT91), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n372), .A2(KEYINPUT91), .A3(new_n374), .A4(new_n638), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n768), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT92), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n768), .A2(KEYINPUT92), .A3(new_n772), .A4(new_n773), .ZN(new_n777));
  AND2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n667), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n776), .A2(new_n777), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n629), .A2(new_n780), .A3(new_n641), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n687), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n691), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(KEYINPUT93), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n781), .A2(new_n779), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n686), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT93), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n782), .A2(new_n787), .A3(new_n691), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n784), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT94), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n778), .A2(new_n695), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n716), .A2(new_n477), .ZN(new_n792));
  INV_X1    g0592(.A(new_n713), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT87), .B(G283), .Z(new_n794));
  AOI22_X1  g0594(.A1(new_n793), .A2(new_n794), .B1(new_n726), .B2(G116), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT88), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n792), .B(new_n796), .C1(G294), .C2(new_n708), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n271), .B1(new_n723), .B2(G303), .ZN(new_n798));
  INV_X1    g0598(.A(G87), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n728), .A2(new_n799), .B1(new_n719), .B2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT89), .Z(new_n802));
  NAND4_X1  g0602(.A1(new_n797), .A2(new_n742), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G137), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n722), .A2(new_n804), .B1(new_n713), .B2(new_n258), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT90), .Z(new_n806));
  INV_X1    g0606(.A(G143), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n806), .B1(new_n807), .B2(new_n707), .C1(new_n393), .C2(new_n725), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT34), .ZN(new_n809));
  INV_X1    g0609(.A(G132), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n719), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n728), .A2(new_n322), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n811), .B(new_n812), .C1(G50), .C2(new_n735), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n809), .A2(new_n271), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n730), .A2(new_n214), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n803), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n752), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n752), .A2(new_n695), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n203), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n791), .A2(new_n692), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n789), .A2(new_n790), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n790), .B1(new_n789), .B2(new_n820), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G384));
  INV_X1    g0625(.A(KEYINPUT100), .ZN(new_n826));
  XOR2_X1   g0626(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n636), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n418), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n421), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n421), .A2(KEYINPUT97), .A3(new_n830), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n831), .A2(new_n412), .B1(new_n832), .B2(KEYINPUT37), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n421), .A2(new_n830), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  NOR4_X1   g0635(.A1(new_n834), .A2(KEYINPUT97), .A3(new_n835), .A4(new_n413), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n830), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n426), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n828), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n830), .B1(new_n417), .B2(new_n425), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n421), .A2(new_n412), .A3(new_n830), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n835), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n421), .A2(new_n830), .A3(KEYINPUT37), .A4(new_n412), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n841), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n826), .B1(new_n840), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n342), .A2(new_n638), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n343), .A2(new_n347), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT95), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n319), .A2(new_n342), .A3(new_n638), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n851), .B1(new_n850), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n780), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT98), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n683), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n681), .A2(KEYINPUT98), .A3(new_n682), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n669), .A2(new_n859), .A3(new_n684), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT99), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT99), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n669), .A2(new_n859), .A3(new_n862), .A4(new_n684), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n855), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n832), .A2(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n842), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n831), .A2(KEYINPUT37), .A3(new_n832), .A4(new_n412), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n827), .B1(new_n868), .B2(new_n841), .ZN(new_n869));
  INV_X1    g0669(.A(new_n845), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n839), .A2(new_n870), .A3(KEYINPUT38), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(KEYINPUT100), .A3(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n848), .A2(KEYINPUT40), .A3(new_n864), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n861), .A2(new_n863), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n846), .B1(new_n841), .B2(new_n845), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n855), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n873), .A2(new_n880), .A3(new_n429), .A4(new_n874), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n873), .A2(new_n880), .A3(G330), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n429), .A2(new_n874), .A3(G330), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n881), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT39), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n840), .B2(new_n847), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n871), .A2(KEYINPUT39), .A3(new_n875), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n343), .A2(new_n638), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n375), .A2(new_n638), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n667), .B2(new_n778), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n853), .A2(new_n854), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n876), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n899), .A2(new_n900), .B1(new_n425), .B2(new_n829), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n893), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n886), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n668), .A2(new_n429), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n612), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n903), .B(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n207), .B2(new_n632), .ZN(new_n907));
  OAI211_X1 g0707(.A(G20), .B(new_n467), .C1(new_n520), .C2(KEYINPUT35), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n578), .B(new_n908), .C1(KEYINPUT35), .C2(new_n520), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT36), .Z(new_n910));
  NAND2_X1  g0710(.A1(new_n382), .A2(G77), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n230), .A2(new_n911), .B1(G50), .B2(new_n322), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(G1), .A3(new_n224), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n907), .A2(new_n910), .A3(new_n913), .ZN(G367));
  NOR2_X1   g0714(.A1(new_n730), .A2(new_n322), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n271), .B1(new_n707), .B2(new_n258), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n915), .B(new_n916), .C1(G50), .C2(new_n726), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n743), .A2(G137), .ZN(new_n918));
  INV_X1    g0718(.A(new_n728), .ZN(new_n919));
  AOI22_X1  g0719(.A1(G159), .A2(new_n793), .B1(new_n919), .B2(G77), .ZN(new_n920));
  AOI22_X1  g0720(.A1(G143), .A2(new_n723), .B1(new_n735), .B2(G58), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n917), .A2(new_n918), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n708), .A2(G303), .B1(G311), .B2(new_n723), .ZN(new_n923));
  INV_X1    g0723(.A(G317), .ZN(new_n924));
  OAI221_X1 g0724(.A(new_n360), .B1(new_n719), .B2(new_n924), .C1(new_n524), .C2(new_n728), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT106), .ZN(new_n926));
  AOI22_X1  g0726(.A1(G294), .A2(new_n793), .B1(new_n726), .B2(new_n794), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n741), .A2(G107), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n923), .A2(new_n926), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n716), .A2(new_n578), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT46), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n922), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT107), .Z(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT47), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n752), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n541), .A2(new_n558), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n638), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n620), .A2(new_n559), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n620), .B2(new_n937), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n939), .A2(new_n698), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n762), .B1(new_n540), .B2(new_n226), .C1(new_n241), .C2(new_n755), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n935), .A2(new_n692), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n652), .B(KEYINPUT41), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n650), .B1(new_n642), .B2(new_n649), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(new_n646), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n688), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n531), .A2(new_n563), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n622), .A2(new_n638), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n509), .A2(new_n622), .A3(new_n638), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n650), .A2(new_n648), .A3(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT45), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n650), .A2(new_n648), .ZN(new_n957));
  INV_X1    g0757(.A(new_n952), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n957), .A2(KEYINPUT44), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(KEYINPUT44), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n955), .A2(new_n956), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n647), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(KEYINPUT105), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT105), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n647), .A2(new_n964), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n961), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n961), .A2(new_n964), .A3(new_n647), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n947), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n688), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n944), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n690), .A2(G1), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n650), .A2(KEYINPUT102), .A3(new_n950), .ZN(new_n974));
  OAI21_X1  g0774(.A(KEYINPUT102), .B1(new_n650), .B2(new_n950), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT103), .ZN(new_n977));
  OR3_X1    g0777(.A1(new_n976), .A2(new_n977), .A3(KEYINPUT42), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(KEYINPUT42), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n952), .B(KEYINPUT101), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(new_n490), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n641), .B1(new_n981), .B2(new_n661), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n977), .B1(new_n976), .B2(KEYINPUT42), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n978), .A2(new_n979), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n962), .A2(new_n980), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT104), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n987), .B(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n986), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n984), .A2(new_n990), .A3(new_n985), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n943), .B1(new_n973), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(G387));
  INV_X1    g0797(.A(new_n946), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n969), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n999), .A2(new_n652), .A3(new_n947), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n642), .A2(new_n698), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(G311), .A2(new_n793), .B1(new_n726), .B2(G303), .ZN(new_n1002));
  INV_X1    g0802(.A(G322), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1002), .B1(new_n1003), .B2(new_n722), .C1(new_n707), .C2(new_n924), .ZN(new_n1004));
  XOR2_X1   g0804(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n735), .A2(G294), .B1(new_n741), .B2(new_n794), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT49), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n271), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n743), .A2(G326), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1006), .A2(KEYINPUT49), .A3(new_n1007), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n919), .A2(G116), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n722), .A2(new_n393), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n253), .A2(new_n793), .B1(new_n726), .B2(G68), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT109), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G97), .B2(new_n919), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n735), .A2(G77), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(KEYINPUT108), .B(G150), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n271), .B1(new_n719), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n540), .A2(new_n730), .ZN(new_n1022));
  AOI211_X1 g0822(.A(new_n1021), .B(new_n1022), .C1(G50), .C2(new_n708), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1018), .A2(new_n1019), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1014), .B1(new_n1015), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n752), .ZN(new_n1026));
  AOI21_X1  g0826(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n253), .A2(new_n202), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n655), .B(new_n1027), .C1(new_n1028), .C2(KEYINPUT50), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(KEYINPUT50), .B2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n754), .B1(new_n238), .B2(new_n457), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n759), .A2(new_n654), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n226), .A2(G107), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n762), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1001), .A2(new_n692), .A3(new_n1026), .A4(new_n1035), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1000), .B(new_n1036), .C1(new_n972), .C2(new_n998), .ZN(G393));
  OAI22_X1  g0837(.A1(new_n254), .A2(new_n725), .B1(new_n807), .B2(new_n719), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n707), .A2(new_n393), .B1(new_n258), .B2(new_n722), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT51), .Z(new_n1040));
  AOI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(G77), .C2(new_n741), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n793), .A2(G50), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n360), .B1(new_n919), .B2(G87), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n735), .A2(G68), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n707), .A2(new_n800), .B1(new_n924), .B2(new_n722), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT52), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n793), .A2(G303), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n271), .B1(new_n741), .B2(G116), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n725), .A2(new_n731), .B1(new_n719), .B2(new_n1003), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n738), .B(new_n1050), .C1(new_n735), .C2(new_n794), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n231), .B(new_n751), .C1(new_n1045), .C2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n692), .B1(new_n980), .B2(new_n698), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n249), .A2(new_n754), .B1(G97), .B2(new_n225), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1053), .B(new_n1054), .C1(new_n762), .C2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n966), .A2(new_n967), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1056), .B1(new_n1057), .B2(new_n971), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n966), .A2(new_n947), .A3(new_n967), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n652), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1058), .B1(new_n1060), .B2(new_n968), .ZN(G390));
  NAND3_X1  g0861(.A1(new_n874), .A2(G330), .A3(new_n877), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(KEYINPUT111), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT111), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n864), .A2(new_n1064), .A3(G330), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n897), .B1(new_n686), .B2(new_n778), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n896), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n686), .A2(new_n897), .A3(new_n778), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n874), .A2(G330), .A3(new_n780), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n897), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n895), .B1(new_n778), .B2(new_n664), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1068), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n612), .A2(new_n884), .A3(new_n904), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n899), .A2(new_n892), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n890), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n891), .B1(new_n1072), .B2(new_n898), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n848), .A3(new_n872), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1082), .A3(new_n1069), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n872), .ZN(new_n1084));
  AOI21_X1  g0884(.A(KEYINPUT100), .B1(new_n869), .B2(new_n871), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1086), .A2(new_n1081), .B1(new_n890), .B2(new_n1079), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1083), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1078), .A2(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1067), .A2(new_n896), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1092), .A2(new_n1076), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(new_n1089), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n1091), .A2(new_n1094), .A3(new_n653), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n691), .B1(new_n818), .B2(new_n254), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT112), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n707), .A2(new_n578), .B1(new_n524), .B2(new_n725), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n812), .B(new_n1098), .C1(G294), .C2(new_n743), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n793), .A2(G107), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n360), .B1(new_n716), .B2(new_n799), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT115), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n723), .A2(G283), .B1(new_n741), .B2(G77), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  XOR2_X1   g0904(.A(KEYINPUT54), .B(G143), .Z(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n1106), .A2(new_n725), .B1(new_n804), .B2(new_n713), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G159), .B2(new_n741), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT113), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n728), .A2(new_n202), .ZN(new_n1110));
  INV_X1    g0910(.A(G125), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n719), .A2(new_n1111), .ZN(new_n1112));
  NOR4_X1   g0912(.A1(new_n1109), .A2(new_n360), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n723), .A2(G128), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(new_n810), .C2(new_n707), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n716), .A2(new_n1020), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1104), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT116), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n1120), .A2(new_n231), .A3(new_n751), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1097), .B(new_n1121), .C1(new_n890), .C2(new_n695), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n1089), .B2(new_n971), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT117), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1095), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(G378));
  AND3_X1   g0926(.A1(new_n295), .A2(new_n269), .A3(new_n829), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n295), .B1(new_n269), .B2(new_n829), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OR3_X1    g0930(.A1(new_n1127), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n882), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1133), .A2(new_n873), .A3(new_n880), .A4(G330), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1135), .A2(new_n902), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n902), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT57), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1076), .B1(new_n1075), .B2(new_n1089), .ZN(new_n1141));
  NOR3_X1   g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(KEYINPUT119), .B1(new_n1142), .B2(new_n653), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1140), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1138), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1135), .A2(new_n902), .A3(new_n1136), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1141), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(new_n1148), .A3(KEYINPUT57), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT119), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1149), .A2(new_n1150), .A3(new_n652), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1143), .A2(new_n1144), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1147), .A2(new_n971), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n573), .A2(new_n726), .B1(G97), .B2(new_n793), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n214), .B2(new_n728), .C1(new_n729), .C2(new_n719), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n915), .B(new_n1155), .C1(G116), .C2(new_n723), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n708), .A2(G107), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n271), .A2(G41), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1156), .A2(new_n1019), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT58), .Z(new_n1160));
  OAI21_X1  g0960(.A(new_n202), .B1(new_n300), .B2(G41), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n708), .A2(G128), .B1(new_n735), .B2(new_n1105), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n722), .A2(new_n1111), .B1(new_n713), .B2(new_n810), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(G150), .B2(new_n741), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1162), .B(new_n1164), .C1(new_n804), .C2(new_n725), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n1165), .A2(KEYINPUT59), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n919), .A2(G159), .ZN(new_n1167));
  AOI21_X1  g0967(.A(G41), .B1(new_n743), .B2(G124), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1166), .A2(new_n255), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  AND2_X1   g0969(.A1(new_n1165), .A2(KEYINPUT59), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1161), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n752), .B1(new_n1160), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n818), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n692), .B1(G50), .B2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT118), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1172), .B(new_n1175), .C1(new_n1133), .C2(new_n696), .ZN(new_n1176));
  AND2_X1   g0976(.A1(new_n1153), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1152), .A2(new_n1177), .ZN(G375));
  OAI21_X1  g0978(.A(new_n692), .B1(G68), .B2(new_n1173), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1022), .B1(new_n708), .B2(G283), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n203), .B2(new_n728), .C1(new_n717), .C2(new_n719), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n722), .A2(new_n731), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n716), .A2(new_n524), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(new_n1181), .A2(new_n271), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n477), .B2(new_n725), .C1(new_n578), .C2(new_n713), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT121), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n707), .A2(new_n804), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n271), .B1(new_n730), .B2(new_n202), .C1(new_n393), .C2(new_n716), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1106), .A2(new_n713), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n728), .A2(new_n214), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n722), .A2(new_n810), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n743), .A2(G128), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n258), .C2(new_n725), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1186), .B1(new_n1187), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1179), .B1(new_n1195), .B2(new_n752), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n897), .A2(new_n695), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT120), .Z(new_n1198));
  AOI22_X1  g0998(.A1(new_n1075), .A2(new_n971), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1068), .A2(new_n1076), .A3(new_n1074), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n944), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1199), .B1(new_n1201), .B2(new_n1093), .ZN(G381));
  INV_X1    g1002(.A(KEYINPUT122), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(G375), .B(new_n1203), .ZN(new_n1204));
  OR2_X1    g1004(.A1(G381), .A2(G384), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(new_n1125), .A3(new_n1206), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(G387), .A2(G396), .A3(G393), .A4(G390), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1207), .A2(new_n1209), .ZN(G407));
  NAND2_X1  g1010(.A1(new_n637), .A2(G213), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT123), .Z(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1204), .A2(new_n1125), .A3(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(G213), .B(new_n1214), .C1(new_n1207), .C2(new_n1209), .ZN(G409));
  INV_X1    g1015(.A(KEYINPUT127), .ZN(new_n1216));
  INV_X1    g1016(.A(G390), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n996), .B2(new_n1217), .ZN(new_n1218));
  XNOR2_X1  g1018(.A(G393), .B(G396), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n994), .B1(new_n970), .B2(new_n972), .ZN(new_n1220));
  OAI21_X1  g1020(.A(G390), .B1(new_n1220), .B2(new_n943), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1219), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1152), .A2(G378), .A3(new_n1177), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1147), .A2(new_n1148), .A3(new_n944), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1139), .B(KEYINPUT124), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1226), .B(new_n1176), .C1(new_n1227), .C2(new_n972), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n1125), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1225), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT60), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1200), .A2(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1068), .A2(KEYINPUT60), .A3(new_n1074), .A4(new_n1076), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1232), .A2(new_n1078), .A3(new_n652), .A4(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(KEYINPUT125), .B(new_n824), .C1(new_n1234), .C2(new_n1199), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT125), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n822), .B2(new_n823), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n823), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(KEYINPUT125), .A3(new_n821), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1234), .A2(new_n1199), .A3(new_n1237), .A4(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1235), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1230), .A2(new_n1211), .A3(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT62), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1213), .B1(new_n1225), .B2(new_n1229), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1244), .A2(new_n1245), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT61), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1233), .B(new_n652), .C1(new_n1076), .C2(new_n1092), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT60), .B1(new_n1092), .B2(new_n1076), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1239), .B(new_n1199), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1237), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1213), .A2(G2897), .ZN(new_n1255));
  AND3_X1   g1055(.A1(new_n1254), .A2(new_n1240), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n637), .A2(G213), .A3(G2897), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(new_n1254), .B2(new_n1240), .ZN(new_n1258));
  OAI21_X1  g1058(.A(KEYINPUT126), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1257), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n1235), .B2(new_n1241), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT126), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1254), .A2(new_n1240), .A3(new_n1255), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1259), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1249), .B1(new_n1246), .B2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1224), .B1(new_n1248), .B2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1242), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1224), .B1(new_n1246), .B2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1230), .A2(new_n1211), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1256), .A2(new_n1258), .A3(KEYINPUT126), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1262), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1268), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1244), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1249), .B(new_n1270), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1267), .A2(new_n1277), .ZN(G405));
  OR3_X1    g1078(.A1(new_n1222), .A2(new_n1223), .A3(new_n1242), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1242), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(G375), .B(G378), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1281), .B(new_n1282), .ZN(G402));
endmodule


