//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT64), .A2(G143), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT64), .A2(G143), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G146), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT64), .A2(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT64), .A2(G143), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n191), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n191), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n202));
  AOI22_X1  g016(.A1(new_n198), .A2(new_n200), .B1(G128), .B2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT67), .B1(new_n195), .B2(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n188), .A2(new_n189), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n199), .B1(new_n207), .B2(new_n191), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n193), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n205), .B(new_n206), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(G134), .B(G137), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT65), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(G134), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(G137), .ZN(new_n216));
  INV_X1    g030(.A(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(KEYINPUT11), .A3(G134), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(G137), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n216), .A2(new_n218), .A3(new_n212), .A4(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n215), .A2(G137), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n217), .A2(G134), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n221), .B(G131), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n213), .A2(new_n220), .A3(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n204), .A2(new_n210), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT68), .ZN(new_n227));
  AND2_X1   g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n190), .A2(new_n192), .A3(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT0), .B(G128), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(new_n198), .B2(new_n200), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT66), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G131), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n220), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n229), .B(new_n237), .C1(new_n208), .C2(new_n231), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n233), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n204), .A2(new_n240), .A3(new_n210), .A4(new_n225), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n227), .A2(KEYINPUT30), .A3(new_n239), .A4(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n239), .A2(KEYINPUT30), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n245), .A2(KEYINPUT69), .A3(new_n227), .A4(new_n241), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n225), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n229), .B1(new_n208), .B2(new_n231), .ZN(new_n250));
  INV_X1    g064(.A(new_n236), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT30), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(G116), .B(G119), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT2), .B(G113), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n247), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n227), .A2(new_n257), .A3(new_n239), .A4(new_n241), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G101), .ZN(new_n263));
  INV_X1    g077(.A(G237), .ZN(new_n264));
  INV_X1    g078(.A(G953), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(new_n265), .A3(G210), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n263), .B(new_n266), .ZN(new_n267));
  XNOR2_X1  g081(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n261), .A2(KEYINPUT31), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n259), .B1(new_n244), .B2(new_n246), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n273), .B1(new_n274), .B2(new_n270), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n252), .A2(new_n258), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n262), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT28), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n239), .A2(new_n226), .A3(new_n257), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT28), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n269), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT71), .B1(new_n276), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n286), .B(new_n283), .C1(new_n272), .C2(new_n275), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n187), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT72), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(KEYINPUT72), .B(new_n187), .C1(new_n285), .C2(new_n287), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT73), .B(KEYINPUT32), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n261), .A2(new_n262), .ZN(new_n294));
  INV_X1    g108(.A(new_n269), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n282), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n297), .B1(new_n278), .B2(KEYINPUT28), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT29), .B1(new_n298), .B2(new_n269), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT74), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n227), .A2(new_n239), .A3(new_n241), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n258), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n262), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n297), .B1(new_n304), .B2(KEYINPUT28), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n269), .A2(KEYINPUT29), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n300), .A2(KEYINPUT74), .ZN(new_n309));
  OAI21_X1  g123(.A(G472), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT31), .B1(new_n261), .B2(new_n271), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n274), .A2(new_n273), .A3(new_n270), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n284), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n286), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n276), .A2(KEYINPUT71), .A3(new_n284), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(KEYINPUT32), .A3(new_n187), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT75), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n316), .A2(new_n319), .A3(KEYINPUT32), .A4(new_n187), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n293), .A2(new_n310), .A3(new_n318), .A4(new_n320), .ZN(new_n321));
  XOR2_X1   g135(.A(KEYINPUT76), .B(G217), .Z(new_n322));
  INV_X1    g136(.A(G902), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(G234), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G125), .B(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT16), .ZN(new_n326));
  INV_X1    g140(.A(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G125), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(KEYINPUT16), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(new_n191), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n331));
  INV_X1    g145(.A(G119), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(G128), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n333), .B(new_n334), .C1(G119), .C2(new_n193), .ZN(new_n335));
  XNOR2_X1  g149(.A(G119), .B(G128), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT24), .B(G110), .Z(new_n337));
  AOI22_X1  g151(.A1(new_n335), .A2(G110), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n330), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n325), .A2(new_n191), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n340), .B(KEYINPUT77), .Z(new_n341));
  OR2_X1    g155(.A1(new_n329), .A2(new_n191), .ZN(new_n342));
  OAI22_X1  g156(.A1(new_n335), .A2(G110), .B1(new_n336), .B2(new_n337), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT78), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n339), .A2(new_n347), .A3(new_n344), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n265), .A2(G221), .A3(G234), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n349), .B(new_n350), .Z(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n346), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n345), .A2(KEYINPUT78), .A3(new_n351), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT25), .B1(new_n355), .B2(new_n323), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT25), .ZN(new_n357));
  AOI211_X1 g171(.A(new_n357), .B(G902), .C1(new_n353), .C2(new_n354), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n324), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n324), .A2(G902), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G104), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(G107), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n363), .A2(G107), .ZN(new_n367));
  XOR2_X1   g181(.A(KEYINPUT80), .B(G107), .Z(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(new_n363), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n366), .B1(new_n369), .B2(new_n365), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT81), .B(G101), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n364), .ZN(new_n374));
  XNOR2_X1  g188(.A(KEYINPUT80), .B(G107), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n374), .B1(new_n375), .B2(G104), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G101), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n378));
  INV_X1    g192(.A(G116), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n379), .A2(KEYINPUT5), .A3(G119), .ZN(new_n380));
  INV_X1    g194(.A(G113), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n256), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n378), .A2(new_n382), .B1(new_n383), .B2(new_n255), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n373), .A2(new_n377), .A3(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(KEYINPUT86), .ZN(new_n386));
  INV_X1    g200(.A(new_n366), .ZN(new_n387));
  INV_X1    g201(.A(new_n367), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n388), .B1(new_n375), .B2(G104), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n387), .B1(new_n389), .B2(KEYINPUT3), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT4), .A3(G101), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n392), .B1(new_n370), .B2(new_n372), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n390), .A2(G101), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n395), .A2(KEYINPUT85), .A3(new_n258), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT85), .B1(new_n395), .B2(new_n258), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n386), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G110), .B(G122), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n399), .B(new_n386), .C1(new_n396), .C2(new_n397), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(KEYINPUT6), .A3(new_n402), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n248), .A2(G125), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n250), .A2(G125), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G224), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(G953), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n406), .B(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n398), .A2(new_n410), .A3(new_n400), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n403), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT7), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n406), .B1(new_n413), .B2(new_n408), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n406), .A2(new_n408), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n414), .B1(new_n415), .B2(new_n413), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n370), .A2(new_n372), .B1(G101), .B2(new_n376), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(new_n384), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n399), .B(KEYINPUT8), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n416), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(G902), .B1(new_n420), .B2(new_n402), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n412), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G210), .B1(G237), .B2(G902), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n412), .A2(new_n423), .A3(new_n421), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G221), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT9), .B(G234), .Z(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT79), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n428), .B1(new_n430), .B2(new_n323), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n265), .A2(G952), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(G234), .B2(G237), .ZN(new_n434));
  AOI211_X1 g248(.A(new_n323), .B(new_n265), .C1(G234), .C2(G237), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(G898), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G214), .B1(G237), .B2(G902), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT84), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n233), .A2(new_n238), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n395), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n190), .A2(new_n192), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n193), .B1(new_n198), .B2(KEYINPUT1), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n205), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n373), .A2(new_n377), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT10), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n417), .A2(KEYINPUT10), .A3(new_n204), .A4(new_n210), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n442), .A2(new_n251), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G140), .ZN(new_n451));
  INV_X1    g265(.A(G227), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G953), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n451), .B(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT83), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT83), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n450), .A2(new_n458), .A3(new_n455), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n446), .B1(new_n417), .B2(new_n248), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n460), .A2(KEYINPUT12), .A3(new_n236), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT12), .B1(new_n460), .B2(new_n236), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n457), .A2(new_n459), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n442), .A2(new_n448), .A3(new_n449), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n236), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n450), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n454), .ZN(new_n468));
  AOI211_X1 g282(.A(G469), .B(G902), .C1(new_n464), .C2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n461), .A2(new_n462), .ZN(new_n470));
  INV_X1    g284(.A(new_n450), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n454), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n456), .A2(KEYINPUT82), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n466), .B1(new_n456), .B2(KEYINPUT82), .ZN(new_n474));
  OAI211_X1 g288(.A(G469), .B(new_n472), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(G469), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n476), .A2(new_n323), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n432), .B(new_n440), .C1(new_n469), .C2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G122), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G116), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT95), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n379), .A2(G122), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(KEYINPUT14), .ZN(new_n487));
  OAI21_X1  g301(.A(G107), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(new_n486), .A3(new_n375), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n196), .A2(new_n197), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G128), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n193), .A2(G143), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n215), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n215), .B1(new_n492), .B2(new_n493), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n495), .A2(KEYINPUT96), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT96), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n492), .A2(new_n493), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(G134), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n499), .B1(new_n501), .B2(new_n496), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n490), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n489), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n375), .B1(new_n484), .B2(new_n486), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n495), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G134), .B1(new_n492), .B2(KEYINPUT13), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n494), .B2(KEYINPUT13), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n322), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n430), .A2(new_n265), .A3(new_n510), .ZN(new_n511));
  OR3_X1    g325(.A1(new_n503), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n503), .B2(new_n509), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT97), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  OAI211_X1 g329(.A(KEYINPUT97), .B(new_n511), .C1(new_n503), .C2(new_n509), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n515), .A2(KEYINPUT98), .A3(new_n323), .A4(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G478), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n517), .A2(new_n519), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n264), .A2(new_n265), .A3(G214), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(new_n201), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n491), .A2(new_n524), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n523), .B1(new_n527), .B2(G131), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(G131), .B2(new_n527), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n525), .A2(new_n526), .A3(new_n523), .A4(new_n212), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT17), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n329), .A2(new_n191), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n527), .A2(KEYINPUT17), .A3(G131), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n342), .A2(new_n533), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n535), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT93), .B1(new_n330), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n532), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n325), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G146), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n341), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(KEYINPUT18), .A2(G131), .ZN(new_n543));
  XOR2_X1   g357(.A(new_n527), .B(new_n543), .Z(new_n544));
  NOR2_X1   g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n539), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(G113), .B(G122), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT92), .B(G104), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n548), .B(new_n549), .Z(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(KEYINPUT94), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n550), .B1(new_n539), .B2(new_n546), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n538), .A2(new_n536), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n546), .B(new_n550), .C1(new_n554), .C2(new_n531), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT94), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n552), .B(new_n323), .C1(new_n553), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G475), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT89), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n529), .B2(new_n530), .ZN(new_n561));
  XOR2_X1   g375(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n325), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(KEYINPUT91), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n563), .A2(KEYINPUT91), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n540), .A2(KEYINPUT19), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n342), .B1(new_n567), .B2(G146), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n561), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n529), .A2(new_n560), .A3(new_n530), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n545), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n555), .B1(new_n571), .B2(new_n550), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT20), .ZN(new_n573));
  NOR2_X1   g387(.A1(G475), .A2(G902), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n574), .ZN(new_n576));
  INV_X1    g390(.A(new_n570), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n577), .A2(new_n561), .A3(new_n568), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n551), .B1(new_n578), .B2(new_n545), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n576), .B1(new_n579), .B2(new_n555), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n575), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n559), .A2(new_n582), .ZN(new_n583));
  NOR4_X1   g397(.A1(new_n427), .A2(new_n480), .A3(new_n522), .A4(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n321), .A2(new_n362), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(new_n371), .ZN(G3));
  OAI21_X1  g400(.A(new_n323), .B1(new_n285), .B2(new_n287), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G472), .ZN(new_n588));
  AND4_X1   g402(.A1(new_n290), .A2(new_n588), .A3(new_n291), .A4(new_n362), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n515), .A2(new_n323), .A3(new_n516), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT100), .B(G478), .Z(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT33), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n515), .A2(new_n593), .A3(new_n516), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT33), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n594), .A2(G478), .A3(new_n323), .A4(new_n595), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n559), .A2(new_n582), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n437), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n425), .A2(KEYINPUT99), .A3(new_n426), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n423), .B1(new_n412), .B2(new_n421), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n439), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n599), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n475), .A2(new_n478), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n464), .A2(new_n468), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n476), .A3(new_n323), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n431), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n589), .A2(new_n604), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT34), .B(G104), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  INV_X1    g425(.A(new_n581), .ZN(new_n612));
  INV_X1    g426(.A(new_n572), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(new_n576), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n580), .A2(new_n581), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n614), .A2(new_n615), .B1(new_n558), .B2(G475), .ZN(new_n616));
  INV_X1    g430(.A(new_n437), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n522), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT101), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n616), .A2(new_n620), .A3(new_n522), .A4(new_n617), .ZN(new_n621));
  AND4_X1   g435(.A1(new_n600), .A2(new_n619), .A3(new_n603), .A4(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(new_n589), .A3(new_n608), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(G107), .Z(new_n624));
  XOR2_X1   g438(.A(KEYINPUT102), .B(KEYINPUT35), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  AND3_X1   g440(.A1(new_n290), .A2(new_n588), .A3(new_n291), .ZN(new_n627));
  INV_X1    g441(.A(new_n324), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n348), .A2(new_n352), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n347), .B1(new_n339), .B2(new_n344), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n354), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n323), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n357), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n355), .A2(KEYINPUT25), .A3(new_n323), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n628), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n352), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n345), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n360), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT103), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n614), .A2(new_n575), .B1(new_n558), .B2(G475), .ZN(new_n642));
  INV_X1    g456(.A(new_n521), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n517), .A2(new_n519), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n359), .A2(new_n646), .A3(new_n639), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n641), .A2(new_n642), .A3(new_n645), .A4(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n427), .A2(new_n480), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n627), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  AND2_X1   g466(.A1(new_n641), .A2(new_n647), .ZN(new_n653));
  INV_X1    g467(.A(G900), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n434), .B1(new_n435), .B2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n653), .A2(new_n616), .A3(new_n656), .ZN(new_n657));
  AND4_X1   g471(.A1(new_n522), .A2(new_n600), .A3(new_n608), .A4(new_n603), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n321), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  OR2_X1    g474(.A1(new_n427), .A2(KEYINPUT38), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n427), .A2(KEYINPUT38), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n359), .A2(new_n639), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n439), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n665), .A2(new_n522), .A3(new_n583), .A4(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n655), .B(KEYINPUT39), .Z(new_n669));
  NAND2_X1  g483(.A1(new_n608), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT40), .Z(new_n671));
  INV_X1    g485(.A(new_n294), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n295), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n323), .B1(new_n304), .B2(new_n269), .ZN(new_n674));
  OAI21_X1  g488(.A(G472), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n293), .A2(new_n318), .A3(new_n320), .A4(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n668), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(new_n207), .ZN(G45));
  AND2_X1   g492(.A1(new_n600), .A2(new_n603), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n598), .A2(new_n655), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n680), .A2(new_n608), .A3(new_n653), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n321), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  NAND2_X1  g497(.A1(new_n606), .A2(new_n323), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G469), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n685), .A2(new_n432), .A3(new_n607), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n321), .A2(new_n362), .A3(new_n604), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NAND4_X1  g503(.A1(new_n321), .A2(new_n362), .A3(new_n622), .A4(new_n686), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  NAND2_X1  g505(.A1(new_n686), .A2(new_n617), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n648), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n321), .A2(new_n693), .A3(new_n679), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G119), .ZN(G21));
  OAI22_X1  g509(.A1(new_n311), .A2(new_n312), .B1(new_n269), .B2(new_n305), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n187), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n587), .B2(G472), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n362), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n600), .A2(new_n603), .A3(new_n522), .A4(new_n583), .ZN(new_n701));
  OR3_X1    g515(.A1(new_n700), .A2(new_n701), .A3(new_n692), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G122), .ZN(G24));
  AND3_X1   g517(.A1(new_n686), .A2(new_n600), .A3(new_n603), .ZN(new_n704));
  AOI21_X1  g518(.A(G902), .B1(new_n314), .B2(new_n315), .ZN(new_n705));
  INV_X1    g519(.A(G472), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n664), .B(new_n697), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(KEYINPUT104), .B1(new_n699), .B2(new_n664), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n680), .B(new_n704), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  NAND3_X1  g526(.A1(new_n427), .A2(new_n608), .A3(new_n666), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n321), .A2(new_n362), .A3(new_n680), .A4(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT32), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n288), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n310), .A2(new_n718), .A3(new_n317), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n362), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n680), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n713), .A2(new_n722), .A3(new_n716), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n715), .A2(new_n716), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n212), .ZN(G33));
  AND3_X1   g539(.A1(new_n616), .A2(new_n522), .A3(new_n656), .ZN(new_n726));
  AND4_X1   g540(.A1(new_n321), .A2(new_n362), .A3(new_n714), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n215), .ZN(G36));
  NAND2_X1  g542(.A1(new_n427), .A2(new_n666), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n642), .A2(KEYINPUT105), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n583), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n596), .A2(new_n592), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n583), .A2(KEYINPUT43), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n734), .A2(KEYINPUT43), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n290), .A2(new_n588), .A3(new_n291), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n737), .A2(KEYINPUT106), .A3(new_n664), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT106), .B1(new_n737), .B2(new_n664), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n729), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n743));
  OAI211_X1 g557(.A(KEYINPUT44), .B(new_n736), .C1(new_n738), .C2(new_n739), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n476), .B1(new_n746), .B2(new_n747), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n477), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n750), .A2(KEYINPUT46), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n607), .B1(new_n750), .B2(KEYINPUT46), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n432), .B(new_n669), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n745), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n743), .B1(new_n742), .B2(new_n744), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G137), .ZN(G39));
  OAI21_X1  g572(.A(new_n432), .B1(new_n751), .B2(new_n752), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(KEYINPUT108), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(KEYINPUT108), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI221_X1 g577(.A(new_n432), .B1(KEYINPUT108), .B2(new_n760), .C1(new_n751), .C2(new_n752), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n729), .ZN(new_n766));
  INV_X1    g580(.A(new_n362), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n767), .A3(new_n680), .ZN(new_n768));
  OR3_X1    g582(.A1(new_n768), .A2(new_n321), .A3(KEYINPUT109), .ZN(new_n769));
  OAI21_X1  g583(.A(KEYINPUT109), .B1(new_n768), .B2(new_n321), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n765), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n327), .ZN(G42));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n608), .A2(new_n665), .A3(new_n656), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n701), .A2(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n676), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n773), .B1(new_n676), .B2(new_n775), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n659), .A2(new_n682), .A3(new_n711), .ZN(new_n779));
  OAI21_X1  g593(.A(KEYINPUT52), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n659), .A2(new_n682), .A3(new_n711), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n676), .A2(new_n775), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT112), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n676), .A2(new_n775), .A3(new_n773), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n781), .A2(new_n782), .A3(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n780), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n715), .A2(new_n716), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n721), .A2(new_n723), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n727), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n707), .A2(new_n708), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n699), .A2(KEYINPUT104), .A3(new_n664), .ZN(new_n793));
  AOI211_X1 g607(.A(new_n722), .B(new_n713), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n795), .B1(new_n643), .B2(new_n644), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n520), .A2(KEYINPUT110), .A3(new_n521), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n713), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n321), .A2(new_n799), .A3(new_n657), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT111), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n321), .A2(new_n799), .A3(new_n802), .A4(new_n657), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n794), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n791), .A2(new_n804), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n687), .A2(new_n690), .A3(new_n694), .A4(new_n702), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n597), .B1(new_n798), .B2(new_n642), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n807), .A2(new_n427), .A3(new_n480), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n589), .A2(new_n808), .B1(new_n627), .B2(new_n649), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n585), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n782), .B1(new_n659), .B2(new_n711), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n813), .A2(KEYINPUT53), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n788), .A2(new_n805), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT53), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n780), .A2(new_n787), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n791), .A2(new_n804), .A3(new_n806), .A4(new_n810), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT54), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n685), .A2(new_n607), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n763), .A2(new_n764), .B1(new_n431), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n736), .A2(new_n434), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n700), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n766), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n823), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n766), .A2(new_n686), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n826), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(new_n710), .B2(new_n709), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n686), .A2(new_n439), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(new_n661), .B2(new_n662), .ZN(new_n834));
  NOR2_X1   g648(.A1(KEYINPUT115), .A2(KEYINPUT50), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n827), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n434), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n830), .A2(new_n767), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n676), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n583), .A2(new_n733), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n827), .A2(new_n834), .ZN(new_n843));
  XOR2_X1   g657(.A(KEYINPUT115), .B(KEYINPUT50), .Z(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n829), .A2(new_n837), .A3(new_n842), .A4(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n825), .A2(new_n823), .A3(new_n828), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n822), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n837), .A2(KEYINPUT116), .A3(new_n842), .A4(new_n845), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n845), .A2(new_n842), .A3(new_n836), .A4(new_n832), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT116), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n825), .A2(new_n828), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n849), .A2(new_n852), .A3(KEYINPUT51), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n831), .A2(new_n721), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT48), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n839), .A2(new_n597), .A3(new_n840), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n433), .B(KEYINPUT117), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n827), .B2(new_n704), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n848), .A2(new_n854), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n585), .A2(new_n809), .A3(KEYINPUT53), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n813), .A2(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n863), .A2(new_n791), .A3(new_n804), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n687), .A2(new_n690), .A3(new_n694), .A4(new_n702), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT113), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n788), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n867), .A2(new_n819), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n821), .A2(new_n861), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT118), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n821), .A2(new_n861), .A3(new_n872), .A4(new_n869), .ZN(new_n873));
  OR2_X1    g687(.A1(G952), .A2(G953), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n824), .B(KEYINPUT49), .Z(new_n876));
  NAND3_X1  g690(.A1(new_n362), .A2(new_n432), .A3(new_n666), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n876), .A2(new_n734), .A3(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n878), .A2(new_n840), .A3(new_n663), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n875), .A2(new_n879), .ZN(G75));
  NOR2_X1   g694(.A1(new_n265), .A2(G952), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n867), .A2(new_n819), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(G210), .A3(G902), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT56), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n403), .A2(new_n411), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n409), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT55), .Z(new_n888));
  AOI21_X1  g702(.A(new_n881), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n888), .B(KEYINPUT119), .Z(new_n890));
  NAND3_X1  g704(.A1(new_n883), .A2(new_n884), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT120), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n883), .A2(KEYINPUT120), .A3(new_n884), .A4(new_n890), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n889), .A2(new_n893), .A3(new_n894), .ZN(G51));
  XOR2_X1   g709(.A(new_n606), .B(KEYINPUT121), .Z(new_n896));
  XNOR2_X1  g710(.A(new_n882), .B(new_n868), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n477), .B(KEYINPUT57), .Z(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n323), .B1(new_n867), .B2(new_n819), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n748), .A3(new_n749), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n881), .B1(new_n899), .B2(new_n901), .ZN(G54));
  AND2_X1   g716(.A1(KEYINPUT58), .A2(G475), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n900), .A2(new_n572), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n572), .B1(new_n900), .B2(new_n903), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n904), .A2(new_n905), .A3(new_n881), .ZN(G60));
  INV_X1    g720(.A(new_n881), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n594), .A2(new_n595), .ZN(new_n908));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT59), .Z(new_n910));
  OR2_X1    g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n907), .B1(new_n897), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n910), .B1(new_n821), .B2(new_n869), .ZN(new_n913));
  INV_X1    g727(.A(new_n908), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT60), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n882), .A2(new_n638), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n918), .B1(new_n867), .B2(new_n819), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n920), .B(new_n907), .C1(new_n355), .C2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n920), .A2(KEYINPUT122), .A3(new_n907), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(KEYINPUT61), .A3(new_n923), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n921), .A2(new_n355), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n881), .B1(new_n921), .B2(new_n638), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n927));
  OAI211_X1 g741(.A(new_n925), .B(new_n926), .C1(KEYINPUT122), .C2(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n924), .A2(new_n928), .ZN(G66));
  OAI21_X1  g743(.A(G953), .B1(new_n436), .B2(new_n407), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n812), .B2(G953), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n886), .B1(G898), .B2(new_n265), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT123), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G69));
  NAND2_X1  g748(.A1(new_n247), .A2(new_n254), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n567), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(G953), .ZN(new_n937));
  INV_X1    g751(.A(new_n807), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n938), .A2(new_n669), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(new_n321), .A3(new_n362), .A4(new_n714), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT124), .B1(new_n757), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n781), .A2(new_n677), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT62), .Z(new_n943));
  OAI211_X1 g757(.A(KEYINPUT124), .B(new_n940), .C1(new_n755), .C2(new_n756), .ZN(new_n944));
  INV_X1    g758(.A(new_n771), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n937), .B1(new_n941), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n265), .A2(G900), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n791), .A2(KEYINPUT125), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n724), .B2(new_n727), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NOR3_X1   g766(.A1(new_n753), .A2(new_n720), .A3(new_n701), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n771), .A2(new_n779), .A3(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n952), .B(new_n954), .C1(new_n755), .C2(new_n756), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n948), .B1(new_n955), .B2(new_n265), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n936), .B1(new_n956), .B2(KEYINPUT126), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n958));
  AOI211_X1 g772(.A(new_n958), .B(new_n948), .C1(new_n955), .C2(new_n265), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n947), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(G953), .B1(new_n452), .B2(new_n654), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT127), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n947), .B(new_n962), .C1(new_n957), .C2(new_n959), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(G72));
  NAND2_X1  g780(.A1(G472), .A2(G902), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT63), .Z(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(new_n955), .B2(new_n811), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n969), .A2(new_n295), .A3(new_n672), .ZN(new_n970));
  INV_X1    g784(.A(new_n968), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n261), .A2(new_n271), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n296), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n881), .B1(new_n820), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n941), .A2(new_n946), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n968), .B1(new_n976), .B2(new_n811), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n975), .B1(new_n977), .B2(new_n673), .ZN(G57));
endmodule


