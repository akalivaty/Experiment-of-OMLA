//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G146), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G143), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n188), .A2(G143), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n197), .B1(new_n190), .B2(G143), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n196), .B1(new_n198), .B2(new_n192), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n188), .A2(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n202), .A3(G143), .ZN(new_n203));
  INV_X1    g017(.A(new_n197), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n203), .A2(new_n196), .A3(new_n204), .A4(new_n192), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n195), .B1(new_n199), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G137), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT11), .A3(G134), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(G137), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G131), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n210), .A2(new_n212), .A3(new_n217), .A4(new_n213), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n214), .A2(KEYINPUT66), .A3(G131), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n187), .B1(new_n207), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n219), .A2(new_n220), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n203), .A2(new_n204), .A3(new_n192), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n225), .A2(new_n205), .B1(new_n191), .B2(new_n194), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(KEYINPUT67), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n203), .A2(new_n204), .A3(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n228), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n231));
  INV_X1    g045(.A(new_n189), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n200), .A2(new_n202), .ZN(new_n233));
  INV_X1    g047(.A(G143), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n230), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n213), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n209), .A2(G137), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n239), .A2(new_n218), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n222), .A2(new_n227), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT30), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT2), .A2(G113), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT68), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT2), .A3(G113), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT2), .ZN(new_n249));
  INV_X1    g063(.A(G113), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n246), .A2(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G116), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT70), .B1(new_n252), .B2(G119), .ZN(new_n253));
  AND2_X1   g067(.A1(KEYINPUT69), .A2(G116), .ZN(new_n254));
  NOR2_X1   g068(.A1(KEYINPUT69), .A2(G116), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n253), .B1(new_n256), .B2(G119), .ZN(new_n257));
  INV_X1    g071(.A(G119), .ZN(new_n258));
  NOR4_X1   g072(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT70), .A4(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n251), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  OR2_X1    g074(.A1(KEYINPUT69), .A2(G116), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT69), .A2(G116), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(G119), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n253), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n246), .A2(new_n248), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n249), .A2(new_n250), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n261), .A2(new_n269), .A3(G119), .A4(new_n262), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n260), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT71), .B1(new_n207), .B2(new_n221), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n226), .A2(new_n274), .A3(new_n220), .A4(new_n219), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n273), .A2(new_n275), .A3(KEYINPUT30), .A4(new_n241), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n244), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  NOR3_X1   g091(.A1(new_n257), .A2(new_n259), .A3(new_n251), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n268), .B1(new_n265), .B2(new_n270), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n241), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n273), .A3(new_n275), .ZN(new_n283));
  NOR2_X1   g097(.A1(G237), .A2(G953), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G210), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT27), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT26), .B(G101), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n277), .A2(new_n283), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT31), .ZN(new_n290));
  INV_X1    g104(.A(new_n288), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT28), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n242), .A2(new_n272), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(new_n283), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n223), .A2(new_n226), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT28), .B1(new_n282), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n291), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT31), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n277), .A2(new_n298), .A3(new_n283), .A4(new_n288), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n290), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(G472), .A2(G902), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n273), .A2(new_n241), .A3(new_n275), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n272), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n292), .B1(new_n305), .B2(new_n283), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n288), .A2(KEYINPUT29), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n306), .A2(new_n296), .A3(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n303), .B1(new_n308), .B2(G902), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n277), .A2(new_n283), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n291), .ZN(new_n311));
  INV_X1    g125(.A(new_n241), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n295), .B2(new_n187), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n280), .B1(new_n313), .B2(new_n227), .ZN(new_n314));
  INV_X1    g128(.A(new_n283), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT28), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n296), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(new_n288), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n311), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G902), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n273), .A2(new_n275), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n322), .A2(new_n282), .B1(new_n304), .B2(new_n272), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n317), .B1(new_n323), .B2(new_n292), .ZN(new_n324));
  OAI211_X1 g138(.A(KEYINPUT73), .B(new_n321), .C1(new_n324), .C2(new_n307), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n309), .A2(new_n320), .A3(new_n325), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n302), .A2(KEYINPUT32), .B1(new_n326), .B2(G472), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n300), .A2(new_n301), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT32), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(KEYINPUT72), .A3(new_n329), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n327), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G125), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT76), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n335), .A2(KEYINPUT76), .A3(G125), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT16), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT16), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n336), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n188), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(G125), .B(G140), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n190), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT24), .B(G110), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(KEYINPUT75), .ZN(new_n349));
  XNOR2_X1  g163(.A(G119), .B(G128), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n258), .B2(G128), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n228), .A2(KEYINPUT23), .A3(G119), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n353), .B(new_n354), .C1(G119), .C2(new_n228), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(G110), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n345), .B(new_n347), .C1(new_n351), .C2(new_n356), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n349), .A2(new_n350), .B1(G110), .B2(new_n355), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n341), .A2(new_n188), .A3(new_n343), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n358), .B1(new_n359), .B2(new_n344), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT22), .B(G137), .ZN(new_n362));
  INV_X1    g176(.A(G953), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(G221), .A3(G234), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n362), .B(new_n364), .ZN(new_n365));
  XOR2_X1   g179(.A(new_n365), .B(KEYINPUT77), .Z(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n357), .A2(new_n360), .A3(new_n365), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G217), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(G234), .B2(new_n321), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n373), .B(KEYINPUT74), .Z(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n321), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n369), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n368), .A2(new_n377), .A3(new_n321), .A4(new_n370), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT25), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n368), .A2(new_n321), .A3(new_n370), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n377), .B1(new_n381), .B2(KEYINPUT79), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n374), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n376), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(G214), .B1(G237), .B2(G902), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(G210), .B1(G237), .B2(G902), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT3), .B1(new_n392), .B2(G107), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n394));
  INV_X1    g208(.A(G107), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(new_n395), .A3(G104), .ZN(new_n396));
  INV_X1    g210(.A(G101), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(G107), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n393), .A2(new_n396), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n392), .A2(G107), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n395), .A2(G104), .ZN(new_n401));
  OAI21_X1  g215(.A(G101), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n260), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT84), .B(KEYINPUT5), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n252), .A2(G119), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G113), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n254), .A2(new_n255), .A3(new_n258), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n270), .B1(new_n410), .B2(new_n253), .ZN(new_n411));
  INV_X1    g225(.A(new_n406), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n405), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n393), .A2(new_n396), .A3(new_n398), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G101), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT4), .A3(new_n399), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT4), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n419), .A3(G101), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n415), .B1(new_n280), .B2(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n418), .A2(new_n420), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(KEYINPUT83), .A3(new_n272), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n414), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G110), .B(G122), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n391), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n280), .A2(new_n421), .A3(new_n415), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT83), .B1(new_n423), .B2(new_n272), .ZN(new_n429));
  OAI22_X1  g243(.A1(new_n428), .A2(new_n429), .B1(new_n405), .B2(new_n413), .ZN(new_n430));
  INV_X1    g244(.A(new_n426), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n226), .B2(new_n337), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n207), .A2(KEYINPUT85), .A3(G125), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n337), .B(new_n230), .C1(new_n231), .C2(new_n235), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n363), .A2(G224), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n430), .A2(new_n391), .A3(new_n431), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n433), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n409), .B1(new_n411), .B2(KEYINPUT5), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT86), .B1(new_n405), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT5), .B1(new_n257), .B2(new_n259), .ZN(new_n445));
  INV_X1    g259(.A(new_n409), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n403), .B1(new_n411), .B2(new_n251), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n403), .B1(new_n413), .B2(new_n279), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n444), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n426), .B(KEYINPUT8), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT7), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n439), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n435), .A2(new_n436), .A3(new_n437), .A4(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n437), .B1(new_n226), .B2(new_n337), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n458), .B1(new_n455), .B2(new_n439), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n454), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AOI211_X1 g274(.A(new_n431), .B(new_n414), .C1(new_n422), .C2(new_n424), .ZN(new_n461));
  OAI211_X1 g275(.A(KEYINPUT87), .B(new_n321), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n442), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n425), .A2(new_n426), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n464), .A2(new_n454), .A3(new_n457), .A4(new_n459), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT87), .B1(new_n465), .B2(new_n321), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n390), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n321), .B1(new_n460), .B2(new_n461), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT87), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n470), .A2(new_n442), .A3(new_n389), .A4(new_n462), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n388), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(G110), .B(G140), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n363), .A2(G227), .ZN(new_n474));
  XOR2_X1   g288(.A(new_n473), .B(new_n474), .Z(new_n475));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n228), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n230), .B1(new_n198), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n404), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n403), .B(new_n230), .C1(new_n231), .C2(new_n235), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n223), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT12), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(KEYINPUT12), .A3(new_n223), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n225), .A2(new_n205), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n487), .A2(new_n195), .A3(new_n420), .A4(new_n418), .ZN(new_n488));
  XOR2_X1   g302(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n489));
  NAND2_X1  g303(.A1(new_n479), .A2(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n399), .A2(new_n402), .A3(KEYINPUT10), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n236), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n488), .A2(new_n490), .A3(new_n221), .A4(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n476), .B1(new_n486), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n481), .A2(KEYINPUT12), .A3(new_n223), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT12), .B1(new_n481), .B2(new_n223), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n476), .B(new_n493), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n475), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n475), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT82), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n479), .A2(new_n489), .B1(new_n236), .B2(new_n491), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n221), .B1(new_n504), .B2(new_n488), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n493), .A2(KEYINPUT82), .A3(new_n500), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n499), .A2(G469), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G469), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(new_n321), .ZN(new_n511));
  AND4_X1   g325(.A1(new_n221), .A2(new_n488), .A3(new_n490), .A4(new_n492), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n475), .B1(new_n512), .B2(new_n505), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n500), .B(new_n493), .C1(new_n495), .C2(new_n496), .ZN(new_n514));
  AOI21_X1  g328(.A(G902), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n511), .B1(new_n515), .B2(new_n510), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n359), .A2(new_n344), .ZN(new_n518));
  INV_X1    g332(.A(G237), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n363), .A3(G214), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(new_n234), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n284), .A2(G143), .A3(G214), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n217), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(KEYINPUT90), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT90), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n525), .B(new_n217), .C1(new_n521), .C2(new_n522), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT17), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n284), .A2(G143), .A3(G214), .ZN(new_n528));
  AOI21_X1  g342(.A(G143), .B1(new_n284), .B2(G214), .ZN(new_n529));
  OAI21_X1  g343(.A(G131), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n525), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n523), .A2(KEYINPUT90), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n521), .A2(new_n217), .A3(new_n522), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n518), .A2(new_n527), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(G113), .B(G122), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(new_n392), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT18), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n521), .B(new_n522), .C1(new_n540), .C2(new_n217), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n539), .A2(new_n541), .B1(new_n523), .B2(KEYINPUT18), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n339), .A2(new_n340), .A3(G146), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT88), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT88), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n339), .A2(new_n340), .A3(new_n545), .A4(G146), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(new_n347), .A3(new_n546), .ZN(new_n547));
  OR2_X1    g361(.A1(new_n541), .A2(new_n539), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n542), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n536), .A2(new_n538), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n538), .B1(new_n536), .B2(new_n549), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n321), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G475), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT92), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n234), .A2(G128), .ZN(new_n555));
  OAI21_X1  g369(.A(G134), .B1(new_n555), .B2(KEYINPUT13), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n234), .A2(G128), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n228), .A2(G143), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n556), .A2(new_n559), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n261), .A2(G122), .A3(new_n262), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n252), .A2(G122), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n562), .A2(new_n395), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n395), .B1(new_n562), .B2(new_n563), .ZN(new_n565));
  OAI22_X1  g379(.A1(new_n560), .A2(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n562), .A2(new_n395), .A3(new_n563), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n557), .A2(new_n558), .A3(G134), .ZN(new_n568));
  AOI21_X1  g382(.A(G134), .B1(new_n557), .B2(new_n558), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT14), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n562), .A2(new_n571), .A3(new_n563), .ZN(new_n572));
  OAI21_X1  g386(.A(G107), .B1(new_n562), .B2(new_n571), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n567), .B(new_n570), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT9), .B(G234), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n575), .A2(new_n372), .A3(G953), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n566), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n566), .B2(new_n574), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n554), .B(new_n321), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G478), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT15), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n579), .B(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT20), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT19), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n346), .A2(KEYINPUT91), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT91), .ZN(new_n588));
  AOI22_X1  g402(.A1(new_n339), .A2(new_n340), .B1(new_n346), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n190), .B(new_n587), .C1(new_n589), .C2(new_n586), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n585), .A2(new_n345), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n549), .ZN(new_n592));
  INV_X1    g406(.A(new_n538), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n536), .A2(new_n538), .A3(new_n549), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(G475), .A2(G902), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n584), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n597), .ZN(new_n599));
  AOI211_X1 g413(.A(KEYINPUT20), .B(new_n599), .C1(new_n594), .C2(new_n595), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n553), .B(new_n583), .C1(new_n598), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n363), .A2(G952), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(G234), .B2(G237), .ZN(new_n603));
  AOI211_X1 g417(.A(new_n321), .B(new_n363), .C1(G234), .C2(G237), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT21), .B(G898), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G221), .B1(new_n575), .B2(G902), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n517), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n472), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n334), .A2(new_n386), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT93), .B(G101), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G3));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT94), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n467), .A2(new_n615), .A3(new_n471), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n387), .B1(new_n471), .B2(new_n615), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AND4_X1   g432(.A1(new_n389), .A2(new_n470), .A3(new_n442), .A4(new_n462), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n388), .B1(new_n619), .B2(KEYINPUT94), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n467), .A2(new_n615), .A3(new_n471), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT95), .ZN(new_n622));
  INV_X1    g436(.A(new_n606), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n580), .A2(new_n321), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  OR2_X1    g439(.A1(new_n577), .A2(new_n578), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n321), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n625), .B1(new_n627), .B2(G478), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n626), .B(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n628), .B1(new_n630), .B2(G478), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n553), .B1(new_n598), .B2(new_n600), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n618), .A2(new_n622), .A3(new_n623), .A4(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(G472), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n300), .B2(new_n321), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n302), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(KEYINPUT81), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n500), .B1(new_n641), .B2(new_n497), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n503), .A2(new_n506), .A3(new_n507), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n642), .A2(new_n643), .A3(new_n510), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n515), .A2(new_n510), .ZN(new_n645));
  INV_X1    g459(.A(new_n511), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n386), .B(new_n608), .C1(new_n644), .C2(new_n647), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n635), .A2(new_n639), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(KEYINPUT34), .B(G104), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G6));
  INV_X1    g465(.A(new_n583), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n652), .B(new_n553), .C1(new_n598), .C2(new_n600), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n618), .A2(new_n622), .A3(new_n623), .A4(new_n654), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n655), .A2(new_n639), .A3(new_n648), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT96), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT35), .B(G107), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  XOR2_X1   g473(.A(new_n361), .B(KEYINPUT97), .Z(new_n660));
  OR2_X1    g474(.A1(new_n367), .A2(KEYINPUT36), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n660), .B(new_n661), .Z(new_n662));
  INV_X1    g476(.A(new_n375), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n382), .A2(new_n385), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n472), .A2(new_n609), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n638), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT37), .B(G110), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G12));
  INV_X1    g484(.A(G900), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n604), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n603), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n653), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n334), .A2(new_n666), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n517), .A2(new_n608), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n618), .A2(new_n622), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n228), .ZN(G30));
  NAND2_X1  g496(.A1(new_n467), .A2(new_n471), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT38), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(new_n685));
  AOI22_X1  g499(.A1(new_n662), .A2(new_n663), .B1(new_n382), .B2(new_n385), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n632), .A2(new_n652), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n686), .A2(new_n387), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n300), .A2(KEYINPUT32), .A3(new_n301), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n323), .A2(new_n291), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n321), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n291), .B1(new_n277), .B2(new_n283), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n332), .A2(new_n696), .A3(new_n333), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n690), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT98), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n690), .A2(KEYINPUT98), .A3(new_n697), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n674), .B(KEYINPUT39), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n679), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n703), .B(KEYINPUT40), .Z(new_n704));
  NAND3_X1  g518(.A1(new_n700), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  NOR2_X1   g520(.A1(new_n633), .A2(new_n675), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n334), .A2(new_n666), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n680), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n188), .ZN(G48));
  OR2_X1    g524(.A1(new_n515), .A2(new_n510), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n645), .ZN(new_n712));
  INV_X1    g526(.A(new_n608), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n334), .A2(new_n386), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n635), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT41), .B(G113), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G15));
  NOR2_X1   g532(.A1(new_n715), .A2(new_n655), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n252), .ZN(G18));
  NAND3_X1  g534(.A1(new_n334), .A2(new_n607), .A3(new_n666), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n618), .A2(new_n622), .A3(new_n714), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n258), .ZN(G21));
  NAND3_X1  g538(.A1(new_n618), .A2(new_n622), .A3(new_n688), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT99), .B1(new_n306), .B2(new_n296), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT99), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n727), .B(new_n317), .C1(new_n323), .C2(new_n292), .ZN(new_n728));
  AND3_X1   g542(.A1(new_n726), .A2(new_n291), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n290), .A2(new_n299), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n301), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT100), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g547(.A(KEYINPUT100), .B(new_n301), .C1(new_n729), .C2(new_n730), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n637), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n712), .A2(new_n713), .A3(new_n606), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n386), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n725), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g552(.A(new_n738), .B(G122), .Z(G24));
  INV_X1    g553(.A(new_n637), .ZN(new_n740));
  INV_X1    g554(.A(new_n734), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n726), .A2(new_n728), .A3(new_n291), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n290), .A3(new_n299), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT100), .B1(new_n743), .B2(new_n301), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n740), .B(new_n666), .C1(new_n741), .C2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT101), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n733), .A2(new_n734), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n748), .A2(KEYINPUT101), .A3(new_n740), .A4(new_n666), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n618), .A2(new_n622), .A3(new_n707), .A4(new_n714), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  XNOR2_X1  g567(.A(new_n508), .B(KEYINPUT103), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(G469), .A3(new_n499), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n511), .B(KEYINPUT102), .Z(new_n756));
  AND2_X1   g570(.A1(new_n645), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n608), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n467), .A2(new_n387), .A3(new_n471), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n761), .A2(new_n707), .ZN(new_n762));
  INV_X1    g576(.A(new_n386), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n327), .B2(new_n330), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(KEYINPUT42), .A3(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n334), .A2(new_n386), .A3(new_n707), .A4(new_n761), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n766), .A2(KEYINPUT104), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT104), .B1(new_n766), .B2(new_n767), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n765), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G131), .ZN(G33));
  NAND4_X1  g585(.A1(new_n334), .A2(new_n386), .A3(new_n676), .A4(new_n761), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G134), .ZN(G36));
  NAND3_X1  g587(.A1(new_n754), .A2(KEYINPUT45), .A3(new_n499), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n774), .A2(KEYINPUT105), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(KEYINPUT105), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT45), .B1(new_n499), .B2(new_n508), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n510), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n775), .A2(new_n776), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT46), .B1(new_n779), .B2(new_n756), .ZN(new_n780));
  INV_X1    g594(.A(new_n645), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(KEYINPUT46), .A3(new_n756), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n713), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n631), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(new_n632), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n786), .B1(KEYINPUT106), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n789));
  OR3_X1    g603(.A1(new_n785), .A2(new_n632), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(KEYINPUT107), .A3(new_n790), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(new_n666), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n788), .A2(new_n790), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT107), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(new_n639), .A3(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT44), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n784), .A2(new_n798), .A3(new_n702), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n792), .A2(KEYINPUT44), .A3(new_n639), .A4(new_n795), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n760), .B(KEYINPUT108), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT109), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n800), .A2(KEYINPUT109), .A3(new_n801), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n799), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(new_n211), .ZN(G39));
  XNOR2_X1  g621(.A(new_n784), .B(KEYINPUT47), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT110), .ZN(new_n809));
  INV_X1    g623(.A(new_n760), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n763), .A3(new_n707), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n334), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n808), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n784), .A2(KEYINPUT47), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT47), .ZN(new_n815));
  AOI211_X1 g629(.A(new_n815), .B(new_n713), .C1(new_n782), .C2(new_n783), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n812), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT110), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G140), .ZN(G42));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n715), .B1(new_n635), .B2(new_n655), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n606), .B1(new_n633), .B2(new_n653), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n683), .A2(new_n387), .A3(new_n823), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n302), .A2(new_n637), .A3(new_n648), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n667), .A2(new_n638), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n826), .B(new_n611), .C1(new_n725), .C2(new_n737), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n822), .A2(new_n827), .A3(new_n723), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n750), .A2(new_n762), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n601), .A2(new_n675), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n760), .A2(new_n686), .A3(new_n678), .A4(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n334), .A2(new_n831), .A3(KEYINPUT113), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT113), .B1(new_n334), .B2(new_n831), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n772), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n828), .A2(new_n770), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n758), .A2(new_n686), .A3(new_n608), .A4(new_n674), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n697), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n838), .B1(new_n725), .B2(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n620), .A2(KEYINPUT95), .A3(new_n621), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT95), .B1(new_n620), .B2(new_n621), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT72), .B1(new_n328), .B2(new_n329), .ZN(new_n846));
  AOI211_X1 g660(.A(new_n331), .B(KEYINPUT32), .C1(new_n300), .C2(new_n301), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n839), .B1(new_n848), .B2(new_n696), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n845), .A2(new_n849), .A3(KEYINPUT114), .A4(new_n688), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n842), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n843), .A2(new_n844), .A3(new_n678), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n686), .B1(new_n848), .B2(new_n327), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n852), .B(new_n853), .C1(new_n676), .C2(new_n707), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n752), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n837), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n842), .A2(new_n850), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(KEYINPUT52), .A3(new_n752), .A4(new_n854), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n836), .A2(new_n859), .A3(KEYINPUT53), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT115), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n856), .A2(new_n862), .A3(new_n858), .ZN(new_n863));
  OAI211_X1 g677(.A(KEYINPUT115), .B(new_n837), .C1(new_n851), .C2(new_n855), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n863), .A2(new_n836), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n860), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n821), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n793), .A2(new_n603), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n810), .A2(new_n714), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n764), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT48), .Z(new_n873));
  XOR2_X1   g687(.A(new_n602), .B(KEYINPUT119), .Z(new_n874));
  NAND2_X1  g688(.A1(new_n735), .A2(new_n386), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n869), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OR4_X1    g691(.A1(new_n763), .A2(new_n697), .A3(new_n870), .A4(new_n673), .ZN(new_n878));
  OAI221_X1 g692(.A(new_n874), .B1(new_n877), .B2(new_n722), .C1(new_n878), .C2(new_n633), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n876), .A2(new_n388), .A3(new_n685), .A4(new_n714), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT50), .Z(new_n882));
  NAND2_X1  g696(.A1(new_n750), .A2(new_n871), .ZN(new_n883));
  OR3_X1    g697(.A1(new_n878), .A2(new_n632), .A3(new_n631), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n882), .A2(KEYINPUT51), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n876), .A2(new_n801), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n814), .A2(new_n816), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n711), .A2(new_n713), .A3(new_n645), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n880), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n808), .A2(KEYINPUT118), .ZN(new_n892));
  OR3_X1    g706(.A1(new_n814), .A2(new_n816), .A3(KEYINPUT118), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n892), .A2(new_n893), .A3(new_n888), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n891), .B1(new_n894), .B2(new_n886), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT51), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n836), .A2(new_n859), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n861), .ZN(new_n899));
  AND4_X1   g713(.A1(KEYINPUT53), .A2(new_n828), .A3(new_n770), .A4(new_n835), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n863), .A3(new_n901), .A4(new_n864), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n900), .A2(new_n863), .A3(new_n864), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT117), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n867), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n865), .A2(new_n861), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n836), .A2(new_n859), .A3(KEYINPUT53), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n909), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n868), .A2(new_n897), .A3(new_n906), .A4(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(G952), .B2(G953), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n786), .B1(KEYINPUT49), .B2(new_n712), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n913), .A2(new_n386), .A3(new_n387), .A4(new_n608), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT111), .Z(new_n915));
  NOR2_X1   g729(.A1(new_n712), .A2(KEYINPUT49), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n916), .B(KEYINPUT112), .Z(new_n917));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n685), .A3(new_n917), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n918), .A2(new_n697), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n912), .A2(new_n919), .ZN(G75));
  NOR2_X1   g734(.A1(new_n363), .A2(G952), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n921), .B(KEYINPUT120), .Z(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n905), .A2(new_n899), .A3(new_n902), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(G210), .A3(G902), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT56), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n433), .A2(new_n441), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(new_n440), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT55), .Z(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n925), .A2(new_n926), .A3(new_n930), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n923), .B1(new_n932), .B2(new_n933), .ZN(G51));
  XOR2_X1   g748(.A(new_n756), .B(KEYINPUT57), .Z(new_n935));
  AOI21_X1  g749(.A(new_n867), .B1(new_n903), .B2(new_n905), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n867), .A2(new_n905), .A3(new_n899), .A4(new_n902), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n513), .A2(new_n514), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n779), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n924), .A2(G902), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n921), .B1(new_n940), .B2(new_n942), .ZN(G54));
  NAND4_X1  g757(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n944));
  INV_X1    g758(.A(new_n596), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n944), .A2(KEYINPUT121), .A3(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n921), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n944), .B2(new_n945), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT121), .B1(new_n944), .B2(new_n945), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(G60));
  INV_X1    g764(.A(new_n630), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n868), .A2(new_n906), .A3(new_n910), .ZN(new_n952));
  XNOR2_X1  g766(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n625), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n951), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n951), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n936), .B2(new_n937), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n922), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n955), .A2(new_n958), .ZN(G63));
  XNOR2_X1  g773(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n372), .A2(new_n321), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n924), .A2(new_n662), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n962), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n964), .B1(new_n903), .B2(new_n905), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n369), .A2(new_n371), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n963), .B(new_n922), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n924), .A2(new_n962), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n369), .B2(new_n371), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n971), .A2(KEYINPUT61), .A3(new_n922), .A4(new_n963), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n969), .A2(new_n972), .ZN(G66));
  INV_X1    g787(.A(new_n605), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n363), .B1(new_n974), .B2(G224), .ZN(new_n975));
  INV_X1    g789(.A(new_n828), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n976), .B2(new_n363), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n928), .B1(G898), .B2(new_n363), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n977), .B(new_n978), .Z(G69));
  AOI21_X1  g793(.A(new_n363), .B1(G227), .B2(G900), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n806), .B1(new_n813), .B2(new_n818), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n770), .A2(new_n772), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT125), .ZN(new_n983));
  INV_X1    g797(.A(new_n725), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n784), .A2(new_n702), .A3(new_n984), .A4(new_n764), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n618), .A2(new_n622), .A3(new_n707), .A4(new_n714), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n747), .B2(new_n749), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n680), .B1(new_n677), .B2(new_n708), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n981), .A2(new_n983), .A3(new_n363), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n244), .A2(new_n276), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n587), .B1(new_n589), .B2(new_n586), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n993), .B(new_n994), .Z(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(G900), .B2(G953), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n980), .B1(new_n997), .B2(KEYINPUT124), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n705), .A2(new_n989), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT62), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  AOI211_X1 g815(.A(new_n703), .B(new_n760), .C1(new_n633), .C2(new_n653), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1002), .A2(new_n334), .A3(new_n386), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n981), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n363), .ZN(new_n1005));
  AOI22_X1  g819(.A1(new_n1005), .A2(new_n995), .B1(new_n992), .B2(new_n996), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n998), .B(new_n1006), .ZN(G72));
  NAND2_X1  g821(.A1(new_n311), .A2(new_n289), .ZN(new_n1008));
  XNOR2_X1  g822(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n636), .A2(new_n321), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n947), .B1(new_n866), .B2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n981), .A2(new_n983), .A3(new_n828), .A4(new_n991), .ZN(new_n1014));
  AOI211_X1 g828(.A(new_n288), .B(new_n310), .C1(new_n1014), .C2(new_n1011), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n981), .A2(new_n1001), .A3(new_n828), .A4(new_n1003), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(KEYINPUT127), .A3(new_n1011), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n1017), .A2(new_n694), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1016), .A2(new_n1011), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT127), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI211_X1 g835(.A(new_n1013), .B(new_n1015), .C1(new_n1018), .C2(new_n1021), .ZN(G57));
endmodule


