

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X2 U548 ( .A(n520), .B(KEYINPUT65), .ZN(n666) );
  INV_X1 U549 ( .A(KEYINPUT28), .ZN(n682) );
  NAND2_X1 U550 ( .A1(n767), .A2(n510), .ZN(n802) );
  AND2_X1 U551 ( .A1(n766), .A2(n765), .ZN(n510) );
  NOR2_X1 U552 ( .A1(n801), .A2(n800), .ZN(n511) );
  NOR2_X1 U553 ( .A1(n749), .A2(n748), .ZN(n512) );
  NOR2_X1 U554 ( .A1(n723), .A2(n722), .ZN(n513) );
  INV_X1 U555 ( .A(n726), .ZN(n690) );
  NAND2_X1 U556 ( .A1(n709), .A2(G8), .ZN(n710) );
  XNOR2_X1 U557 ( .A(n710), .B(KEYINPUT96), .ZN(n712) );
  NOR2_X1 U558 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U559 ( .A(KEYINPUT99), .B(KEYINPUT32), .ZN(n740) );
  NAND2_X1 U560 ( .A1(n676), .A2(n769), .ZN(n726) );
  INV_X1 U561 ( .A(n811), .ZN(n801) );
  AND2_X1 U562 ( .A1(n521), .A2(G2104), .ZN(n878) );
  NOR2_X1 U563 ( .A1(G2104), .A2(n521), .ZN(n881) );
  NOR2_X1 U564 ( .A1(G651), .A2(n623), .ZN(n631) );
  INV_X1 U565 ( .A(KEYINPUT85), .ZN(n669) );
  AND2_X1 U566 ( .A1(n519), .A2(n518), .ZN(n675) );
  INV_X1 U567 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U568 ( .A1(G101), .A2(n878), .ZN(n514) );
  XNOR2_X1 U569 ( .A(KEYINPUT64), .B(n514), .ZN(n516) );
  INV_X1 U570 ( .A(KEYINPUT23), .ZN(n515) );
  XNOR2_X1 U571 ( .A(n516), .B(n515), .ZN(n519) );
  NOR2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  XOR2_X2 U573 ( .A(KEYINPUT17), .B(n517), .Z(n877) );
  NAND2_X1 U574 ( .A1(G137), .A2(n877), .ZN(n518) );
  NAND2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  NAND2_X1 U576 ( .A1(G113), .A2(n666), .ZN(n523) );
  NAND2_X1 U577 ( .A1(G125), .A2(n881), .ZN(n522) );
  AND2_X1 U578 ( .A1(n523), .A2(n522), .ZN(n673) );
  AND2_X1 U579 ( .A1(n675), .A2(n673), .ZN(G160) );
  INV_X1 U580 ( .A(G651), .ZN(n527) );
  NOR2_X1 U581 ( .A1(G543), .A2(n527), .ZN(n524) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n524), .Z(n630) );
  NAND2_X1 U583 ( .A1(G64), .A2(n630), .ZN(n526) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n623) );
  NAND2_X1 U585 ( .A1(G52), .A2(n631), .ZN(n525) );
  NAND2_X1 U586 ( .A1(n526), .A2(n525), .ZN(n532) );
  NOR2_X1 U587 ( .A1(G651), .A2(G543), .ZN(n626) );
  NAND2_X1 U588 ( .A1(G90), .A2(n626), .ZN(n529) );
  NOR2_X1 U589 ( .A1(n623), .A2(n527), .ZN(n627) );
  NAND2_X1 U590 ( .A1(G77), .A2(n627), .ZN(n528) );
  NAND2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U592 ( .A(KEYINPUT9), .B(n530), .Z(n531) );
  NOR2_X1 U593 ( .A1(n532), .A2(n531), .ZN(G171) );
  NAND2_X1 U594 ( .A1(G99), .A2(n878), .ZN(n539) );
  NAND2_X1 U595 ( .A1(G111), .A2(n666), .ZN(n534) );
  NAND2_X1 U596 ( .A1(G135), .A2(n877), .ZN(n533) );
  NAND2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n537) );
  NAND2_X1 U598 ( .A1(n881), .A2(G123), .ZN(n535) );
  XOR2_X1 U599 ( .A(KEYINPUT18), .B(n535), .Z(n536) );
  NOR2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U602 ( .A(n540), .B(KEYINPUT76), .ZN(n924) );
  XNOR2_X1 U603 ( .A(n924), .B(G2096), .ZN(n541) );
  OR2_X1 U604 ( .A1(G2100), .A2(n541), .ZN(G156) );
  INV_X1 U605 ( .A(G120), .ZN(G236) );
  INV_X1 U606 ( .A(G69), .ZN(G235) );
  INV_X1 U607 ( .A(G108), .ZN(G238) );
  INV_X1 U608 ( .A(G82), .ZN(G220) );
  NAND2_X1 U609 ( .A1(G65), .A2(n630), .ZN(n543) );
  NAND2_X1 U610 ( .A1(G53), .A2(n631), .ZN(n542) );
  NAND2_X1 U611 ( .A1(n543), .A2(n542), .ZN(n547) );
  NAND2_X1 U612 ( .A1(G91), .A2(n626), .ZN(n545) );
  NAND2_X1 U613 ( .A1(G78), .A2(n627), .ZN(n544) );
  NAND2_X1 U614 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n685) );
  INV_X1 U616 ( .A(n685), .ZN(G299) );
  NAND2_X1 U617 ( .A1(G88), .A2(n626), .ZN(n549) );
  NAND2_X1 U618 ( .A1(G75), .A2(n627), .ZN(n548) );
  NAND2_X1 U619 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U620 ( .A1(G62), .A2(n630), .ZN(n551) );
  NAND2_X1 U621 ( .A1(G50), .A2(n631), .ZN(n550) );
  NAND2_X1 U622 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U623 ( .A1(n553), .A2(n552), .ZN(G166) );
  NAND2_X1 U624 ( .A1(G63), .A2(n630), .ZN(n555) );
  NAND2_X1 U625 ( .A1(G51), .A2(n631), .ZN(n554) );
  NAND2_X1 U626 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U627 ( .A(KEYINPUT6), .B(n556), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n627), .A2(G76), .ZN(n557) );
  XNOR2_X1 U629 ( .A(KEYINPUT74), .B(n557), .ZN(n561) );
  XOR2_X1 U630 ( .A(KEYINPUT4), .B(KEYINPUT73), .Z(n559) );
  NAND2_X1 U631 ( .A1(G89), .A2(n626), .ZN(n558) );
  XNOR2_X1 U632 ( .A(n559), .B(n558), .ZN(n560) );
  NAND2_X1 U633 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U634 ( .A(n562), .B(KEYINPUT5), .Z(n563) );
  NOR2_X1 U635 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U636 ( .A(KEYINPUT7), .B(n565), .Z(n566) );
  XOR2_X1 U637 ( .A(KEYINPUT75), .B(n566), .Z(G168) );
  XOR2_X1 U638 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U639 ( .A1(G94), .A2(G452), .ZN(n567) );
  XOR2_X1 U640 ( .A(KEYINPUT68), .B(n567), .Z(G173) );
  NAND2_X1 U641 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U642 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U643 ( .A(G223), .ZN(n833) );
  NAND2_X1 U644 ( .A1(n833), .A2(G567), .ZN(n569) );
  XOR2_X1 U645 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U646 ( .A1(G56), .A2(n630), .ZN(n570) );
  XOR2_X1 U647 ( .A(KEYINPUT14), .B(n570), .Z(n576) );
  NAND2_X1 U648 ( .A1(n626), .A2(G81), .ZN(n571) );
  XNOR2_X1 U649 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U650 ( .A1(G68), .A2(n627), .ZN(n572) );
  NAND2_X1 U651 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U652 ( .A(KEYINPUT13), .B(n574), .Z(n575) );
  NOR2_X1 U653 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U654 ( .A1(n631), .A2(G43), .ZN(n577) );
  NAND2_X1 U655 ( .A1(n578), .A2(n577), .ZN(n993) );
  INV_X1 U656 ( .A(G860), .ZN(n600) );
  OR2_X1 U657 ( .A1(n993), .A2(n600), .ZN(G153) );
  XOR2_X1 U658 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  INV_X1 U659 ( .A(G868), .ZN(n590) );
  NOR2_X1 U660 ( .A1(G301), .A2(n590), .ZN(n588) );
  NAND2_X1 U661 ( .A1(n631), .A2(G54), .ZN(n585) );
  NAND2_X1 U662 ( .A1(G66), .A2(n630), .ZN(n580) );
  NAND2_X1 U663 ( .A1(G79), .A2(n627), .ZN(n579) );
  NAND2_X1 U664 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U665 ( .A1(G92), .A2(n626), .ZN(n581) );
  XNOR2_X1 U666 ( .A(KEYINPUT71), .B(n581), .ZN(n582) );
  NOR2_X1 U667 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U668 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U669 ( .A(KEYINPUT15), .B(n586), .Z(n994) );
  NOR2_X1 U670 ( .A1(G868), .A2(n994), .ZN(n587) );
  NOR2_X1 U671 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U672 ( .A(KEYINPUT72), .B(n589), .ZN(G284) );
  NOR2_X1 U673 ( .A1(G286), .A2(n590), .ZN(n592) );
  NOR2_X1 U674 ( .A1(G868), .A2(G299), .ZN(n591) );
  NOR2_X1 U675 ( .A1(n592), .A2(n591), .ZN(G297) );
  NAND2_X1 U676 ( .A1(n600), .A2(G559), .ZN(n593) );
  INV_X1 U677 ( .A(n994), .ZN(n598) );
  NAND2_X1 U678 ( .A1(n593), .A2(n598), .ZN(n594) );
  XNOR2_X1 U679 ( .A(n594), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n993), .ZN(n597) );
  NAND2_X1 U681 ( .A1(G868), .A2(n598), .ZN(n595) );
  NOR2_X1 U682 ( .A1(G559), .A2(n595), .ZN(n596) );
  NOR2_X1 U683 ( .A1(n597), .A2(n596), .ZN(G282) );
  XOR2_X1 U684 ( .A(KEYINPUT77), .B(KEYINPUT80), .Z(n602) );
  NAND2_X1 U685 ( .A1(G559), .A2(n598), .ZN(n599) );
  XOR2_X1 U686 ( .A(n993), .B(n599), .Z(n643) );
  NAND2_X1 U687 ( .A1(n643), .A2(n600), .ZN(n601) );
  XNOR2_X1 U688 ( .A(n602), .B(n601), .ZN(n611) );
  NAND2_X1 U689 ( .A1(G67), .A2(n630), .ZN(n604) );
  NAND2_X1 U690 ( .A1(G55), .A2(n631), .ZN(n603) );
  NAND2_X1 U691 ( .A1(n604), .A2(n603), .ZN(n610) );
  NAND2_X1 U692 ( .A1(n627), .A2(G80), .ZN(n605) );
  XNOR2_X1 U693 ( .A(n605), .B(KEYINPUT78), .ZN(n607) );
  NAND2_X1 U694 ( .A1(G93), .A2(n626), .ZN(n606) );
  NAND2_X1 U695 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U696 ( .A(KEYINPUT79), .B(n608), .Z(n609) );
  NOR2_X1 U697 ( .A1(n610), .A2(n609), .ZN(n645) );
  XOR2_X1 U698 ( .A(n611), .B(n645), .Z(G145) );
  NAND2_X1 U699 ( .A1(G61), .A2(n630), .ZN(n613) );
  NAND2_X1 U700 ( .A1(G86), .A2(n626), .ZN(n612) );
  NAND2_X1 U701 ( .A1(n613), .A2(n612), .ZN(n616) );
  NAND2_X1 U702 ( .A1(n627), .A2(G73), .ZN(n614) );
  XOR2_X1 U703 ( .A(KEYINPUT2), .B(n614), .Z(n615) );
  NOR2_X1 U704 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U705 ( .A(KEYINPUT81), .B(n617), .Z(n619) );
  NAND2_X1 U706 ( .A1(n631), .A2(G48), .ZN(n618) );
  NAND2_X1 U707 ( .A1(n619), .A2(n618), .ZN(G305) );
  NAND2_X1 U708 ( .A1(G49), .A2(n631), .ZN(n621) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n620) );
  NAND2_X1 U710 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U711 ( .A1(n630), .A2(n622), .ZN(n625) );
  NAND2_X1 U712 ( .A1(n623), .A2(G87), .ZN(n624) );
  NAND2_X1 U713 ( .A1(n625), .A2(n624), .ZN(G288) );
  NAND2_X1 U714 ( .A1(G85), .A2(n626), .ZN(n629) );
  NAND2_X1 U715 ( .A1(G72), .A2(n627), .ZN(n628) );
  NAND2_X1 U716 ( .A1(n629), .A2(n628), .ZN(n636) );
  NAND2_X1 U717 ( .A1(G60), .A2(n630), .ZN(n633) );
  NAND2_X1 U718 ( .A1(G47), .A2(n631), .ZN(n632) );
  NAND2_X1 U719 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U720 ( .A(KEYINPUT66), .B(n634), .ZN(n635) );
  NOR2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U722 ( .A(n637), .B(KEYINPUT67), .ZN(G290) );
  XNOR2_X1 U723 ( .A(G288), .B(KEYINPUT19), .ZN(n639) );
  XNOR2_X1 U724 ( .A(n685), .B(G166), .ZN(n638) );
  XNOR2_X1 U725 ( .A(n639), .B(n638), .ZN(n640) );
  XOR2_X1 U726 ( .A(n645), .B(n640), .Z(n641) );
  XNOR2_X1 U727 ( .A(G305), .B(n641), .ZN(n642) );
  XNOR2_X1 U728 ( .A(n642), .B(G290), .ZN(n904) );
  XNOR2_X1 U729 ( .A(n643), .B(n904), .ZN(n644) );
  NAND2_X1 U730 ( .A1(n644), .A2(G868), .ZN(n647) );
  OR2_X1 U731 ( .A1(G868), .A2(n645), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n647), .A2(n646), .ZN(G295) );
  NAND2_X1 U733 ( .A1(G2084), .A2(G2078), .ZN(n648) );
  XOR2_X1 U734 ( .A(KEYINPUT20), .B(n648), .Z(n649) );
  NAND2_X1 U735 ( .A1(G2090), .A2(n649), .ZN(n650) );
  XNOR2_X1 U736 ( .A(KEYINPUT21), .B(n650), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n651), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U738 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U739 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U740 ( .A1(G220), .A2(G219), .ZN(n652) );
  XOR2_X1 U741 ( .A(KEYINPUT22), .B(n652), .Z(n653) );
  NOR2_X1 U742 ( .A1(G218), .A2(n653), .ZN(n654) );
  NAND2_X1 U743 ( .A1(G96), .A2(n654), .ZN(n838) );
  NAND2_X1 U744 ( .A1(G2106), .A2(n838), .ZN(n660) );
  NOR2_X1 U745 ( .A1(G235), .A2(G236), .ZN(n655) );
  XOR2_X1 U746 ( .A(KEYINPUT82), .B(n655), .Z(n656) );
  NOR2_X1 U747 ( .A1(G238), .A2(n656), .ZN(n657) );
  NAND2_X1 U748 ( .A1(G57), .A2(n657), .ZN(n837) );
  NAND2_X1 U749 ( .A1(G567), .A2(n837), .ZN(n658) );
  XOR2_X1 U750 ( .A(KEYINPUT83), .B(n658), .Z(n659) );
  NAND2_X1 U751 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U752 ( .A(KEYINPUT84), .B(n661), .Z(G319) );
  INV_X1 U753 ( .A(G319), .ZN(n663) );
  NAND2_X1 U754 ( .A1(G661), .A2(G483), .ZN(n662) );
  NOR2_X1 U755 ( .A1(n663), .A2(n662), .ZN(n836) );
  NAND2_X1 U756 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U757 ( .A1(G138), .A2(n877), .ZN(n665) );
  NAND2_X1 U758 ( .A1(G102), .A2(n878), .ZN(n664) );
  NAND2_X1 U759 ( .A1(n665), .A2(n664), .ZN(n672) );
  NAND2_X1 U760 ( .A1(G126), .A2(n881), .ZN(n668) );
  NAND2_X1 U761 ( .A1(G114), .A2(n666), .ZN(n667) );
  NAND2_X1 U762 ( .A1(n668), .A2(n667), .ZN(n670) );
  XNOR2_X1 U763 ( .A(n670), .B(n669), .ZN(n671) );
  NOR2_X1 U764 ( .A1(n672), .A2(n671), .ZN(G164) );
  INV_X1 U765 ( .A(G166), .ZN(G303) );
  AND2_X1 U766 ( .A1(G40), .A2(n673), .ZN(n674) );
  NAND2_X1 U767 ( .A1(n675), .A2(n674), .ZN(n768) );
  XNOR2_X1 U768 ( .A(KEYINPUT91), .B(n768), .ZN(n676) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n769) );
  NAND2_X1 U770 ( .A1(n690), .A2(G2072), .ZN(n677) );
  XNOR2_X1 U771 ( .A(KEYINPUT27), .B(n677), .ZN(n680) );
  NAND2_X1 U772 ( .A1(G1956), .A2(n726), .ZN(n678) );
  XNOR2_X1 U773 ( .A(KEYINPUT93), .B(n678), .ZN(n679) );
  NOR2_X1 U774 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U775 ( .A(n681), .B(KEYINPUT94), .ZN(n684) );
  NOR2_X1 U776 ( .A1(n684), .A2(n685), .ZN(n683) );
  XNOR2_X1 U777 ( .A(n683), .B(n682), .ZN(n701) );
  NAND2_X1 U778 ( .A1(n685), .A2(n684), .ZN(n699) );
  INV_X1 U779 ( .A(G1996), .ZN(n943) );
  NOR2_X1 U780 ( .A1(n726), .A2(n943), .ZN(n686) );
  XOR2_X1 U781 ( .A(n686), .B(KEYINPUT26), .Z(n688) );
  NAND2_X1 U782 ( .A1(n726), .A2(G1341), .ZN(n687) );
  NAND2_X1 U783 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U784 ( .A1(n993), .A2(n689), .ZN(n694) );
  NAND2_X1 U785 ( .A1(G1348), .A2(n726), .ZN(n692) );
  NAND2_X1 U786 ( .A1(G2067), .A2(n690), .ZN(n691) );
  NAND2_X1 U787 ( .A1(n692), .A2(n691), .ZN(n695) );
  NOR2_X1 U788 ( .A1(n994), .A2(n695), .ZN(n693) );
  OR2_X1 U789 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n994), .A2(n695), .ZN(n696) );
  NAND2_X1 U791 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U794 ( .A(KEYINPUT29), .B(n702), .ZN(n703) );
  INV_X1 U795 ( .A(n703), .ZN(n708) );
  OR2_X1 U796 ( .A1(n690), .A2(G1961), .ZN(n705) );
  XNOR2_X1 U797 ( .A(G2078), .B(KEYINPUT25), .ZN(n942) );
  NAND2_X1 U798 ( .A1(n690), .A2(n942), .ZN(n704) );
  NAND2_X1 U799 ( .A1(n705), .A2(n704), .ZN(n714) );
  NAND2_X1 U800 ( .A1(G171), .A2(n714), .ZN(n706) );
  XNOR2_X1 U801 ( .A(n706), .B(KEYINPUT92), .ZN(n707) );
  NAND2_X1 U802 ( .A1(n708), .A2(n707), .ZN(n734) );
  INV_X1 U803 ( .A(KEYINPUT31), .ZN(n718) );
  NAND2_X1 U804 ( .A1(G8), .A2(n726), .ZN(n749) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n749), .ZN(n722) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n726), .ZN(n721) );
  NOR2_X1 U807 ( .A1(n722), .A2(n721), .ZN(n709) );
  XOR2_X1 U808 ( .A(KEYINPUT30), .B(KEYINPUT95), .Z(n711) );
  XNOR2_X1 U809 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U810 ( .A1(G168), .A2(n713), .ZN(n716) );
  NOR2_X1 U811 ( .A1(G171), .A2(n714), .ZN(n715) );
  XNOR2_X1 U812 ( .A(n718), .B(n717), .ZN(n732) );
  NAND2_X1 U813 ( .A1(n734), .A2(n732), .ZN(n720) );
  INV_X1 U814 ( .A(KEYINPUT97), .ZN(n719) );
  XNOR2_X1 U815 ( .A(n720), .B(n719), .ZN(n724) );
  AND2_X1 U816 ( .A1(G8), .A2(n721), .ZN(n723) );
  AND2_X1 U817 ( .A1(n724), .A2(n513), .ZN(n743) );
  INV_X1 U818 ( .A(G8), .ZN(n731) );
  BUF_X1 U819 ( .A(n749), .Z(n764) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n764), .ZN(n725) );
  XNOR2_X1 U821 ( .A(n725), .B(KEYINPUT98), .ZN(n728) );
  NOR2_X1 U822 ( .A1(n726), .A2(G2090), .ZN(n727) );
  NOR2_X1 U823 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U824 ( .A1(n729), .A2(G303), .ZN(n730) );
  OR2_X1 U825 ( .A1(n731), .A2(n730), .ZN(n735) );
  AND2_X1 U826 ( .A1(n732), .A2(n735), .ZN(n733) );
  NAND2_X1 U827 ( .A1(n734), .A2(n733), .ZN(n739) );
  INV_X1 U828 ( .A(n735), .ZN(n737) );
  AND2_X1 U829 ( .A1(G286), .A2(G8), .ZN(n736) );
  OR2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n741) );
  XNOR2_X1 U832 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n757) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n997) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U836 ( .A1(n997), .A2(n744), .ZN(n745) );
  XOR2_X1 U837 ( .A(KEYINPUT100), .B(n745), .Z(n746) );
  NOR2_X1 U838 ( .A1(n757), .A2(n746), .ZN(n747) );
  XNOR2_X1 U839 ( .A(n747), .B(KEYINPUT101), .ZN(n750) );
  NAND2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n998) );
  INV_X1 U841 ( .A(n998), .ZN(n748) );
  AND2_X1 U842 ( .A1(n750), .A2(n512), .ZN(n751) );
  NOR2_X1 U843 ( .A1(n751), .A2(KEYINPUT33), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n997), .A2(KEYINPUT33), .ZN(n752) );
  OR2_X1 U845 ( .A1(n752), .A2(n764), .ZN(n753) );
  XOR2_X1 U846 ( .A(G1981), .B(G305), .Z(n986) );
  NAND2_X1 U847 ( .A1(n753), .A2(n986), .ZN(n754) );
  NOR2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n756) );
  INV_X1 U849 ( .A(n756), .ZN(n767) );
  INV_X1 U850 ( .A(n757), .ZN(n760) );
  NOR2_X1 U851 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U852 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U853 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U854 ( .A1(n761), .A2(n764), .ZN(n766) );
  NOR2_X1 U855 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XOR2_X1 U856 ( .A(n762), .B(KEYINPUT24), .Z(n763) );
  OR2_X1 U857 ( .A1(n764), .A2(n763), .ZN(n765) );
  NOR2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n817) );
  XNOR2_X1 U859 ( .A(G2067), .B(KEYINPUT37), .ZN(n770) );
  XOR2_X1 U860 ( .A(n770), .B(KEYINPUT86), .Z(n813) );
  NAND2_X1 U861 ( .A1(G140), .A2(n877), .ZN(n772) );
  NAND2_X1 U862 ( .A1(G104), .A2(n878), .ZN(n771) );
  NAND2_X1 U863 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U864 ( .A(KEYINPUT34), .B(n773), .ZN(n779) );
  NAND2_X1 U865 ( .A1(n666), .A2(G116), .ZN(n774) );
  XOR2_X1 U866 ( .A(KEYINPUT87), .B(n774), .Z(n776) );
  NAND2_X1 U867 ( .A1(n881), .A2(G128), .ZN(n775) );
  NAND2_X1 U868 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U869 ( .A(KEYINPUT35), .B(n777), .Z(n778) );
  NOR2_X1 U870 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U871 ( .A(KEYINPUT36), .B(n780), .Z(n895) );
  AND2_X1 U872 ( .A1(n813), .A2(n895), .ZN(n934) );
  NAND2_X1 U873 ( .A1(n817), .A2(n934), .ZN(n811) );
  NAND2_X1 U874 ( .A1(n878), .A2(G105), .ZN(n782) );
  XNOR2_X1 U875 ( .A(KEYINPUT90), .B(KEYINPUT38), .ZN(n781) );
  XNOR2_X1 U876 ( .A(n782), .B(n781), .ZN(n789) );
  NAND2_X1 U877 ( .A1(G117), .A2(n666), .ZN(n784) );
  NAND2_X1 U878 ( .A1(G141), .A2(n877), .ZN(n783) );
  NAND2_X1 U879 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G129), .A2(n881), .ZN(n785) );
  XNOR2_X1 U881 ( .A(KEYINPUT89), .B(n785), .ZN(n786) );
  NOR2_X1 U882 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U883 ( .A1(n789), .A2(n788), .ZN(n899) );
  NAND2_X1 U884 ( .A1(G1996), .A2(n899), .ZN(n798) );
  NAND2_X1 U885 ( .A1(G119), .A2(n881), .ZN(n791) );
  NAND2_X1 U886 ( .A1(G95), .A2(n878), .ZN(n790) );
  NAND2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n877), .A2(G131), .ZN(n792) );
  XOR2_X1 U889 ( .A(KEYINPUT88), .B(n792), .Z(n793) );
  NOR2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n796) );
  NAND2_X1 U891 ( .A1(n666), .A2(G107), .ZN(n795) );
  NAND2_X1 U892 ( .A1(n796), .A2(n795), .ZN(n888) );
  NAND2_X1 U893 ( .A1(G1991), .A2(n888), .ZN(n797) );
  NAND2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n922) );
  NAND2_X1 U895 ( .A1(n817), .A2(n922), .ZN(n804) );
  XNOR2_X1 U896 ( .A(G1986), .B(G290), .ZN(n990) );
  NAND2_X1 U897 ( .A1(n817), .A2(n990), .ZN(n799) );
  NAND2_X1 U898 ( .A1(n804), .A2(n799), .ZN(n800) );
  NAND2_X1 U899 ( .A1(n802), .A2(n511), .ZN(n803) );
  XNOR2_X1 U900 ( .A(n803), .B(KEYINPUT102), .ZN(n819) );
  NOR2_X1 U901 ( .A1(G1996), .A2(n899), .ZN(n915) );
  INV_X1 U902 ( .A(n804), .ZN(n807) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n805) );
  NOR2_X1 U904 ( .A1(G1991), .A2(n888), .ZN(n918) );
  NOR2_X1 U905 ( .A1(n805), .A2(n918), .ZN(n806) );
  NOR2_X1 U906 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U907 ( .A(KEYINPUT103), .B(n808), .Z(n809) );
  NOR2_X1 U908 ( .A1(n915), .A2(n809), .ZN(n810) );
  XNOR2_X1 U909 ( .A(KEYINPUT39), .B(n810), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n812), .A2(n811), .ZN(n815) );
  NOR2_X1 U911 ( .A1(n895), .A2(n813), .ZN(n814) );
  XOR2_X1 U912 ( .A(KEYINPUT104), .B(n814), .Z(n932) );
  NAND2_X1 U913 ( .A1(n815), .A2(n932), .ZN(n816) );
  NAND2_X1 U914 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n822) );
  XOR2_X1 U916 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n820) );
  XNOR2_X1 U917 ( .A(KEYINPUT40), .B(n820), .ZN(n821) );
  XNOR2_X1 U918 ( .A(n822), .B(n821), .ZN(G329) );
  XOR2_X1 U919 ( .A(G2454), .B(G2435), .Z(n824) );
  XNOR2_X1 U920 ( .A(G2438), .B(G2427), .ZN(n823) );
  XNOR2_X1 U921 ( .A(n824), .B(n823), .ZN(n831) );
  XOR2_X1 U922 ( .A(KEYINPUT107), .B(G2446), .Z(n826) );
  XNOR2_X1 U923 ( .A(G2443), .B(G2430), .ZN(n825) );
  XNOR2_X1 U924 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U925 ( .A(n827), .B(G2451), .Z(n829) );
  XNOR2_X1 U926 ( .A(G1341), .B(G1348), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n830) );
  XNOR2_X1 U928 ( .A(n831), .B(n830), .ZN(n832) );
  NAND2_X1 U929 ( .A1(n832), .A2(G14), .ZN(n908) );
  XOR2_X1 U930 ( .A(KEYINPUT108), .B(n908), .Z(G401) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n833), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U933 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U935 ( .A1(n836), .A2(n835), .ZN(G188) );
  NOR2_X1 U936 ( .A1(n838), .A2(n837), .ZN(G325) );
  XNOR2_X1 U937 ( .A(KEYINPUT109), .B(G325), .ZN(G261) );
  XOR2_X1 U938 ( .A(G1976), .B(G1971), .Z(n840) );
  XNOR2_X1 U939 ( .A(G1986), .B(G1961), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(n850) );
  XOR2_X1 U941 ( .A(KEYINPUT111), .B(KEYINPUT113), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1996), .B(KEYINPUT41), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U944 ( .A(G1981), .B(G1956), .Z(n844) );
  XNOR2_X1 U945 ( .A(G1991), .B(G1966), .ZN(n843) );
  XNOR2_X1 U946 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U947 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U948 ( .A(KEYINPUT112), .B(G2474), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U950 ( .A(n850), .B(n849), .Z(G229) );
  XOR2_X1 U951 ( .A(G2096), .B(KEYINPUT43), .Z(n852) );
  XNOR2_X1 U952 ( .A(G2090), .B(KEYINPUT110), .ZN(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U954 ( .A(n853), .B(G2678), .Z(n855) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2072), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U957 ( .A(KEYINPUT42), .B(G2100), .Z(n857) );
  XNOR2_X1 U958 ( .A(G2084), .B(G2078), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(G227) );
  NAND2_X1 U961 ( .A1(G124), .A2(n881), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n860), .B(KEYINPUT114), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n861), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U964 ( .A1(G112), .A2(n666), .ZN(n862) );
  NAND2_X1 U965 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G136), .A2(n877), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G100), .A2(n878), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U969 ( .A1(n867), .A2(n866), .ZN(G162) );
  NAND2_X1 U970 ( .A1(n878), .A2(G106), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n868), .B(KEYINPUT116), .ZN(n870) );
  NAND2_X1 U972 ( .A1(G142), .A2(n877), .ZN(n869) );
  NAND2_X1 U973 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n871), .B(KEYINPUT45), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G118), .A2(n666), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G130), .A2(n881), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n874), .B(KEYINPUT115), .ZN(n875) );
  NOR2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n890) );
  NAND2_X1 U980 ( .A1(G139), .A2(n877), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G103), .A2(n878), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U983 ( .A1(G115), .A2(n666), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G127), .A2(n881), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U986 ( .A(KEYINPUT47), .B(n884), .ZN(n885) );
  XNOR2_X1 U987 ( .A(KEYINPUT117), .B(n885), .ZN(n886) );
  NOR2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n925) );
  XOR2_X1 U989 ( .A(n888), .B(n925), .Z(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n894) );
  XOR2_X1 U991 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n892) );
  XNOR2_X1 U992 ( .A(n924), .B(KEYINPUT118), .ZN(n891) );
  XNOR2_X1 U993 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U994 ( .A(n894), .B(n893), .Z(n897) );
  XNOR2_X1 U995 ( .A(G160), .B(n895), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n901) );
  XOR2_X1 U997 ( .A(G164), .B(G162), .Z(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U1001 ( .A(G171), .B(G286), .Z(n903) );
  XNOR2_X1 U1002 ( .A(n994), .B(n903), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n993), .B(n904), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n907), .ZN(G397) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n908), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(G229), .A2(G227), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(G225) );
  XNOR2_X1 U1012 ( .A(KEYINPUT119), .B(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G96), .ZN(G221) );
  INV_X1 U1015 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1016 ( .A(G2090), .B(G162), .Z(n914) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1018 ( .A(KEYINPUT51), .B(n916), .Z(n920) );
  XOR2_X1 U1019 ( .A(G160), .B(G2084), .Z(n917) );
  NOR2_X1 U1020 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n930) );
  XOR2_X1 U1024 ( .A(G2072), .B(n925), .Z(n927) );
  XOR2_X1 U1025 ( .A(G164), .B(G2078), .Z(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1027 ( .A(KEYINPUT50), .B(n928), .Z(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1031 ( .A(KEYINPUT52), .B(n935), .Z(n936) );
  NOR2_X1 U1032 ( .A1(KEYINPUT55), .A2(n936), .ZN(n937) );
  XOR2_X1 U1033 ( .A(KEYINPUT120), .B(n937), .Z(n938) );
  NAND2_X1 U1034 ( .A1(n938), .A2(G29), .ZN(n1015) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(G1991), .B(G25), .ZN(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n950) );
  XOR2_X1 U1038 ( .A(G2072), .B(G33), .Z(n941) );
  NAND2_X1 U1039 ( .A1(n941), .A2(G28), .ZN(n948) );
  XOR2_X1 U1040 ( .A(n942), .B(G27), .Z(n945) );
  XOR2_X1 U1041 ( .A(n943), .B(G32), .Z(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n946), .B(KEYINPUT121), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(KEYINPUT53), .B(n951), .ZN(n955) );
  XOR2_X1 U1047 ( .A(G34), .B(KEYINPUT122), .Z(n953) );
  XNOR2_X1 U1048 ( .A(G2084), .B(KEYINPUT54), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(n953), .B(n952), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G35), .B(G2090), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1053 ( .A(KEYINPUT55), .B(n958), .Z(n959) );
  NOR2_X1 U1054 ( .A1(G29), .A2(n959), .ZN(n1013) );
  XOR2_X1 U1055 ( .A(G1986), .B(G24), .Z(n963) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G22), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(G23), .B(G1976), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT125), .B(KEYINPUT58), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(n965), .B(n964), .ZN(n978) );
  XNOR2_X1 U1062 ( .A(G1966), .B(G21), .ZN(n976) );
  XOR2_X1 U1063 ( .A(G1348), .B(KEYINPUT59), .Z(n966) );
  XNOR2_X1 U1064 ( .A(G4), .B(n966), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(G19), .B(G1341), .ZN(n967) );
  NOR2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(G1956), .B(G20), .ZN(n970) );
  XNOR2_X1 U1068 ( .A(G1981), .B(G6), .ZN(n969) );
  NOR2_X1 U1069 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1071 ( .A(n973), .B(KEYINPUT60), .ZN(n974) );
  XNOR2_X1 U1072 ( .A(KEYINPUT124), .B(n974), .ZN(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(G5), .B(G1961), .ZN(n979) );
  NOR2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1077 ( .A(KEYINPUT61), .B(n981), .Z(n982) );
  NOR2_X1 U1078 ( .A1(G16), .A2(n982), .ZN(n1009) );
  XOR2_X1 U1079 ( .A(G16), .B(KEYINPUT56), .Z(n1007) );
  XNOR2_X1 U1080 ( .A(G166), .B(G1971), .ZN(n983) );
  XNOR2_X1 U1081 ( .A(n983), .B(KEYINPUT123), .ZN(n985) );
  XOR2_X1 U1082 ( .A(G171), .B(G1961), .Z(n984) );
  NOR2_X1 U1083 ( .A1(n985), .A2(n984), .ZN(n992) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G168), .ZN(n987) );
  NAND2_X1 U1085 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1086 ( .A(KEYINPUT57), .B(n988), .Z(n989) );
  NOR2_X1 U1087 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1088 ( .A1(n992), .A2(n991), .ZN(n1005) );
  XNOR2_X1 U1089 ( .A(n993), .B(G1341), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(n994), .B(G1348), .ZN(n995) );
  NOR2_X1 U1091 ( .A1(n996), .A2(n995), .ZN(n1003) );
  INV_X1 U1092 ( .A(n997), .ZN(n999) );
  NAND2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1001) );
  XNOR2_X1 U1094 ( .A(G1956), .B(G299), .ZN(n1000) );
  NOR2_X1 U1095 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1096 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(KEYINPUT126), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(G11), .A2(n1011), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(n1016), .B(KEYINPUT62), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(KEYINPUT127), .B(n1017), .ZN(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

