//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n449, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT67), .B(G108), .Z(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT68), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g023(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n449));
  AND2_X1   g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n449), .B(new_n450), .ZN(G223));
  NAND2_X1  g026(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n450), .A2(G2106), .ZN(G217));
  OR4_X1    g028(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G235), .A3(G237), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT70), .ZN(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  NAND2_X1  g035(.A1(new_n455), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  OAI211_X1 g047(.A(G137), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n473));
  INV_X1    g048(.A(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT72), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n474), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  OR2_X1    g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  AOI21_X1  g061(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n482), .A2(new_n484), .B1(G136), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n467), .A2(new_n468), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT71), .B1(new_n489), .B2(new_n466), .ZN(new_n490));
  XNOR2_X1  g065(.A(KEYINPUT3), .B(G2104), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G124), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n488), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT73), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n496), .B(new_n497), .ZN(G162));
  OAI211_X1 g073(.A(G126), .B(G2105), .C1(new_n467), .C2(new_n468), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n500), .A2(new_n502), .A3(G2104), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n506), .B1(new_n467), .B2(new_n468), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n506), .B(new_n509), .C1(new_n468), .C2(new_n467), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n504), .B1(new_n508), .B2(new_n510), .ZN(G164));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G50), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n514), .A2(new_n515), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G62), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n525), .B1(new_n518), .B2(new_n519), .ZN(new_n526));
  NAND2_X1  g101(.A1(G75), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g103(.A(G651), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n512), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n522), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G88), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n533), .A2(KEYINPUT74), .A3(new_n529), .A4(new_n517), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n531), .A2(new_n534), .ZN(G166));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  INV_X1    g112(.A(new_n516), .ZN(new_n538));
  INV_X1    g113(.A(G51), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n520), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n521), .A2(G89), .ZN(new_n542));
  NAND2_X1  g117(.A1(G63), .A2(G651), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n540), .A2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  AOI22_X1  g121(.A1(new_n520), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G651), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n516), .A2(G52), .ZN(new_n550));
  INV_X1    g125(.A(G90), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n522), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(G171));
  AOI22_X1  g128(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n548), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n516), .A2(G43), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n522), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT75), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n566));
  INV_X1    g141(.A(G91), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n522), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT76), .A4(G91), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n541), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n568), .A2(new_n569), .B1(new_n572), .B2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n516), .A2(G53), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT9), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(G299));
  NAND2_X1  g151(.A1(G171), .A2(KEYINPUT77), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n578), .B1(new_n549), .B2(new_n552), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G301));
  INV_X1    g156(.A(KEYINPUT78), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n531), .A2(new_n534), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n582), .B1(new_n531), .B2(new_n534), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(G303));
  NAND2_X1  g160(.A1(new_n532), .A2(G87), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n516), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  AOI22_X1  g164(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n548), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n516), .A2(G48), .ZN(new_n592));
  INV_X1    g167(.A(G86), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n522), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(G305));
  AOI22_X1  g171(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n548), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n516), .A2(G47), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n522), .B2(new_n600), .ZN(new_n601));
  OR3_X1    g176(.A1(new_n598), .A2(new_n601), .A3(KEYINPUT79), .ZN(new_n602));
  OAI21_X1  g177(.A(KEYINPUT79), .B1(new_n598), .B2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(G290));
  AND3_X1   g179(.A1(new_n520), .A2(new_n521), .A3(G92), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n541), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n516), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n580), .ZN(G284));
  XOR2_X1   g188(.A(G284), .B(KEYINPUT80), .Z(G321));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G299), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(new_n615), .B2(G168), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(new_n615), .B2(G168), .ZN(G280));
  INV_X1    g193(.A(new_n611), .ZN(new_n619));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G860), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT81), .ZN(G148));
  INV_X1    g197(.A(new_n559), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(new_n615), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n611), .A2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n491), .A2(new_n475), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2100), .ZN(new_n632));
  INV_X1    g207(.A(new_n494), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G123), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n635), .B1(new_n636), .B2(G2105), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(G135), .B2(new_n487), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n631), .A2(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(G2096), .ZN(new_n642));
  NAND4_X1  g217(.A1(new_n632), .A2(new_n640), .A3(new_n641), .A4(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2430), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n647), .A2(KEYINPUT14), .ZN(new_n648));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n645), .A2(new_n646), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G1341), .B(G1348), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2443), .B(G2446), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n658), .B(new_n659), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n654), .A2(new_n660), .A3(new_n656), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n665), .A2(G14), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n664), .ZN(new_n667));
  INV_X1    g242(.A(new_n663), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n666), .A2(new_n669), .ZN(G401));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT17), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT86), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n673), .B1(new_n671), .B2(KEYINPUT85), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(KEYINPUT85), .B2(new_n671), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n680), .A3(new_n675), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n674), .A2(new_n671), .A3(new_n673), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT18), .Z(new_n683));
  NAND3_X1  g258(.A1(new_n677), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(G2096), .B(G2100), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G227));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1956), .B(G2474), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT87), .ZN(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT88), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n693), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n698), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT20), .ZN(new_n701));
  INV_X1    g276(.A(G1981), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n697), .A2(new_n693), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n695), .A2(new_n696), .ZN(new_n704));
  MUX2_X1   g279(.A(new_n693), .B(new_n703), .S(new_n704), .Z(new_n705));
  NAND3_X1  g280(.A1(new_n701), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n702), .B1(new_n701), .B2(new_n705), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n691), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n701), .A2(new_n705), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G1981), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n711), .A2(G1986), .A3(new_n706), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n709), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n714), .B1(new_n709), .B2(new_n712), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n690), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n709), .A2(new_n712), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(new_n713), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n709), .A2(new_n712), .A3(new_n714), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n719), .A2(new_n689), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n717), .A2(new_n721), .ZN(G229));
  NAND3_X1  g297(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT25), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n487), .A2(G139), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT95), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n491), .A2(G127), .ZN(new_n729));
  AND2_X1   g304(.A1(G115), .A2(G2104), .ZN(new_n730));
  OAI21_X1  g305(.A(G2105), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  MUX2_X1   g307(.A(G33), .B(new_n732), .S(G29), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G2072), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT31), .B(G11), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT96), .B(G28), .Z(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(KEYINPUT30), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(KEYINPUT30), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI221_X1 g315(.A(new_n735), .B1(new_n737), .B2(new_n740), .C1(new_n639), .C2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(G16), .ZN(new_n742));
  NOR2_X1   g317(.A1(G168), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n742), .B2(G21), .ZN(new_n744));
  INV_X1    g319(.A(G1966), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n741), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G34), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n747), .A2(KEYINPUT24), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(KEYINPUT24), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n739), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G160), .B2(new_n739), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(G2084), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n742), .A2(G5), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G171), .B2(new_n742), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n752), .B1(new_n754), .B2(G1961), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(G1961), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G2084), .B2(new_n751), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n746), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n739), .A2(G32), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n633), .A2(G129), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n475), .A2(G105), .ZN(new_n761));
  NAND3_X1  g336(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT26), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n761), .B(new_n763), .C1(G141), .C2(new_n487), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n760), .A2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n759), .B1(new_n766), .B2(new_n739), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT27), .Z(new_n768));
  AOI21_X1  g343(.A(new_n758), .B1(new_n768), .B2(G1996), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n739), .A2(G27), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G164), .B2(new_n739), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT97), .B(G2078), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n745), .B2(new_n744), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n733), .A2(G2072), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n768), .A2(G1996), .ZN(new_n777));
  AND4_X1   g352(.A1(new_n734), .A2(new_n769), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(KEYINPUT98), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n739), .A2(G35), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G162), .B2(new_n739), .ZN(new_n781));
  INV_X1    g356(.A(G2090), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n619), .A2(G16), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G4), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT93), .B(G1348), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n742), .A2(G19), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n559), .B2(new_n742), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G1341), .Z(new_n792));
  NAND2_X1  g367(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n787), .A2(new_n788), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n742), .A2(G20), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT23), .Z(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G299), .B2(G16), .ZN(new_n797));
  INV_X1    g372(.A(G1956), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n739), .A2(G26), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT28), .Z(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G116), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G2105), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT94), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n487), .A2(G140), .ZN(new_n806));
  INV_X1    g381(.A(G128), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n805), .B(new_n806), .C1(new_n494), .C2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n801), .B1(new_n808), .B2(G29), .ZN(new_n809));
  INV_X1    g384(.A(G2067), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n793), .A2(new_n794), .A3(new_n799), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n779), .A2(new_n785), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n778), .A2(KEYINPUT98), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(G16), .A2(G22), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G166), .B2(G16), .ZN(new_n817));
  INV_X1    g392(.A(G1971), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT91), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n820), .ZN(new_n822));
  NOR2_X1   g397(.A1(G6), .A2(G16), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n595), .B2(G16), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT32), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n702), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n742), .A2(G23), .ZN(new_n827));
  INV_X1    g402(.A(G288), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(new_n742), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT33), .B(G1976), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n821), .A2(new_n822), .A3(new_n826), .A4(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n832), .A2(KEYINPUT34), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n834), .A2(KEYINPUT92), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n739), .A2(G25), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n633), .A2(G119), .ZN(new_n837));
  OAI21_X1  g412(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n838));
  INV_X1    g413(.A(G107), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(G2105), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G131), .B2(new_n487), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n836), .B1(new_n843), .B2(new_n739), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT35), .B(G1991), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n742), .A2(G24), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(G290), .B2(G16), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n848), .B2(new_n691), .ZN(new_n849));
  AOI211_X1 g424(.A(new_n835), .B(new_n849), .C1(new_n691), .C2(new_n848), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n832), .A2(KEYINPUT34), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n833), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n852), .A2(KEYINPUT92), .A3(new_n834), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n834), .A2(KEYINPUT92), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n815), .A2(new_n853), .A3(new_n855), .ZN(G150));
  INV_X1    g431(.A(G150), .ZN(G311));
  AOI22_X1  g432(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(new_n548), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n516), .A2(G55), .ZN(new_n860));
  INV_X1    g435(.A(G93), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n522), .B2(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(G860), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(KEYINPUT100), .ZN(new_n866));
  OR3_X1    g441(.A1(new_n859), .A2(new_n862), .A3(KEYINPUT100), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n559), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n623), .A2(new_n863), .A3(KEYINPUT100), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT38), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n611), .A2(new_n620), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n874));
  INV_X1    g449(.A(G860), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OR3_X1    g451(.A1(new_n873), .A2(KEYINPUT101), .A3(KEYINPUT39), .ZN(new_n877));
  OAI21_X1  g452(.A(KEYINPUT101), .B1(new_n873), .B2(KEYINPUT39), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n879), .A2(KEYINPUT102), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(KEYINPUT102), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n865), .B1(new_n880), .B2(new_n881), .ZN(G145));
  XNOR2_X1  g457(.A(G162), .B(G160), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT103), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(new_n639), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n883), .A2(KEYINPUT103), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(KEYINPUT103), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n886), .A2(new_n887), .B1(new_n634), .B2(new_n638), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n732), .B(new_n808), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n487), .A2(G142), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n466), .A2(G118), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n894), .B1(new_n633), .B2(G130), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n842), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n890), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n508), .A2(new_n510), .ZN(new_n898));
  INV_X1    g473(.A(new_n504), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n765), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n630), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n897), .A2(new_n902), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n889), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n903), .B(new_n904), .C1(new_n885), .C2(new_n888), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n909), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g485(.A(G290), .B(G305), .ZN(new_n911));
  XNOR2_X1  g486(.A(G166), .B(G288), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n611), .A2(G299), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n611), .A2(G299), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT41), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n870), .B(new_n625), .Z(new_n924));
  OR2_X1    g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n918), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n926), .B1(new_n925), .B2(new_n927), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n915), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n925), .A2(new_n927), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(KEYINPUT42), .ZN(new_n932));
  INV_X1    g507(.A(new_n915), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n930), .A2(new_n935), .A3(G868), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT104), .B1(new_n863), .B2(new_n615), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n930), .A2(new_n935), .A3(KEYINPUT104), .A4(G868), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(G295));
  AND2_X1   g515(.A1(new_n938), .A2(new_n939), .ZN(G331));
  AOI21_X1  g516(.A(G286), .B1(new_n577), .B2(new_n579), .ZN(new_n942));
  NOR2_X1   g517(.A1(G168), .A2(G171), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n870), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n868), .B(new_n869), .C1(new_n942), .C2(new_n943), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n920), .A2(new_n922), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n919), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n915), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n951), .B(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(KEYINPUT105), .B1(new_n950), .B2(new_n915), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n933), .A2(new_n955), .A3(new_n949), .A4(new_n947), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n954), .A2(new_n956), .A3(new_n907), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n953), .A2(KEYINPUT43), .A3(new_n957), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n954), .A2(new_n956), .A3(new_n907), .A4(new_n951), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT44), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n953), .A2(new_n957), .A3(new_n960), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n962), .A2(new_n967), .ZN(G397));
  XNOR2_X1  g543(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(G164), .B2(G1384), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n472), .A2(new_n478), .A3(G40), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n808), .B(new_n810), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n974), .B2(new_n766), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT126), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n973), .A2(G1996), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(KEYINPUT125), .B2(KEYINPUT46), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT125), .B(KEYINPUT46), .Z(new_n979));
  OAI211_X1 g554(.A(new_n976), .B(new_n978), .C1(new_n977), .C2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT47), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n843), .A2(new_n845), .ZN(new_n982));
  INV_X1    g557(.A(G1996), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n765), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n974), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n982), .B1(new_n985), .B2(new_n972), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n808), .A2(G2067), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n973), .B1(new_n988), .B2(KEYINPUT124), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n989), .B1(KEYINPUT124), .B2(new_n988), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n973), .A2(G290), .A3(G1986), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT48), .Z(new_n992));
  XOR2_X1   g567(.A(new_n842), .B(new_n845), .Z(new_n993));
  NOR2_X1   g568(.A1(new_n985), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n992), .B1(new_n973), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n981), .A2(new_n990), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n573), .A2(new_n998), .A3(new_n575), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n998), .B1(new_n573), .B2(new_n575), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1384), .ZN(new_n1002));
  INV_X1    g577(.A(new_n510), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n509), .B1(new_n491), .B2(new_n506), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1002), .B1(new_n1005), .B2(new_n504), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n971), .B1(new_n1006), .B2(new_n969), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1002), .A2(KEYINPUT45), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1008), .B(new_n1010), .C1(new_n1005), .C2(new_n504), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT108), .B1(G164), .B2(new_n1009), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT56), .B(G2072), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1007), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G40), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n471), .A2(new_n477), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(G1384), .B1(new_n898), .B2(new_n899), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1016), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n900), .A2(new_n1018), .A3(new_n1002), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT111), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1017), .A2(new_n1022), .A3(new_n1018), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1019), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1001), .B(new_n1014), .C1(new_n1024), .C2(G1956), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1017), .A2(new_n1016), .A3(new_n810), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n1020), .A3(new_n1016), .ZN(new_n1028));
  AOI211_X1 g603(.A(KEYINPUT116), .B(new_n1026), .C1(new_n788), .C2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n788), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1026), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1029), .A2(new_n1033), .A3(new_n611), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n971), .B1(new_n1006), .B2(KEYINPUT50), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1022), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1036));
  NOR4_X1   g611(.A1(G164), .A2(KEYINPUT111), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n798), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1001), .B1(new_n1039), .B2(new_n1014), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1025), .B1(new_n1034), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT61), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1025), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1042), .B1(new_n1043), .B2(new_n1040), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n970), .A2(new_n1012), .A3(new_n1016), .A4(new_n1011), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(G1996), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1008), .B1(new_n900), .B2(new_n1010), .ZN(new_n1048));
  AOI211_X1 g623(.A(KEYINPUT108), .B(new_n1009), .C1(new_n898), .C2(new_n899), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1050), .A2(KEYINPUT117), .A3(new_n983), .A4(new_n1007), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT58), .B(G1341), .Z(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1006), .B2(new_n971), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1047), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n623), .B1(new_n1055), .B2(KEYINPUT59), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1055), .A2(KEYINPUT59), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1054), .B(new_n1056), .C1(new_n1055), .C2(KEYINPUT59), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1014), .B1(new_n1024), .B2(G1956), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1001), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(KEYINPUT61), .A3(new_n1025), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1044), .A2(new_n1059), .A3(new_n1060), .A4(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT60), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1066));
  INV_X1    g641(.A(new_n788), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1067), .B1(new_n1035), .B2(new_n1020), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT116), .B1(new_n1068), .B2(new_n1026), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1031), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT60), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1066), .A2(new_n1072), .A3(new_n619), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT60), .B(new_n611), .C1(new_n1029), .C2(new_n1033), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1041), .B1(new_n1065), .B2(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n1077));
  INV_X1    g652(.A(G8), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1016), .B1(new_n1017), .B2(KEYINPUT45), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT113), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1006), .A2(new_n969), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1082), .B(new_n1016), .C1(new_n1017), .C2(KEYINPUT45), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n745), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1028), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT114), .B(G2084), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1078), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G286), .A2(G8), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(G286), .A2(KEYINPUT119), .A3(G8), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT121), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1077), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1094), .A2(KEYINPUT51), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1089), .B2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1084), .A2(new_n745), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1100), .A2(KEYINPUT122), .A3(new_n1078), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1096), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1100), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1094), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT49), .ZN(new_n1106));
  OAI21_X1  g681(.A(G1981), .B1(new_n591), .B2(new_n594), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n591), .A2(new_n594), .A3(G1981), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n595), .A2(new_n702), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(KEYINPUT49), .A3(new_n1107), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1078), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n828), .A2(G1976), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1113), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(KEYINPUT52), .ZN(new_n1117));
  INV_X1    g692(.A(G1976), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT52), .B1(G288), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n1113), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1114), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n584), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n531), .A2(new_n534), .A3(new_n582), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1122), .A2(G8), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n583), .A2(new_n584), .A3(new_n1078), .ZN(new_n1126));
  AND2_X1   g701(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1125), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1086), .A2(new_n782), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1046), .A2(new_n818), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1078), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1121), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT112), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1038), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1035), .B(KEYINPUT112), .C1(new_n1037), .C2(new_n1036), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1134), .A2(new_n782), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1078), .B1(new_n1136), .B2(new_n1130), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1132), .B1(new_n1137), .B2(new_n1128), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT53), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1046), .B2(G2078), .ZN(new_n1140));
  INV_X1    g715(.A(G1961), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1028), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1139), .A2(G2078), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1050), .A2(new_n1007), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(G171), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1080), .A2(new_n1081), .A3(new_n1083), .A4(new_n1143), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1140), .A2(new_n1147), .A3(G301), .A4(new_n1142), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1146), .A2(KEYINPUT54), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1140), .A2(new_n1147), .A3(new_n1142), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n580), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1140), .A2(G301), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT54), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1138), .A2(new_n1149), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1076), .A2(new_n1105), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1157));
  NOR2_X1   g732(.A1(G288), .A2(G1976), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT110), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1111), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1113), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1161), .B1(new_n1162), .B2(new_n1121), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT115), .B(KEYINPUT63), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1089), .A2(G168), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1138), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1165), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1167), .A2(KEYINPUT63), .A3(new_n1132), .A4(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1163), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  AND3_X1   g745(.A1(new_n1155), .A2(new_n1156), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1156), .B1(new_n1155), .B2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1138), .A2(new_n1151), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1089), .A2(new_n1098), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT122), .B1(new_n1100), .B2(new_n1078), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1174), .A2(new_n1175), .A3(new_n1097), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1176), .A2(new_n1096), .B1(new_n1094), .B2(new_n1103), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1173), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1105), .A2(KEYINPUT62), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1171), .A2(new_n1172), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g757(.A(G290), .B(new_n691), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n973), .B1(new_n994), .B2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n997), .B1(new_n1182), .B2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g760(.A1(G227), .A2(new_n464), .ZN(new_n1187));
  AOI21_X1  g761(.A(new_n1187), .B1(new_n666), .B2(new_n669), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n717), .A2(new_n721), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g765(.A1(new_n717), .A2(new_n721), .A3(new_n1188), .A4(KEYINPUT127), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g767(.A(new_n909), .B1(new_n963), .B2(new_n964), .ZN(new_n1194));
  AND2_X1   g768(.A1(new_n1193), .A2(new_n1194), .ZN(G308));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(G225));
endmodule


