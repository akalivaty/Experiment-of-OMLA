//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(new_n201), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n213), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n212), .B1(new_n219), .B2(KEYINPUT0), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(KEYINPUT0), .B2(new_n219), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT64), .Z(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  INV_X1    g0025(.A(G87), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n213), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  INV_X1    g0028(.A(G77), .ZN(new_n229));
  INV_X1    g0029(.A(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G107), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n228), .B1(new_n229), .B2(new_n230), .C1(new_n231), .C2(new_n218), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n214), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT1), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n222), .A2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n239), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  OAI21_X1  g0052(.A(KEYINPUT67), .B1(new_n214), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT67), .ZN(new_n254));
  NAND4_X1  g0054(.A1(new_n254), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n253), .A2(new_n209), .A3(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n252), .A2(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI22_X1  g0058(.A1(new_n258), .A2(new_n229), .B1(new_n210), .B2(G68), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(new_n202), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n256), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  XOR2_X1   g0063(.A(new_n263), .B(KEYINPUT11), .Z(new_n264));
  INV_X1    g0064(.A(new_n256), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G1), .B2(new_n210), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n224), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n268), .A2(new_n210), .A3(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n224), .ZN(new_n270));
  XOR2_X1   g0070(.A(new_n270), .B(KEYINPUT12), .Z(new_n271));
  INV_X1    g0071(.A(KEYINPUT70), .ZN(new_n272));
  OR3_X1    g0072(.A1(new_n267), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n272), .B1(new_n267), .B2(new_n271), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n264), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT3), .B(G33), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n276), .A2(G232), .A3(G1698), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(G226), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G97), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G238), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT66), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(G1), .B(G13), .C1(new_n252), .C2(new_n285), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G41), .A2(G45), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT66), .B1(new_n293), .B2(G1), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n291), .A2(new_n292), .A3(new_n294), .A4(G274), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT13), .B1(new_n284), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n296), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT13), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n298), .A2(new_n299), .A3(new_n283), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G200), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n275), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n301), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G190), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT71), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n303), .A2(KEYINPUT71), .A3(new_n305), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n295), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(G226), .B2(new_n288), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n276), .A2(G222), .A3(new_n278), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n276), .A2(G1698), .ZN(new_n314));
  INV_X1    g0114(.A(G223), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n313), .B1(new_n229), .B2(new_n276), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n282), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n312), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(G169), .B2(new_n318), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n260), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT68), .ZN(new_n324));
  INV_X1    g0124(.A(G58), .ZN(new_n325));
  OR3_X1    g0125(.A1(new_n325), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n322), .B1(new_n327), .B2(new_n258), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n256), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT69), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n256), .A2(new_n269), .ZN(new_n331));
  INV_X1    g0131(.A(G1), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n202), .B1(new_n332), .B2(G20), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n331), .A2(new_n333), .B1(new_n202), .B2(new_n269), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n329), .A2(KEYINPUT69), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n321), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n282), .A2(new_n287), .A3(new_n230), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n276), .A2(G232), .A3(new_n278), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n341), .B1(new_n231), .B2(new_n276), .C1(new_n314), .C2(new_n225), .ZN(new_n342));
  AOI211_X1 g0142(.A(new_n340), .B(new_n311), .C1(new_n342), .C2(new_n282), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n319), .ZN(new_n344));
  INV_X1    g0144(.A(new_n323), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT15), .B(G87), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n346), .B1(new_n258), .B2(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(new_n256), .B1(new_n229), .B2(new_n269), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n229), .B2(new_n266), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n344), .B(new_n350), .C1(G169), .C2(new_n343), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n350), .B1(new_n343), .B2(G190), .ZN(new_n352));
  INV_X1    g0152(.A(G200), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n343), .ZN(new_n354));
  AND4_X1   g0154(.A1(new_n310), .A2(new_n339), .A3(new_n351), .A4(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n301), .A2(new_n319), .ZN(new_n356));
  NOR2_X1   g0156(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n301), .A2(G169), .ZN(new_n359));
  NAND2_X1  g0159(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n359), .A2(new_n360), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n358), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n275), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT10), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT9), .B1(new_n335), .B2(new_n336), .ZN(new_n367));
  INV_X1    g0167(.A(new_n336), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT9), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n368), .A2(new_n369), .A3(new_n330), .A4(new_n334), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n353), .B1(new_n312), .B2(new_n317), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(G190), .B2(new_n318), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n366), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(new_n366), .A3(new_n373), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n355), .B(new_n365), .C1(new_n374), .C2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT18), .ZN(new_n378));
  INV_X1    g0178(.A(new_n327), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n269), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n266), .B2(new_n379), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT3), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n382), .B1(new_n383), .B2(G33), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n252), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(G33), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n210), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT7), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(new_n387), .A3(new_n210), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(G68), .A3(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n325), .A2(new_n224), .ZN(new_n394));
  OAI21_X1  g0194(.A(G20), .B1(new_n394), .B2(new_n201), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n260), .A2(G159), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(KEYINPUT16), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n224), .B1(new_n388), .B2(KEYINPUT7), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n397), .B1(new_n402), .B2(new_n392), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT75), .A3(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n390), .B1(new_n276), .B2(G20), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n386), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n210), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n410), .A3(G68), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n398), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n265), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n381), .B1(new_n405), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n288), .A2(G232), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n416), .A2(new_n295), .ZN(new_n417));
  INV_X1    g0217(.A(G226), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G1698), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(G223), .B2(G1698), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n387), .A2(new_n420), .B1(new_n252), .B2(new_n226), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n282), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n423), .A2(KEYINPUT76), .A3(G179), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT76), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n417), .A2(new_n422), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(new_n319), .ZN(new_n427));
  AOI21_X1  g0227(.A(G169), .B1(new_n417), .B2(new_n422), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n424), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g0230(.A(KEYINPUT77), .B(new_n378), .C1(new_n415), .C2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n399), .A2(new_n400), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT75), .B1(new_n403), .B2(KEYINPUT16), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n414), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n381), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n353), .B1(new_n417), .B2(new_n422), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(G190), .B2(new_n426), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n415), .A2(KEYINPUT17), .A3(new_n437), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n431), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n426), .A2(new_n425), .A3(new_n319), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT76), .B1(new_n423), .B2(G179), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n443), .B1(new_n444), .B2(new_n428), .ZN(new_n445));
  INV_X1    g0245(.A(new_n414), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n446), .B1(new_n401), .B2(new_n404), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n447), .B2(new_n381), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n378), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n445), .B(KEYINPUT18), .C1(new_n447), .C2(new_n381), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n442), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n377), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT23), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n210), .B2(G107), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n231), .A2(KEYINPUT23), .A3(G20), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G116), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(G20), .B2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n384), .A2(new_n385), .A3(new_n210), .A4(new_n386), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT22), .B1(new_n461), .B2(new_n226), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n276), .A2(new_n463), .A3(new_n210), .A4(G87), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n460), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT24), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI211_X1 g0267(.A(KEYINPUT24), .B(new_n460), .C1(new_n462), .C2(new_n464), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n256), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n269), .A2(new_n231), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n470), .B(KEYINPUT25), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n252), .A2(G1), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n256), .A2(new_n269), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n471), .B1(G107), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n332), .B(G45), .C1(new_n285), .C2(KEYINPUT5), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT79), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n286), .A2(G1), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G41), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n479), .A2(KEYINPUT79), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n285), .A2(KEYINPUT5), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(G264), .A3(new_n292), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT87), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n476), .A2(new_n477), .B1(KEYINPUT5), .B2(new_n285), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n282), .B1(new_n487), .B2(new_n482), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT87), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(G264), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n292), .A2(G274), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n487), .A3(new_n482), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n217), .A2(G1698), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n494), .B1(G250), .B2(G1698), .ZN(new_n495));
  INV_X1    g0295(.A(G294), .ZN(new_n496));
  OAI22_X1  g0296(.A1(new_n387), .A2(new_n495), .B1(new_n252), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT86), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT86), .ZN(new_n499));
  OAI221_X1 g0299(.A(new_n499), .B1(new_n252), .B2(new_n496), .C1(new_n387), .C2(new_n495), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n282), .A3(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n491), .A2(new_n319), .A3(new_n493), .A4(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(new_n486), .A3(new_n493), .A4(new_n490), .ZN(new_n503));
  INV_X1    g0303(.A(G169), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n475), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT88), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT88), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n475), .A2(new_n502), .A3(new_n508), .A4(new_n505), .ZN(new_n509));
  INV_X1    g0309(.A(new_n475), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n503), .A2(new_n353), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(G190), .B2(new_n503), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n507), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G116), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n332), .A2(new_n516), .A3(G13), .A4(G20), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT84), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n517), .B(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n473), .B2(G116), .ZN(new_n520));
  AOI21_X1  g0320(.A(G20), .B1(new_n252), .B2(G97), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n521), .A2(new_n522), .B1(G20), .B2(new_n516), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n256), .A2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT20), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n256), .A2(new_n523), .A3(KEYINPUT20), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n218), .A2(G1698), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(G257), .B2(G1698), .ZN(new_n532));
  INV_X1    g0332(.A(G303), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n387), .A2(new_n532), .B1(new_n533), .B2(new_n276), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n282), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n484), .A2(G270), .A3(new_n292), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(new_n493), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT83), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT83), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n535), .A2(new_n536), .A3(new_n539), .A4(new_n493), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(G190), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n530), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(G200), .B2(new_n541), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n538), .A2(G169), .A3(new_n529), .A4(new_n540), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT21), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n537), .A2(new_n319), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n545), .A2(new_n546), .B1(new_n529), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n541), .A2(KEYINPUT21), .A3(G169), .A4(new_n529), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n544), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n261), .A2(new_n229), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n231), .A2(KEYINPUT6), .A3(G97), .ZN(new_n553));
  XOR2_X1   g0353(.A(G97), .B(G107), .Z(new_n554));
  OAI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(KEYINPUT6), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n552), .B1(new_n555), .B2(G20), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n406), .A2(new_n410), .A3(G107), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n256), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n473), .A2(G97), .ZN(new_n560));
  INV_X1    g0360(.A(new_n269), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n561), .A2(G97), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n559), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n407), .A2(new_n386), .A3(G250), .A4(G1698), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n522), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT4), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n230), .A2(G1698), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n384), .A2(new_n385), .A3(new_n568), .A4(new_n386), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n566), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  AND2_X1   g0370(.A1(KEYINPUT4), .A2(G244), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n407), .A2(new_n386), .A3(new_n571), .A4(new_n278), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT78), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT78), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n276), .A2(new_n574), .A3(new_n278), .A4(new_n571), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n292), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n484), .A2(G257), .A3(new_n292), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n493), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n577), .A2(new_n319), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n569), .A2(new_n567), .ZN(new_n581));
  INV_X1    g0381(.A(new_n566), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n576), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n282), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n478), .A2(new_n482), .A3(new_n483), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n488), .A2(G257), .B1(new_n585), .B2(new_n492), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n504), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n564), .B1(new_n580), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n265), .B1(new_n556), .B2(new_n557), .ZN(new_n589));
  INV_X1    g0389(.A(new_n560), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n589), .A2(new_n590), .A3(new_n562), .ZN(new_n591));
  OAI21_X1  g0391(.A(G200), .B1(new_n577), .B2(new_n579), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n584), .A2(G190), .A3(new_n586), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT82), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n230), .A2(G1698), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(G238), .B2(G1698), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n459), .B1(new_n387), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n282), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n479), .A2(G274), .ZN(new_n601));
  OAI21_X1  g0401(.A(G250), .B1(new_n286), .B2(G1), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n282), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n353), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  AOI211_X1 g0405(.A(new_n542), .B(new_n603), .C1(new_n599), .C2(new_n282), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n347), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n608), .A2(new_n561), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT19), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n210), .B1(new_n280), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(G97), .ZN(new_n612));
  AND4_X1   g0412(.A1(KEYINPUT80), .A2(new_n226), .A3(new_n612), .A4(new_n231), .ZN(new_n613));
  NOR2_X1   g0413(.A1(G87), .A2(G97), .ZN(new_n614));
  AOI21_X1  g0414(.A(KEYINPUT80), .B1(new_n614), .B2(new_n231), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n611), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT81), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(new_n210), .A3(G68), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n610), .B1(new_n258), .B2(new_n612), .ZN(new_n621));
  OAI211_X1 g0421(.A(KEYINPUT81), .B(new_n611), .C1(new_n613), .C2(new_n615), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n618), .A2(new_n620), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n609), .B1(new_n623), .B2(new_n256), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n473), .A2(G87), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n607), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n600), .A2(new_n319), .A3(new_n604), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n603), .B1(new_n599), .B2(new_n282), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n627), .B1(G169), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n473), .A2(new_n608), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n624), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n596), .B1(new_n626), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n624), .A2(new_n630), .ZN(new_n633));
  INV_X1    g0433(.A(new_n629), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n607), .A2(new_n624), .A3(new_n625), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(KEYINPUT82), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n595), .B1(new_n632), .B2(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n454), .A2(new_n515), .A3(new_n551), .A4(new_n638), .ZN(G372));
  INV_X1    g0439(.A(KEYINPUT89), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n580), .B2(new_n587), .ZN(new_n641));
  OAI21_X1  g0441(.A(G169), .B1(new_n577), .B2(new_n579), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n584), .A2(G179), .A3(new_n586), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(KEYINPUT89), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n641), .A2(new_n564), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n635), .A2(new_n636), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n645), .A2(KEYINPUT26), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n588), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n626), .A2(new_n631), .A3(new_n596), .ZN(new_n649));
  AOI21_X1  g0449(.A(KEYINPUT82), .B1(new_n635), .B2(new_n636), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n647), .B1(KEYINPUT26), .B2(new_n651), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n503), .A2(G190), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n475), .B1(new_n653), .B2(new_n511), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n654), .A2(new_n595), .A3(new_n646), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n506), .A2(new_n548), .A3(new_n549), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n631), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n652), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n454), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n449), .A2(new_n451), .ZN(new_n660));
  INV_X1    g0460(.A(new_n351), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n363), .A2(new_n364), .B1(new_n306), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n440), .A2(new_n441), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT90), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n376), .B2(new_n374), .ZN(new_n666));
  INV_X1    g0466(.A(new_n374), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(KEYINPUT90), .A3(new_n375), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n338), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n659), .A2(new_n670), .ZN(G369));
  NAND3_X1  g0471(.A1(new_n332), .A2(new_n210), .A3(G13), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n530), .A2(new_n678), .ZN(new_n679));
  MUX2_X1   g0479(.A(new_n551), .B(new_n550), .S(new_n679), .Z(new_n680));
  AND2_X1   g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n510), .A2(new_n678), .ZN(new_n682));
  OAI22_X1  g0482(.A1(new_n514), .A2(new_n682), .B1(new_n506), .B2(new_n678), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n550), .A2(new_n678), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n515), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n506), .A2(new_n677), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT91), .Z(G399));
  OR3_X1    g0492(.A1(new_n216), .A2(KEYINPUT92), .A3(G41), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT92), .B1(new_n216), .B2(G41), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n613), .A2(new_n615), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n516), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n698), .A3(G1), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n207), .B2(new_n695), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n677), .B1(new_n652), .B2(new_n657), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n507), .A2(new_n509), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n655), .B1(new_n704), .B2(new_n550), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n626), .A2(new_n631), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n642), .A2(new_n643), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n591), .B1(new_n707), .B2(new_n640), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n706), .A2(new_n708), .A3(KEYINPUT26), .A4(new_n644), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n705), .B(new_n635), .C1(KEYINPUT93), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(KEYINPUT93), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT26), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(new_n651), .ZN(new_n713));
  OAI211_X1 g0513(.A(KEYINPUT29), .B(new_n678), .C1(new_n710), .C2(new_n713), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n703), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n491), .A2(new_n501), .A3(new_n628), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n577), .A2(new_n579), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n547), .A4(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n719), .A2(G179), .A3(new_n628), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(new_n503), .A3(new_n541), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT30), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n719), .A2(new_n547), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n717), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n720), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n726), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n727));
  AOI21_X1  g0527(.A(KEYINPUT31), .B1(new_n726), .B2(new_n677), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n515), .A2(new_n551), .A3(new_n638), .A4(new_n678), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n716), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n715), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n701), .B1(new_n732), .B2(G1), .ZN(G364));
  INV_X1    g0533(.A(new_n695), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n268), .A2(G20), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n332), .B1(new_n735), .B2(G45), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n681), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(G330), .B2(new_n680), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n738), .B(KEYINPUT95), .Z(new_n743));
  NAND2_X1  g0543(.A1(new_n276), .A2(new_n215), .ZN(new_n744));
  INV_X1    g0544(.A(G355), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n744), .A2(new_n745), .B1(G116), .B2(new_n215), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n247), .A2(new_n286), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n619), .A2(new_n216), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n749), .B1(new_n286), .B2(new_n208), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n746), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n209), .B1(G20), .B2(new_n504), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n743), .B1(new_n751), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n755), .ZN(new_n759));
  XOR2_X1   g0559(.A(KEYINPUT33), .B(G317), .Z(new_n760));
  NOR2_X1   g0560(.A1(new_n319), .A2(new_n353), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n210), .A2(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n319), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n762), .ZN(new_n765));
  INV_X1    g0565(.A(G311), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n760), .A2(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n210), .A2(new_n542), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n769), .A2(new_n353), .A3(G179), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n533), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n768), .A2(new_n764), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n767), .B(new_n772), .C1(G322), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n210), .B1(new_n776), .B2(G190), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n496), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n762), .A2(new_n776), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n276), .B(new_n778), .C1(G329), .C2(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n768), .A2(new_n761), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT97), .Z(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G326), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n762), .A2(new_n319), .A3(G200), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT96), .Z(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G283), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n775), .A2(new_n781), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n771), .A2(new_n226), .B1(new_n773), .B2(new_n325), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n763), .A2(new_n224), .B1(new_n765), .B2(new_n229), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n276), .B1(new_n777), .B2(new_n612), .C1(new_n782), .C2(new_n202), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G159), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n779), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n787), .A2(G107), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n793), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n759), .B1(new_n789), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n758), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n754), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n680), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n741), .A2(new_n742), .A3(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT98), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  INV_X1    g0605(.A(new_n743), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n755), .A2(new_n752), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(new_n229), .B2(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G294), .A2(new_n774), .B1(new_n780), .B2(G311), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n809), .B(new_n408), .C1(new_n231), .C2(new_n771), .ZN(new_n810));
  INV_X1    g0610(.A(new_n787), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n226), .ZN(new_n812));
  INV_X1    g0612(.A(new_n777), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n810), .B(new_n812), .C1(G97), .C2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n763), .ZN(new_n815));
  INV_X1    g0615(.A(new_n765), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G283), .A2(new_n815), .B1(new_n816), .B2(G116), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n817), .B1(new_n533), .B2(new_n782), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT99), .Z(new_n819));
  NOR2_X1   g0619(.A1(new_n811), .A2(new_n224), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n777), .A2(new_n325), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n771), .A2(new_n202), .B1(new_n779), .B2(new_n822), .ZN(new_n823));
  NOR4_X1   g0623(.A1(new_n820), .A2(new_n387), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G143), .A2(new_n774), .B1(new_n816), .B2(G159), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  INV_X1    g0626(.A(G150), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n782), .C1(new_n827), .C2(new_n763), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT34), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n814), .A2(new_n819), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n351), .A2(new_n677), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n350), .A2(new_n677), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n354), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n833), .B2(new_n351), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n808), .B1(new_n759), .B2(new_n830), .C1(new_n834), .C2(new_n753), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT100), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n702), .B2(new_n834), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n588), .A2(new_n594), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(new_n513), .A3(new_n706), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n506), .A2(new_n548), .A3(new_n549), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n635), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n706), .A2(new_n708), .A3(new_n712), .A4(new_n644), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n588), .B1(new_n632), .B2(new_n637), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(new_n712), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n678), .B(new_n834), .C1(new_n841), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(KEYINPUT100), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n837), .A2(new_n846), .B1(new_n702), .B2(new_n834), .ZN(new_n847));
  INV_X1    g0647(.A(new_n731), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n738), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n847), .A2(new_n848), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n835), .B1(new_n850), .B2(new_n851), .ZN(G384));
  OR2_X1    g0652(.A1(new_n555), .A2(KEYINPUT35), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n555), .A2(KEYINPUT35), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n853), .A2(G116), .A3(new_n211), .A4(new_n854), .ZN(new_n855));
  XOR2_X1   g0655(.A(new_n855), .B(KEYINPUT36), .Z(new_n856));
  OR3_X1    g0656(.A1(new_n207), .A2(new_n229), .A3(new_n394), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n202), .A2(G68), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n332), .B(G13), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n393), .A2(new_n398), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n265), .B1(new_n861), .B2(new_n413), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n432), .B2(new_n433), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n435), .ZN(new_n864));
  INV_X1    g0664(.A(new_n675), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n431), .A2(new_n440), .A3(new_n441), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT101), .B1(new_n415), .B2(new_n675), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT101), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n872), .B(new_n865), .C1(new_n447), .C2(new_n381), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n448), .A2(new_n438), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n864), .A2(new_n445), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n866), .A2(new_n878), .A3(new_n438), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n870), .A2(new_n881), .A3(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n874), .A2(new_n876), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT37), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(KEYINPUT103), .A3(new_n877), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n448), .A2(new_n438), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n873), .B2(new_n871), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT103), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(new_n888), .A3(new_n875), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n449), .A2(new_n451), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n873), .B(new_n871), .C1(new_n890), .C2(new_n663), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n885), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n882), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n834), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n729), .B2(new_n730), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n364), .A2(new_n677), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n306), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n365), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n363), .B1(new_n308), .B2(new_n309), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n899), .B1(new_n900), .B2(new_n897), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT40), .B1(new_n894), .B2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n902), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n877), .A2(new_n880), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n866), .B1(new_n442), .B2(new_n452), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n893), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n870), .A2(new_n881), .A3(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n904), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n903), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT105), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n729), .A2(new_n730), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n454), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(G330), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n915), .B2(new_n913), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n845), .A2(KEYINPUT100), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n658), .A2(new_n836), .A3(new_n678), .A4(new_n834), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n831), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n870), .B2(new_n881), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n882), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n901), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n660), .A2(new_n865), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT102), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n365), .A2(new_n677), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT103), .B1(new_n887), .B2(new_n875), .ZN(new_n928));
  INV_X1    g0728(.A(new_n877), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n891), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n889), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n893), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT104), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n932), .A2(new_n933), .A3(new_n934), .A4(new_n908), .ZN(new_n935));
  INV_X1    g0735(.A(new_n663), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n874), .B1(new_n936), .B2(new_n660), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n888), .B1(new_n883), .B2(KEYINPUT37), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n937), .B1(new_n938), .B2(new_n877), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT38), .B1(new_n939), .B2(new_n889), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n940), .A2(KEYINPUT39), .A3(new_n882), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT39), .B1(new_n882), .B2(new_n921), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT104), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n927), .B(new_n935), .C1(new_n941), .C2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n831), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n837), .B2(new_n846), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(new_n909), .A3(new_n901), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT102), .ZN(new_n948));
  INV_X1    g0748(.A(new_n925), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n926), .A2(new_n944), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n454), .A2(new_n715), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n952), .A2(new_n670), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n917), .A2(new_n954), .B1(new_n332), .B2(new_n735), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n917), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n860), .B1(new_n955), .B2(new_n956), .ZN(G367));
  OR3_X1    g0757(.A1(new_n683), .A2(KEYINPUT109), .A3(new_n687), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT109), .B1(new_n683), .B2(new_n687), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n958), .A2(new_n688), .A3(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(new_n681), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n732), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n838), .B1(new_n591), .B2(new_n678), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n708), .A2(new_n644), .A3(new_n677), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n688), .B2(new_n689), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n967), .A2(KEYINPUT44), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(KEYINPUT44), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT108), .ZN(new_n970));
  OR3_X1    g0770(.A1(new_n968), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT45), .ZN(new_n972));
  INV_X1    g0772(.A(new_n966), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n972), .B1(new_n690), .B2(new_n973), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n688), .A2(KEYINPUT45), .A3(new_n689), .A4(new_n966), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n969), .A2(new_n970), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n685), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n971), .A2(new_n684), .A3(new_n976), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n963), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(new_n732), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n695), .B(KEYINPUT41), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n736), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n966), .A2(new_n704), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n678), .B1(new_n984), .B2(new_n648), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n966), .A2(new_n515), .A3(new_n687), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT107), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n624), .A2(new_n625), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n677), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n706), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n631), .A2(new_n992), .A3(new_n677), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(KEYINPUT106), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT106), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT43), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n989), .A2(new_n991), .A3(new_n996), .A4(new_n999), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n989), .A2(new_n991), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n996), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1000), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n684), .A2(new_n973), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n983), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n756), .B1(new_n215), .B2(new_n347), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n243), .B2(new_n748), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n806), .A2(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G150), .A2(new_n774), .B1(new_n816), .B2(G50), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n229), .B2(new_n786), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G143), .B2(new_n784), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n777), .A2(new_n224), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n408), .B1(new_n815), .B2(G159), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n770), .A2(G58), .B1(G137), .B2(new_n780), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n770), .A2(G116), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT46), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT111), .Z(new_n1023));
  AOI22_X1  g0823(.A1(new_n1020), .A2(new_n1021), .B1(G294), .B2(new_n815), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT112), .Z(new_n1026));
  AOI22_X1  g0826(.A1(new_n784), .A2(G311), .B1(G303), .B2(new_n774), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT110), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT110), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n387), .B1(new_n231), .B2(new_n777), .ZN(new_n1030));
  INV_X1    g0830(.A(G283), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n786), .A2(new_n612), .B1(new_n765), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(G317), .C2(new_n780), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1028), .A2(new_n1029), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1019), .B1(new_n1026), .B2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT113), .Z(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT47), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1011), .B1(new_n801), .B2(new_n997), .C1(new_n1037), .C2(new_n759), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1008), .A2(new_n1038), .ZN(G387));
  OR2_X1    g0839(.A1(new_n683), .A2(new_n801), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n698), .A2(new_n744), .B1(G107), .B2(new_n215), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n749), .B1(new_n239), .B2(G45), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n697), .A2(KEYINPUT114), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n697), .A2(KEYINPUT114), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n323), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1041), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n743), .B1(new_n1049), .B2(new_n757), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n771), .A2(new_n229), .B1(new_n773), .B2(new_n202), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G68), .B2(new_n816), .ZN(new_n1052));
  XOR2_X1   g0852(.A(KEYINPUT115), .B(G150), .Z(new_n1053));
  OAI22_X1  g0853(.A1(new_n794), .A2(new_n782), .B1(new_n1053), .B2(new_n779), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n387), .B(new_n1054), .C1(new_n608), .C2(new_n813), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n379), .A2(new_n815), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n787), .A2(G97), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1052), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G311), .A2(new_n815), .B1(new_n816), .B2(G303), .ZN(new_n1059));
  INV_X1    g0859(.A(G317), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n1060), .B2(new_n773), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(KEYINPUT116), .B(G322), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1061), .B1(new_n784), .B2(new_n1062), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1063), .A2(KEYINPUT48), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n771), .A2(new_n496), .B1(new_n777), .B2(new_n1031), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1063), .B2(KEYINPUT48), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(KEYINPUT49), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n786), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1068), .A2(G116), .B1(new_n780), .B2(G326), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(new_n387), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT49), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1058), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1050), .B1(new_n1072), .B2(new_n755), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n961), .A2(new_n737), .B1(new_n1040), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n962), .A2(new_n734), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n732), .A2(new_n961), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(G393));
  INV_X1    g0877(.A(KEYINPUT117), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n979), .A2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(new_n978), .Z(new_n1080));
  OAI211_X1 g0880(.A(new_n734), .B(new_n980), .C1(new_n1080), .C2(new_n963), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n973), .A2(new_n754), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n756), .B1(new_n612), .B2(new_n215), .C1(new_n749), .C2(new_n250), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n743), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n812), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n770), .A2(G68), .B1(G143), .B2(new_n780), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n815), .A2(G50), .B1(new_n816), .B2(new_n345), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n387), .B1(new_n813), .B2(G77), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n782), .A2(new_n827), .B1(new_n773), .B2(new_n794), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT51), .Z(new_n1091));
  OAI22_X1  g0891(.A1(new_n782), .A2(new_n1060), .B1(new_n773), .B2(new_n766), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT52), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n797), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n770), .A2(G283), .B1(new_n780), .B2(new_n1062), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n276), .B1(new_n816), .B2(G294), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n815), .A2(G303), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n813), .A2(G116), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1089), .A2(new_n1091), .B1(new_n1096), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1084), .B1(new_n1102), .B2(new_n755), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1080), .A2(new_n737), .B1(new_n1082), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1081), .A2(new_n1104), .ZN(G390));
  OAI21_X1  g0905(.A(new_n935), .B1(new_n941), .B2(new_n943), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n927), .B1(new_n946), .B2(new_n901), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n896), .A2(G330), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1110), .A2(new_n923), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n901), .B(KEYINPUT118), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n833), .A2(new_n351), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n678), .B(new_n1114), .C1(new_n710), .C2(new_n713), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n945), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n927), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n894), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1109), .A2(new_n1112), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n933), .B1(new_n909), .B2(KEYINPUT39), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n932), .A2(new_n934), .A3(new_n908), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1107), .B1(new_n1124), .B2(new_n935), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1111), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1121), .A2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1128), .A2(new_n736), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1106), .A2(new_n752), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n806), .B1(new_n327), .B2(new_n807), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n1131), .A2(KEYINPUT120), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1131), .A2(KEYINPUT120), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n771), .A2(new_n1053), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT53), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n813), .A2(G159), .ZN(new_n1136));
  INV_X1    g0936(.A(G128), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n782), .A2(new_n1137), .B1(new_n763), .B2(new_n826), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n408), .B(new_n1138), .C1(G132), .C2(new_n774), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n786), .A2(new_n202), .B1(new_n765), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G125), .B2(new_n780), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1135), .A2(new_n1136), .A3(new_n1139), .A4(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n820), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n813), .A2(G77), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n782), .A2(new_n1031), .B1(new_n765), .B2(new_n612), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n276), .B(new_n1146), .C1(G87), .C2(new_n770), .ZN(new_n1147));
  OAI22_X1  g0947(.A1(new_n773), .A2(new_n516), .B1(new_n779), .B2(new_n496), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G107), .B2(new_n815), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n759), .B1(new_n1143), .B2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1132), .A2(new_n1133), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1129), .B1(new_n1130), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n454), .A2(new_n731), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n952), .A2(new_n1154), .A3(new_n670), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1111), .A2(new_n1116), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n731), .A2(KEYINPUT119), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n895), .B1(new_n731), .B2(KEYINPUT119), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1156), .B1(new_n1159), .B2(new_n1113), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n901), .B1(new_n896), .B2(G330), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n946), .B1(new_n1161), .B2(new_n1111), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1155), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1128), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1121), .A2(new_n1127), .A3(new_n1163), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n734), .A3(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1153), .A2(new_n1167), .ZN(G378));
  NAND2_X1  g0968(.A1(new_n951), .A2(KEYINPUT122), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n666), .A2(new_n668), .A3(new_n339), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n337), .A2(new_n675), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1171), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n666), .A2(new_n668), .A3(new_n339), .A4(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1175), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n896), .A2(new_n910), .A3(new_n901), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n922), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n904), .B1(new_n940), .B2(new_n882), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1181), .B2(KEYINPUT40), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1178), .B1(new_n1182), .B2(new_n716), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1178), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n912), .A2(G330), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1183), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1169), .A2(new_n1186), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n951), .A2(KEYINPUT122), .A3(new_n1183), .A4(new_n1185), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n737), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n807), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n738), .B1(G50), .B2(new_n1191), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT121), .Z(new_n1193));
  INV_X1    g0993(.A(G125), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n782), .A2(new_n1194), .B1(new_n763), .B2(new_n822), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1140), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n770), .A2(new_n1196), .B1(G137), .B2(new_n816), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n1137), .B2(new_n773), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1195), .B(new_n1198), .C1(G150), .C2(new_n813), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1068), .A2(G159), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G33), .B(G41), .C1(new_n780), .C2(G124), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n770), .A2(G77), .B1(new_n608), .B2(new_n816), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n786), .A2(new_n325), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G107), .B2(new_n774), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1206), .A2(new_n1208), .A3(new_n1016), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n387), .A2(new_n285), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n815), .A2(G97), .B1(new_n780), .B2(G283), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n516), .B2(new_n782), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT58), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1213), .A2(KEYINPUT58), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1210), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1216));
  AND4_X1   g1016(.A1(new_n1205), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1193), .B1(new_n759), .B2(new_n1217), .C1(new_n1184), .C2(new_n753), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1190), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT57), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n948), .B1(new_n947), .B2(new_n949), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1224), .A2(new_n944), .A3(new_n1183), .A4(new_n1185), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1184), .B1(new_n912), .B2(G330), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n716), .B(new_n1178), .C1(new_n903), .C2(new_n911), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n951), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1221), .B1(new_n1225), .B2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1155), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1166), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n695), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT57), .B1(new_n1189), .B2(new_n1231), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1232), .B1(new_n1233), .B2(KEYINPUT123), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1166), .A2(new_n1230), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1221), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT123), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1220), .B1(new_n1234), .B2(new_n1239), .ZN(G375));
  NAND2_X1  g1040(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1155), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n982), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1164), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1241), .A2(KEYINPUT124), .A3(new_n737), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT124), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1242), .B2(new_n736), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n743), .B1(G68), .B2(new_n1191), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n771), .A2(new_n794), .B1(new_n782), .B2(new_n822), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1207), .B(new_n1250), .C1(G150), .C2(new_n816), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n773), .A2(new_n826), .B1(new_n779), .B2(new_n1137), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n815), .B2(new_n1196), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n387), .B1(new_n813), .B2(G50), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n771), .A2(new_n612), .B1(new_n779), .B2(new_n533), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n276), .B(new_n1256), .C1(G283), .C2(new_n774), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1257), .B1(new_n347), .B2(new_n777), .C1(new_n229), .C2(new_n811), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(G116), .A2(new_n815), .B1(new_n816), .B2(G107), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n496), .B2(new_n782), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT125), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1255), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1249), .B1(new_n1262), .B2(new_n755), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1113), .B2(new_n753), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1245), .A2(new_n1246), .A3(new_n1248), .A4(new_n1264), .ZN(G381));
  NAND2_X1  g1065(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n734), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1238), .B2(new_n1237), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1233), .A2(KEYINPUT123), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1219), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(G378), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  OR4_X1    g1072(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1273));
  OR4_X1    g1073(.A1(G387), .A2(new_n1272), .A3(G381), .A4(new_n1273), .ZN(G407));
  OAI211_X1 g1074(.A(G407), .B(G213), .C1(G343), .C2(new_n1272), .ZN(G409));
  NAND2_X1  g1075(.A1(new_n676), .A2(G213), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1225), .A2(new_n1228), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n737), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1153), .A2(new_n1167), .A3(new_n1218), .A4(new_n1278), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1235), .A2(new_n1236), .A3(new_n982), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1276), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1242), .A2(KEYINPUT60), .A3(new_n1155), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n734), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1164), .A2(KEYINPUT60), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1284), .B1(new_n1243), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(G384), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1248), .A2(new_n1246), .A3(new_n1264), .ZN(new_n1288));
  OR3_X1    g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1287), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n1282), .B(new_n1291), .C1(new_n1270), .C2(new_n1271), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT127), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1292), .A2(new_n1293), .A3(KEYINPUT62), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1282), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n676), .A2(G213), .A3(G2897), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1289), .A2(new_n1290), .A3(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1281), .B1(G375), .B2(G378), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .A4(new_n1291), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1294), .A2(new_n1300), .A3(new_n1304), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1081), .A2(new_n1104), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G387), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1038), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1308), .B1(new_n983), .B2(new_n1007), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(G390), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1309), .A2(G390), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1312), .A2(KEYINPUT126), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n804), .B(G393), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1311), .B1(new_n1313), .B2(new_n1315), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1307), .A2(new_n1310), .A3(KEYINPUT126), .A4(new_n1314), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1305), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1292), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT126), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1307), .A2(new_n1322), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n1323), .A2(new_n1314), .B1(new_n1310), .B2(new_n1307), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1317), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1301), .A2(KEYINPUT63), .A3(new_n1291), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1300), .A2(new_n1321), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1319), .A2(new_n1328), .ZN(G405));
  NAND2_X1  g1129(.A1(G375), .A2(G378), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1272), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1326), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1318), .A2(new_n1272), .A3(new_n1330), .ZN(new_n1333));
  AND3_X1   g1133(.A1(new_n1332), .A2(new_n1333), .A3(new_n1291), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1291), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(G402));
endmodule


