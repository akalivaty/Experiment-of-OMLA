

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(n555), .A2(n554), .ZN(n892) );
  OR2_X1 U556 ( .A1(n771), .A2(n770), .ZN(n772) );
  AND2_X1 U557 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U558 ( .A1(n985), .A2(n730), .ZN(n736) );
  XNOR2_X1 U559 ( .A(n755), .B(KEYINPUT101), .ZN(n756) );
  XNOR2_X1 U560 ( .A(n757), .B(n756), .ZN(n758) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n747) );
  XNOR2_X1 U562 ( .A(n748), .B(n747), .ZN(n753) );
  XOR2_X1 U563 ( .A(KEYINPUT98), .B(n720), .Z(n725) );
  NAND2_X1 U564 ( .A1(n724), .A2(n725), .ZN(n766) );
  NAND2_X1 U565 ( .A1(G8), .A2(n766), .ZN(n807) );
  NOR2_X1 U566 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U567 ( .A1(G543), .A2(G651), .ZN(n660) );
  NAND2_X1 U568 ( .A1(G89), .A2(n660), .ZN(n524) );
  XOR2_X1 U569 ( .A(KEYINPUT75), .B(n524), .Z(n525) );
  XNOR2_X1 U570 ( .A(n525), .B(KEYINPUT4), .ZN(n527) );
  XOR2_X1 U571 ( .A(KEYINPUT0), .B(G543), .Z(n639) );
  INV_X1 U572 ( .A(G651), .ZN(n529) );
  NOR2_X1 U573 ( .A1(n639), .A2(n529), .ZN(n657) );
  NAND2_X1 U574 ( .A1(G76), .A2(n657), .ZN(n526) );
  NAND2_X1 U575 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U576 ( .A(n528), .B(KEYINPUT5), .ZN(n538) );
  XNOR2_X1 U577 ( .A(KEYINPUT6), .B(KEYINPUT77), .ZN(n536) );
  NOR2_X1 U578 ( .A1(G543), .A2(n529), .ZN(n530) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n530), .Z(n652) );
  NAND2_X1 U580 ( .A1(n652), .A2(G63), .ZN(n531) );
  XNOR2_X1 U581 ( .A(n531), .B(KEYINPUT76), .ZN(n534) );
  NOR2_X1 U582 ( .A1(n639), .A2(G651), .ZN(n532) );
  XNOR2_X1 U583 ( .A(KEYINPUT64), .B(n532), .ZN(n653) );
  NAND2_X1 U584 ( .A1(G51), .A2(n653), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U586 ( .A(n536), .B(n535), .ZN(n537) );
  NAND2_X1 U587 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U588 ( .A(KEYINPUT7), .B(n539), .ZN(G168) );
  XOR2_X1 U589 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U590 ( .A1(G64), .A2(n652), .ZN(n540) );
  XNOR2_X1 U591 ( .A(n540), .B(KEYINPUT68), .ZN(n543) );
  NAND2_X1 U592 ( .A1(n653), .A2(G52), .ZN(n541) );
  XOR2_X1 U593 ( .A(KEYINPUT69), .B(n541), .Z(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n548) );
  NAND2_X1 U595 ( .A1(G90), .A2(n660), .ZN(n545) );
  NAND2_X1 U596 ( .A1(G77), .A2(n657), .ZN(n544) );
  NAND2_X1 U597 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U598 ( .A(KEYINPUT9), .B(n546), .Z(n547) );
  NOR2_X1 U599 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U600 ( .A(KEYINPUT70), .B(n549), .ZN(G171) );
  INV_X1 U601 ( .A(G171), .ZN(G301) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U603 ( .A(G2105), .ZN(n554) );
  XOR2_X1 U604 ( .A(KEYINPUT65), .B(G2104), .Z(n555) );
  AND2_X1 U605 ( .A1(n554), .A2(n555), .ZN(n895) );
  NAND2_X1 U606 ( .A1(n895), .A2(G102), .ZN(n552) );
  NOR2_X1 U607 ( .A1(G2105), .A2(G2104), .ZN(n550) );
  XOR2_X2 U608 ( .A(KEYINPUT17), .B(n550), .Z(n897) );
  NAND2_X1 U609 ( .A1(n897), .A2(G138), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U611 ( .A(KEYINPUT92), .B(n553), .Z(n557) );
  NAND2_X1 U612 ( .A1(n892), .A2(G126), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n557), .A2(n556), .ZN(n560) );
  AND2_X1 U614 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U615 ( .A1(G114), .A2(n891), .ZN(n558) );
  XNOR2_X1 U616 ( .A(KEYINPUT91), .B(n558), .ZN(n559) );
  NOR2_X1 U617 ( .A1(n560), .A2(n559), .ZN(n685) );
  BUF_X1 U618 ( .A(n685), .Z(G164) );
  INV_X1 U619 ( .A(G57), .ZN(G237) );
  NAND2_X1 U620 ( .A1(n657), .A2(G75), .ZN(n561) );
  XNOR2_X1 U621 ( .A(n561), .B(KEYINPUT86), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G88), .A2(n660), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U624 ( .A(KEYINPUT87), .B(n564), .ZN(n569) );
  NAND2_X1 U625 ( .A1(G62), .A2(n652), .ZN(n566) );
  NAND2_X1 U626 ( .A1(G50), .A2(n653), .ZN(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U628 ( .A(KEYINPUT85), .B(n567), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(G303) );
  NAND2_X1 U630 ( .A1(G137), .A2(n897), .ZN(n570) );
  XNOR2_X1 U631 ( .A(n570), .B(KEYINPUT66), .ZN(n573) );
  NAND2_X1 U632 ( .A1(G101), .A2(n895), .ZN(n571) );
  XOR2_X1 U633 ( .A(KEYINPUT23), .B(n571), .Z(n572) );
  NAND2_X1 U634 ( .A1(n573), .A2(n572), .ZN(n689) );
  NAND2_X1 U635 ( .A1(G113), .A2(n891), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G125), .A2(n892), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n687) );
  NOR2_X1 U638 ( .A1(n689), .A2(n687), .ZN(G160) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U640 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U641 ( .A(G223), .ZN(n831) );
  NAND2_X1 U642 ( .A1(n831), .A2(G567), .ZN(n577) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n577), .Z(G234) );
  NAND2_X1 U644 ( .A1(G56), .A2(n652), .ZN(n578) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n578), .Z(n584) );
  NAND2_X1 U646 ( .A1(n660), .A2(G81), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n579), .B(KEYINPUT12), .ZN(n581) );
  NAND2_X1 U648 ( .A1(G68), .A2(n657), .ZN(n580) );
  NAND2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U650 ( .A(KEYINPUT13), .B(n582), .Z(n583) );
  NOR2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G43), .A2(n653), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n985) );
  INV_X1 U654 ( .A(G860), .ZN(n609) );
  OR2_X1 U655 ( .A1(n985), .A2(n609), .ZN(G153) );
  NAND2_X1 U656 ( .A1(G79), .A2(n657), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G54), .A2(n653), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n594) );
  NAND2_X1 U659 ( .A1(n660), .A2(G92), .ZN(n589) );
  XNOR2_X1 U660 ( .A(n589), .B(KEYINPUT72), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G66), .A2(n652), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U663 ( .A(n592), .B(KEYINPUT73), .Z(n593) );
  NOR2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U665 ( .A(KEYINPUT15), .B(n595), .Z(n596) );
  XNOR2_X1 U666 ( .A(KEYINPUT74), .B(n596), .ZN(n737) );
  INV_X1 U667 ( .A(n737), .ZN(n974) );
  NOR2_X1 U668 ( .A1(n974), .A2(G868), .ZN(n598) );
  INV_X1 U669 ( .A(G868), .ZN(n667) );
  NOR2_X1 U670 ( .A1(G301), .A2(n667), .ZN(n597) );
  NOR2_X1 U671 ( .A1(n598), .A2(n597), .ZN(G284) );
  NAND2_X1 U672 ( .A1(G91), .A2(n660), .ZN(n600) );
  NAND2_X1 U673 ( .A1(G78), .A2(n657), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U675 ( .A1(G65), .A2(n652), .ZN(n601) );
  XNOR2_X1 U676 ( .A(KEYINPUT71), .B(n601), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n605) );
  NAND2_X1 U678 ( .A1(G53), .A2(n653), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(G299) );
  NOR2_X1 U680 ( .A1(G286), .A2(n667), .ZN(n606) );
  XNOR2_X1 U681 ( .A(n606), .B(KEYINPUT78), .ZN(n608) );
  NOR2_X1 U682 ( .A1(G299), .A2(G868), .ZN(n607) );
  NOR2_X1 U683 ( .A1(n608), .A2(n607), .ZN(G297) );
  NAND2_X1 U684 ( .A1(n609), .A2(G559), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n610), .A2(n737), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(G868), .A2(n985), .ZN(n614) );
  NAND2_X1 U688 ( .A1(n737), .A2(G868), .ZN(n612) );
  NOR2_X1 U689 ( .A1(G559), .A2(n612), .ZN(n613) );
  NOR2_X1 U690 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U691 ( .A1(G135), .A2(n897), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G111), .A2(n891), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n892), .A2(G123), .ZN(n617) );
  XOR2_X1 U695 ( .A(KEYINPUT18), .B(n617), .Z(n618) );
  NOR2_X1 U696 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n895), .A2(G99), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n1010) );
  XNOR2_X1 U699 ( .A(G2096), .B(n1010), .ZN(n622) );
  NOR2_X1 U700 ( .A1(n622), .A2(G2100), .ZN(n623) );
  XNOR2_X1 U701 ( .A(n623), .B(KEYINPUT79), .ZN(G156) );
  NAND2_X1 U702 ( .A1(n653), .A2(G48), .ZN(n630) );
  NAND2_X1 U703 ( .A1(G86), .A2(n660), .ZN(n625) );
  NAND2_X1 U704 ( .A1(G61), .A2(n652), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n657), .A2(G73), .ZN(n626) );
  XOR2_X1 U707 ( .A(KEYINPUT2), .B(n626), .Z(n627) );
  NOR2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n631), .B(KEYINPUT84), .ZN(G305) );
  INV_X1 U711 ( .A(G303), .ZN(G166) );
  NAND2_X1 U712 ( .A1(G72), .A2(n657), .ZN(n633) );
  NAND2_X1 U713 ( .A1(G47), .A2(n653), .ZN(n632) );
  NAND2_X1 U714 ( .A1(n633), .A2(n632), .ZN(n637) );
  NAND2_X1 U715 ( .A1(G85), .A2(n660), .ZN(n635) );
  NAND2_X1 U716 ( .A1(G60), .A2(n652), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U718 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U719 ( .A(n638), .B(KEYINPUT67), .ZN(G290) );
  NAND2_X1 U720 ( .A1(G74), .A2(G651), .ZN(n641) );
  NAND2_X1 U721 ( .A1(G87), .A2(n639), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U723 ( .A1(n652), .A2(n642), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n653), .A2(G49), .ZN(n643) );
  XOR2_X1 U725 ( .A(KEYINPUT83), .B(n643), .Z(n644) );
  NAND2_X1 U726 ( .A1(n645), .A2(n644), .ZN(G288) );
  XOR2_X1 U727 ( .A(KEYINPUT19), .B(KEYINPUT88), .Z(n647) );
  INV_X1 U728 ( .A(G299), .ZN(n978) );
  XNOR2_X1 U729 ( .A(n978), .B(G166), .ZN(n646) );
  XNOR2_X1 U730 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U731 ( .A(G305), .B(n648), .ZN(n649) );
  XNOR2_X1 U732 ( .A(n649), .B(G290), .ZN(n651) );
  XOR2_X1 U733 ( .A(n985), .B(G288), .Z(n650) );
  XNOR2_X1 U734 ( .A(n651), .B(n650), .ZN(n665) );
  NAND2_X1 U735 ( .A1(G67), .A2(n652), .ZN(n655) );
  NAND2_X1 U736 ( .A1(G55), .A2(n653), .ZN(n654) );
  NAND2_X1 U737 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U738 ( .A(n656), .B(KEYINPUT81), .ZN(n659) );
  NAND2_X1 U739 ( .A1(G80), .A2(n657), .ZN(n658) );
  NAND2_X1 U740 ( .A1(n659), .A2(n658), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n660), .A2(G93), .ZN(n661) );
  XOR2_X1 U742 ( .A(KEYINPUT80), .B(n661), .Z(n662) );
  NOR2_X1 U743 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U744 ( .A(KEYINPUT82), .B(n664), .Z(n839) );
  XOR2_X1 U745 ( .A(n665), .B(n839), .Z(n862) );
  NAND2_X1 U746 ( .A1(G559), .A2(n737), .ZN(n837) );
  XNOR2_X1 U747 ( .A(n862), .B(n837), .ZN(n666) );
  NOR2_X1 U748 ( .A1(n667), .A2(n666), .ZN(n669) );
  NOR2_X1 U749 ( .A1(n839), .A2(G868), .ZN(n668) );
  NOR2_X1 U750 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XNOR2_X1 U752 ( .A(n670), .B(KEYINPUT20), .ZN(n671) );
  XNOR2_X1 U753 ( .A(n671), .B(KEYINPUT89), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n672), .A2(G2090), .ZN(n673) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U756 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U757 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U758 ( .A1(G132), .A2(G82), .ZN(n675) );
  XNOR2_X1 U759 ( .A(n675), .B(KEYINPUT22), .ZN(n676) );
  XNOR2_X1 U760 ( .A(n676), .B(KEYINPUT90), .ZN(n677) );
  NOR2_X1 U761 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U762 ( .A1(G96), .A2(n678), .ZN(n841) );
  NAND2_X1 U763 ( .A1(n841), .A2(G2106), .ZN(n682) );
  NAND2_X1 U764 ( .A1(G69), .A2(G120), .ZN(n679) );
  NOR2_X1 U765 ( .A1(G237), .A2(n679), .ZN(n680) );
  NAND2_X1 U766 ( .A1(G108), .A2(n680), .ZN(n842) );
  NAND2_X1 U767 ( .A1(n842), .A2(G567), .ZN(n681) );
  NAND2_X1 U768 ( .A1(n682), .A2(n681), .ZN(n843) );
  NAND2_X1 U769 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U770 ( .A1(n843), .A2(n683), .ZN(n836) );
  NAND2_X1 U771 ( .A1(n836), .A2(G36), .ZN(G176) );
  XOR2_X1 U772 ( .A(KEYINPUT93), .B(G1986), .Z(n684) );
  XNOR2_X1 U773 ( .A(G290), .B(n684), .ZN(n976) );
  NOR2_X1 U774 ( .A1(n685), .A2(G1384), .ZN(n724) );
  INV_X1 U775 ( .A(G40), .ZN(n686) );
  OR2_X1 U776 ( .A1(n687), .A2(n686), .ZN(n688) );
  OR2_X1 U777 ( .A1(n689), .A2(n688), .ZN(n720) );
  NOR2_X1 U778 ( .A1(n724), .A2(n720), .ZN(n826) );
  NAND2_X1 U779 ( .A1(n976), .A2(n826), .ZN(n815) );
  NAND2_X1 U780 ( .A1(G131), .A2(n897), .ZN(n691) );
  NAND2_X1 U781 ( .A1(G95), .A2(n895), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n691), .A2(n690), .ZN(n695) );
  NAND2_X1 U783 ( .A1(G107), .A2(n891), .ZN(n693) );
  NAND2_X1 U784 ( .A1(G119), .A2(n892), .ZN(n692) );
  NAND2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n694) );
  OR2_X1 U786 ( .A1(n695), .A2(n694), .ZN(n876) );
  AND2_X1 U787 ( .A1(n876), .A2(G1991), .ZN(n704) );
  NAND2_X1 U788 ( .A1(G141), .A2(n897), .ZN(n697) );
  NAND2_X1 U789 ( .A1(G117), .A2(n891), .ZN(n696) );
  NAND2_X1 U790 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n895), .A2(G105), .ZN(n698) );
  XOR2_X1 U792 ( .A(KEYINPUT38), .B(n698), .Z(n699) );
  NOR2_X1 U793 ( .A1(n700), .A2(n699), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n892), .A2(G129), .ZN(n701) );
  NAND2_X1 U795 ( .A1(n702), .A2(n701), .ZN(n874) );
  AND2_X1 U796 ( .A1(G1996), .A2(n874), .ZN(n703) );
  NOR2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n1015) );
  INV_X1 U798 ( .A(n826), .ZN(n705) );
  NOR2_X1 U799 ( .A1(n1015), .A2(n705), .ZN(n818) );
  INV_X1 U800 ( .A(n818), .ZN(n719) );
  XNOR2_X1 U801 ( .A(G2067), .B(KEYINPUT37), .ZN(n823) );
  XNOR2_X1 U802 ( .A(KEYINPUT35), .B(KEYINPUT97), .ZN(n710) );
  NAND2_X1 U803 ( .A1(n891), .A2(G116), .ZN(n706) );
  XNOR2_X1 U804 ( .A(n706), .B(KEYINPUT96), .ZN(n708) );
  NAND2_X1 U805 ( .A1(G128), .A2(n892), .ZN(n707) );
  NAND2_X1 U806 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U807 ( .A(n710), .B(n709), .ZN(n717) );
  NAND2_X1 U808 ( .A1(n897), .A2(G140), .ZN(n711) );
  XNOR2_X1 U809 ( .A(KEYINPUT95), .B(n711), .ZN(n714) );
  NAND2_X1 U810 ( .A1(n895), .A2(G104), .ZN(n712) );
  XOR2_X1 U811 ( .A(KEYINPUT94), .B(n712), .Z(n713) );
  NOR2_X1 U812 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U813 ( .A(KEYINPUT34), .B(n715), .Z(n716) );
  NOR2_X1 U814 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U815 ( .A(KEYINPUT36), .B(n718), .ZN(n905) );
  NOR2_X1 U816 ( .A1(n823), .A2(n905), .ZN(n1024) );
  NAND2_X1 U817 ( .A1(n826), .A2(n1024), .ZN(n821) );
  NAND2_X1 U818 ( .A1(n719), .A2(n821), .ZN(n813) );
  INV_X1 U819 ( .A(n766), .ZN(n749) );
  NAND2_X1 U820 ( .A1(n749), .A2(G2072), .ZN(n721) );
  XNOR2_X1 U821 ( .A(n721), .B(KEYINPUT27), .ZN(n723) );
  INV_X1 U822 ( .A(G1956), .ZN(n977) );
  NOR2_X1 U823 ( .A1(n977), .A2(n749), .ZN(n722) );
  NOR2_X1 U824 ( .A1(n723), .A2(n722), .ZN(n743) );
  NAND2_X1 U825 ( .A1(n743), .A2(n978), .ZN(n742) );
  AND2_X1 U826 ( .A1(n724), .A2(G1996), .ZN(n726) );
  XOR2_X1 U827 ( .A(n727), .B(KEYINPUT26), .Z(n729) );
  NAND2_X1 U828 ( .A1(n766), .A2(G1341), .ZN(n728) );
  NAND2_X1 U829 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U830 ( .A1(n737), .A2(n736), .ZN(n735) );
  AND2_X1 U831 ( .A1(n766), .A2(G1348), .ZN(n731) );
  XNOR2_X1 U832 ( .A(n731), .B(KEYINPUT99), .ZN(n733) );
  NAND2_X1 U833 ( .A1(n749), .A2(G2067), .ZN(n732) );
  NAND2_X1 U834 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U835 ( .A1(n735), .A2(n734), .ZN(n739) );
  OR2_X1 U836 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U837 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U838 ( .A(n740), .B(KEYINPUT100), .ZN(n741) );
  NAND2_X1 U839 ( .A1(n742), .A2(n741), .ZN(n746) );
  NOR2_X1 U840 ( .A1(n743), .A2(n978), .ZN(n744) );
  XOR2_X1 U841 ( .A(n744), .B(KEYINPUT28), .Z(n745) );
  NAND2_X1 U842 ( .A1(n746), .A2(n745), .ZN(n748) );
  XNOR2_X1 U843 ( .A(KEYINPUT25), .B(G2078), .ZN(n930) );
  NOR2_X1 U844 ( .A1(n766), .A2(n930), .ZN(n751) );
  INV_X1 U845 ( .A(G1961), .ZN(n946) );
  NOR2_X1 U846 ( .A1(n749), .A2(n946), .ZN(n750) );
  NOR2_X1 U847 ( .A1(n751), .A2(n750), .ZN(n759) );
  NAND2_X1 U848 ( .A1(G171), .A2(n759), .ZN(n752) );
  NAND2_X1 U849 ( .A1(n753), .A2(n752), .ZN(n764) );
  NOR2_X1 U850 ( .A1(G1966), .A2(n807), .ZN(n776) );
  NOR2_X1 U851 ( .A1(G2084), .A2(n766), .ZN(n777) );
  NOR2_X1 U852 ( .A1(n776), .A2(n777), .ZN(n754) );
  NAND2_X1 U853 ( .A1(G8), .A2(n754), .ZN(n757) );
  INV_X1 U854 ( .A(KEYINPUT30), .ZN(n755) );
  NOR2_X1 U855 ( .A1(G168), .A2(n758), .ZN(n761) );
  NOR2_X1 U856 ( .A1(n759), .A2(G171), .ZN(n760) );
  NOR2_X1 U857 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U858 ( .A(KEYINPUT31), .B(n762), .Z(n763) );
  NAND2_X1 U859 ( .A1(n764), .A2(n763), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n774), .A2(G286), .ZN(n765) );
  XNOR2_X1 U861 ( .A(n765), .B(KEYINPUT103), .ZN(n771) );
  NOR2_X1 U862 ( .A1(G1971), .A2(n807), .ZN(n768) );
  NOR2_X1 U863 ( .A1(G2090), .A2(n766), .ZN(n767) );
  NOR2_X1 U864 ( .A1(n768), .A2(n767), .ZN(n769) );
  AND2_X1 U865 ( .A1(G303), .A2(n769), .ZN(n770) );
  NAND2_X1 U866 ( .A1(n772), .A2(G8), .ZN(n773) );
  XNOR2_X1 U867 ( .A(n773), .B(KEYINPUT32), .ZN(n782) );
  INV_X1 U868 ( .A(n774), .ZN(n775) );
  NOR2_X1 U869 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U870 ( .A1(G8), .A2(n777), .ZN(n778) );
  NAND2_X1 U871 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U872 ( .A(KEYINPUT102), .B(n780), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n803) );
  NOR2_X1 U874 ( .A1(G1976), .A2(G288), .ZN(n980) );
  NOR2_X1 U875 ( .A1(G1971), .A2(G303), .ZN(n783) );
  NOR2_X1 U876 ( .A1(n980), .A2(n783), .ZN(n785) );
  INV_X1 U877 ( .A(KEYINPUT33), .ZN(n784) );
  AND2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U879 ( .A1(n803), .A2(n786), .ZN(n800) );
  NAND2_X1 U880 ( .A1(G288), .A2(G1976), .ZN(n787) );
  XOR2_X1 U881 ( .A(KEYINPUT104), .B(n787), .Z(n982) );
  OR2_X1 U882 ( .A1(KEYINPUT105), .A2(n982), .ZN(n788) );
  NOR2_X1 U883 ( .A1(n788), .A2(n807), .ZN(n789) );
  OR2_X1 U884 ( .A1(KEYINPUT33), .A2(n789), .ZN(n796) );
  INV_X1 U885 ( .A(KEYINPUT105), .ZN(n791) );
  NAND2_X1 U886 ( .A1(n980), .A2(KEYINPUT33), .ZN(n790) );
  NAND2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n793) );
  NAND2_X1 U888 ( .A1(n980), .A2(KEYINPUT105), .ZN(n792) );
  NAND2_X1 U889 ( .A1(n793), .A2(n792), .ZN(n794) );
  OR2_X1 U890 ( .A1(n807), .A2(n794), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n798) );
  XOR2_X1 U892 ( .A(G305), .B(G1981), .Z(n994) );
  INV_X1 U893 ( .A(n994), .ZN(n797) );
  NOR2_X1 U894 ( .A1(n798), .A2(n797), .ZN(n799) );
  AND2_X1 U895 ( .A1(n800), .A2(n799), .ZN(n811) );
  NOR2_X1 U896 ( .A1(G2090), .A2(G303), .ZN(n801) );
  NAND2_X1 U897 ( .A1(G8), .A2(n801), .ZN(n802) );
  NAND2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n804), .A2(n807), .ZN(n809) );
  NOR2_X1 U900 ( .A1(G305), .A2(G1981), .ZN(n805) );
  XOR2_X1 U901 ( .A(n805), .B(KEYINPUT24), .Z(n806) );
  OR2_X1 U902 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U905 ( .A1(n815), .A2(n814), .ZN(n829) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n874), .ZN(n1017) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n876), .ZN(n1013) );
  NOR2_X1 U909 ( .A1(n816), .A2(n1013), .ZN(n817) );
  NOR2_X1 U910 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U911 ( .A1(n1017), .A2(n819), .ZN(n820) );
  XNOR2_X1 U912 ( .A(KEYINPUT39), .B(n820), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n822), .A2(n821), .ZN(n824) );
  NAND2_X1 U914 ( .A1(n823), .A2(n905), .ZN(n1021) );
  NAND2_X1 U915 ( .A1(n824), .A2(n1021), .ZN(n825) );
  NAND2_X1 U916 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U917 ( .A(KEYINPUT106), .B(n827), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U919 ( .A(n830), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U920 ( .A1(G2106), .A2(n831), .ZN(G217) );
  NAND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n833) );
  INV_X1 U922 ( .A(G661), .ZN(n832) );
  NOR2_X1 U923 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U924 ( .A(n834), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U926 ( .A1(n836), .A2(n835), .ZN(G188) );
  XNOR2_X1 U928 ( .A(n985), .B(n837), .ZN(n838) );
  NOR2_X1 U929 ( .A1(n838), .A2(G860), .ZN(n840) );
  XOR2_X1 U930 ( .A(n840), .B(n839), .Z(G145) );
  INV_X1 U931 ( .A(G132), .ZN(G219) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G82), .ZN(G220) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  INV_X1 U937 ( .A(n843), .ZN(G319) );
  XNOR2_X1 U938 ( .A(G1961), .B(KEYINPUT41), .ZN(n853) );
  XOR2_X1 U939 ( .A(G1986), .B(G1976), .Z(n845) );
  XNOR2_X1 U940 ( .A(G1956), .B(G1971), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U942 ( .A(G1991), .B(G1981), .Z(n847) );
  XNOR2_X1 U943 ( .A(G1966), .B(G1996), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U945 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U946 ( .A(KEYINPUT110), .B(G2474), .ZN(n850) );
  XNOR2_X1 U947 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U948 ( .A(n853), .B(n852), .ZN(G229) );
  XOR2_X1 U949 ( .A(G2100), .B(G2096), .Z(n855) );
  XNOR2_X1 U950 ( .A(KEYINPUT42), .B(G2678), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U952 ( .A(KEYINPUT43), .B(G2090), .Z(n857) );
  XNOR2_X1 U953 ( .A(G2072), .B(G2067), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U955 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U956 ( .A(G2078), .B(G2084), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n861), .B(n860), .ZN(G227) );
  XOR2_X1 U958 ( .A(n862), .B(G286), .Z(n864) );
  XNOR2_X1 U959 ( .A(G301), .B(n974), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n864), .B(n863), .ZN(n865) );
  NOR2_X1 U961 ( .A1(G37), .A2(n865), .ZN(G397) );
  NAND2_X1 U962 ( .A1(G124), .A2(n892), .ZN(n866) );
  XNOR2_X1 U963 ( .A(n866), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G112), .A2(n891), .ZN(n867) );
  XOR2_X1 U965 ( .A(KEYINPUT111), .B(n867), .Z(n868) );
  NAND2_X1 U966 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U967 ( .A1(G136), .A2(n897), .ZN(n871) );
  NAND2_X1 U968 ( .A1(G100), .A2(n895), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U970 ( .A1(n873), .A2(n872), .ZN(G162) );
  XNOR2_X1 U971 ( .A(G160), .B(n874), .ZN(n875) );
  XNOR2_X1 U972 ( .A(n875), .B(n1010), .ZN(n880) );
  XOR2_X1 U973 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n878) );
  XOR2_X1 U974 ( .A(G164), .B(n876), .Z(n877) );
  XNOR2_X1 U975 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U976 ( .A(n880), .B(n879), .ZN(n890) );
  NAND2_X1 U977 ( .A1(G139), .A2(n897), .ZN(n882) );
  NAND2_X1 U978 ( .A1(G103), .A2(n895), .ZN(n881) );
  NAND2_X1 U979 ( .A1(n882), .A2(n881), .ZN(n887) );
  NAND2_X1 U980 ( .A1(G115), .A2(n891), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G127), .A2(n892), .ZN(n883) );
  NAND2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U985 ( .A(KEYINPUT113), .B(n888), .ZN(n1005) );
  XNOR2_X1 U986 ( .A(n1005), .B(G162), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n904) );
  NAND2_X1 U988 ( .A1(G118), .A2(n891), .ZN(n894) );
  NAND2_X1 U989 ( .A1(G130), .A2(n892), .ZN(n893) );
  NAND2_X1 U990 ( .A1(n894), .A2(n893), .ZN(n902) );
  NAND2_X1 U991 ( .A1(n895), .A2(G106), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n896), .B(KEYINPUT112), .ZN(n899) );
  NAND2_X1 U993 ( .A1(G142), .A2(n897), .ZN(n898) );
  NAND2_X1 U994 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U995 ( .A(n900), .B(KEYINPUT45), .Z(n901) );
  NOR2_X1 U996 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U997 ( .A(n904), .B(n903), .Z(n906) );
  XOR2_X1 U998 ( .A(n906), .B(n905), .Z(n907) );
  NOR2_X1 U999 ( .A1(G37), .A2(n907), .ZN(n908) );
  XNOR2_X1 U1000 ( .A(KEYINPUT114), .B(n908), .ZN(G395) );
  XNOR2_X1 U1001 ( .A(G2451), .B(G2427), .ZN(n918) );
  XOR2_X1 U1002 ( .A(G2430), .B(G2443), .Z(n910) );
  XNOR2_X1 U1003 ( .A(G2435), .B(G2438), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(n910), .B(n909), .ZN(n914) );
  XOR2_X1 U1005 ( .A(G2454), .B(KEYINPUT107), .Z(n912) );
  XNOR2_X1 U1006 ( .A(G1341), .B(G1348), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1008 ( .A(n914), .B(n913), .Z(n916) );
  XNOR2_X1 U1009 ( .A(G2446), .B(KEYINPUT108), .ZN(n915) );
  XNOR2_X1 U1010 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(n918), .B(n917), .ZN(n919) );
  NAND2_X1 U1012 ( .A1(n919), .A2(G14), .ZN(n925) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n925), .ZN(n922) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n920), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(G397), .A2(G395), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G96), .ZN(G221) );
  INV_X1 U1021 ( .A(G108), .ZN(G238) );
  INV_X1 U1022 ( .A(n925), .ZN(G401) );
  XOR2_X1 U1023 ( .A(KEYINPUT118), .B(G29), .Z(n945) );
  XOR2_X1 U1024 ( .A(G2084), .B(G34), .Z(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT54), .B(n926), .ZN(n941) );
  XNOR2_X1 U1026 ( .A(G2090), .B(G35), .ZN(n939) );
  XOR2_X1 U1027 ( .A(G25), .B(G1991), .Z(n927) );
  NAND2_X1 U1028 ( .A1(n927), .A2(G28), .ZN(n936) );
  XNOR2_X1 U1029 ( .A(G2072), .B(G33), .ZN(n929) );
  XNOR2_X1 U1030 ( .A(G2067), .B(G26), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n934) );
  XOR2_X1 U1032 ( .A(n930), .B(G27), .Z(n932) );
  XNOR2_X1 U1033 ( .A(G1996), .B(G32), .ZN(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(KEYINPUT53), .B(n937), .ZN(n938) );
  NOR2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(n942), .B(KEYINPUT55), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(KEYINPUT117), .B(n943), .ZN(n944) );
  NAND2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n1035) );
  XNOR2_X1 U1043 ( .A(KEYINPUT122), .B(G5), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(n947), .B(n946), .ZN(n969) );
  XOR2_X1 U1045 ( .A(G1966), .B(G21), .Z(n956) );
  XNOR2_X1 U1046 ( .A(G1986), .B(G24), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(G1971), .B(G22), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(n948), .B(KEYINPUT124), .ZN(n950) );
  XNOR2_X1 U1049 ( .A(G23), .B(G1976), .ZN(n949) );
  NOR2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1051 ( .A(KEYINPUT125), .B(n951), .ZN(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1053 ( .A(KEYINPUT58), .B(n954), .ZN(n955) );
  NAND2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n967) );
  XNOR2_X1 U1055 ( .A(G20), .B(n977), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(G1341), .B(G19), .ZN(n958) );
  XNOR2_X1 U1057 ( .A(G1981), .B(G6), .ZN(n957) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1060 ( .A(KEYINPUT59), .B(G1348), .Z(n961) );
  XNOR2_X1 U1061 ( .A(G4), .B(n961), .ZN(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1063 ( .A(KEYINPUT123), .B(n964), .ZN(n965) );
  XNOR2_X1 U1064 ( .A(KEYINPUT60), .B(n965), .ZN(n966) );
  NOR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(n970), .B(KEYINPUT126), .ZN(n971) );
  XOR2_X1 U1068 ( .A(KEYINPUT61), .B(n971), .Z(n973) );
  XNOR2_X1 U1069 ( .A(G16), .B(KEYINPUT121), .ZN(n972) );
  NAND2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n1002) );
  XNOR2_X1 U1071 ( .A(KEYINPUT56), .B(G16), .ZN(n1000) );
  XNOR2_X1 U1072 ( .A(G1348), .B(n974), .ZN(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n990) );
  XNOR2_X1 U1074 ( .A(n978), .B(n977), .ZN(n979) );
  NOR2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(G1961), .B(G301), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(G1341), .B(n985), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(KEYINPUT120), .B(n986), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1083 ( .A(G1971), .B(G303), .Z(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT119), .B(n991), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G168), .ZN(n995) );
  NAND2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(n996), .B(KEYINPUT57), .ZN(n997) );
  NAND2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1003), .B(KEYINPUT127), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(G11), .ZN(n1033) );
  XNOR2_X1 U1094 ( .A(G2072), .B(KEYINPUT116), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(n1006), .B(n1005), .ZN(n1008) );
  XOR2_X1 U1096 ( .A(G164), .B(G2078), .Z(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1098 ( .A(KEYINPUT50), .B(n1009), .Z(n1027) );
  XNOR2_X1 U1099 ( .A(G160), .B(G2084), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1020) );
  XOR2_X1 U1103 ( .A(G2090), .B(G162), .Z(n1016) );
  NOR2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(n1018), .B(KEYINPUT51), .ZN(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(KEYINPUT115), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1110 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1111 ( .A(KEYINPUT52), .B(n1028), .Z(n1029) );
  NOR2_X1 U1112 ( .A1(KEYINPUT55), .A2(n1029), .ZN(n1031) );
  INV_X1 U1113 ( .A(G29), .ZN(n1030) );
  NOR2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1115 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1116 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1036), .Z(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

