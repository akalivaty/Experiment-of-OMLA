//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT74), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G64gat), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n206), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n207), .A2(G92gat), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(G92gat), .B1(new_n207), .B2(new_n208), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G169gat), .Z(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G176gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n213), .A2(KEYINPUT23), .A3(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT25), .ZN(new_n220));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(KEYINPUT24), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n223), .B1(G183gat), .B2(G190gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n222), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G169gat), .B2(G176gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  AND2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n219), .A2(new_n220), .A3(new_n227), .A4(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G190gat), .ZN(new_n233));
  AND2_X1   g032(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT28), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT27), .B(G183gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT28), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n239), .A3(new_n233), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT26), .ZN(new_n241));
  INV_X1    g040(.A(G169gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n214), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n243), .A2(new_n230), .A3(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n237), .A2(new_n240), .A3(new_n245), .A4(new_n221), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n223), .A2(G183gat), .A3(G190gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n221), .A2(KEYINPUT24), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(new_n225), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n242), .A2(new_n214), .A3(KEYINPUT23), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n250), .A2(new_n229), .A3(new_n230), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT25), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n232), .A2(new_n246), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G226gat), .A2(G233gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n254), .B(KEYINPUT73), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT29), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n258), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G197gat), .B(G204gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT22), .ZN(new_n262));
  NAND2_X1  g061(.A1(G211gat), .A2(G218gat), .ZN(new_n263));
  OR2_X1    g062(.A1(G211gat), .A2(G218gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n265), .A2(KEYINPUT71), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(KEYINPUT71), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT22), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n263), .B1(new_n264), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(new_n261), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(new_n273), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n257), .A2(new_n260), .A3(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n271), .B(KEYINPUT72), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n276), .B1(new_n267), .B2(new_n266), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n253), .A2(new_n259), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n254), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n253), .A2(new_n258), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n212), .B1(new_n275), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT75), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT30), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n258), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n278), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n287), .A2(new_n277), .A3(new_n256), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n253), .A2(new_n258), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n255), .B1(new_n253), .B2(new_n259), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n274), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n211), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT30), .B1(new_n292), .B2(KEYINPUT75), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n288), .A2(new_n291), .A3(new_n211), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n285), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G225gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G127gat), .B(G134gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299));
  INV_X1    g098(.A(G120gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G113gat), .ZN(new_n301));
  INV_X1    g100(.A(G113gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G120gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n298), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(G134gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G127gat), .ZN(new_n307));
  INV_X1    g106(.A(G127gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G134gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT67), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT67), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n298), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT1), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT66), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n316), .B1(new_n301), .B2(new_n303), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n303), .A3(new_n316), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n314), .A2(new_n315), .A3(new_n320), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n307), .A2(new_n309), .A3(new_n312), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n312), .B1(new_n307), .B2(new_n309), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n299), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n301), .A2(new_n303), .A3(new_n316), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(new_n317), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT68), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n305), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(G141gat), .B(G148gat), .Z(new_n329));
  INV_X1    g128(.A(G155gat), .ZN(new_n330));
  INV_X1    g129(.A(G162gat), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT2), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G155gat), .B(G162gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n329), .A2(new_n334), .A3(new_n332), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n328), .A2(new_n339), .ZN(new_n340));
  AOI211_X1 g139(.A(new_n305), .B(new_n338), .C1(new_n321), .C2(new_n327), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n297), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT78), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(KEYINPUT78), .B(new_n297), .C1(new_n340), .C2(new_n341), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n347));
  INV_X1    g146(.A(new_n337), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n334), .B1(new_n329), .B2(new_n332), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT3), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT3), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n351), .A3(new_n337), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n347), .B1(new_n328), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n328), .A2(new_n339), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n297), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT4), .ZN(new_n357));
  AND3_X1   g156(.A1(new_n356), .A2(KEYINPUT77), .A3(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT77), .B1(new_n356), .B2(new_n357), .ZN(new_n359));
  OAI211_X1 g158(.A(KEYINPUT5), .B(new_n346), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n361));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n363), .B(new_n364), .Z(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n355), .A2(new_n367), .A3(KEYINPUT4), .ZN(new_n368));
  INV_X1    g167(.A(new_n305), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT68), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n315), .B1(new_n314), .B2(new_n320), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(new_n350), .A3(new_n352), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n321), .A2(new_n327), .ZN(new_n374));
  INV_X1    g173(.A(new_n347), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n374), .A2(new_n369), .A3(new_n339), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT80), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n378), .B1(new_n328), .B2(new_n339), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n368), .B(new_n373), .C1(new_n377), .C2(new_n379), .ZN(new_n380));
  OR3_X1    g179(.A1(new_n380), .A2(KEYINPUT5), .A3(new_n297), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n360), .A2(new_n366), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT6), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n366), .B1(new_n360), .B2(new_n381), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n360), .A2(new_n381), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(KEYINPUT6), .A3(new_n365), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n295), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n253), .B(new_n369), .C1(new_n371), .C2(new_n370), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n253), .B1(new_n374), .B2(new_n369), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(G227gat), .A3(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G15gat), .B(G43gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(G71gat), .ZN(new_n399));
  INV_X1    g198(.A(G99gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n395), .A2(KEYINPUT32), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT69), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n404), .B1(new_n392), .B2(new_n393), .ZN(new_n405));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n253), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n372), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n408), .A2(KEYINPUT69), .A3(new_n391), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n405), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT34), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT70), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n410), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT34), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n416), .B(new_n406), .C1(new_n392), .C2(new_n393), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n403), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n410), .A2(KEYINPUT70), .A3(KEYINPUT34), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT70), .B1(new_n410), .B2(KEYINPUT34), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n403), .B(new_n417), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n402), .B1(new_n418), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n417), .B1(new_n419), .B2(new_n420), .ZN(new_n424));
  INV_X1    g223(.A(new_n403), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n402), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n427), .A3(new_n421), .ZN(new_n428));
  INV_X1    g227(.A(new_n352), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n277), .B1(KEYINPUT29), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n273), .A2(KEYINPUT82), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT82), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n276), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n433), .A3(new_n265), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT3), .B1(new_n434), .B2(new_n259), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n430), .B1(new_n435), .B2(new_n339), .ZN(new_n436));
  INV_X1    g235(.A(G228gat), .ZN(new_n437));
  INV_X1    g236(.A(G233gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT83), .B(G22gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT3), .B1(new_n274), .B2(new_n259), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n441), .B(new_n430), .C1(new_n442), .C2(new_n339), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G78gat), .B(G106gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT31), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(G50gat), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n439), .A2(new_n443), .ZN(new_n448));
  INV_X1    g247(.A(G22gat), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n444), .B(new_n447), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n447), .B(KEYINPUT81), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n440), .B1(new_n439), .B2(new_n443), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n423), .A2(new_n428), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n202), .B1(new_n390), .B2(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n426), .A2(new_n427), .A3(new_n421), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n427), .B1(new_n426), .B2(new_n421), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n295), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n387), .A2(new_n365), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(new_n383), .A3(new_n382), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n461), .B1(new_n463), .B2(new_n388), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n460), .A2(new_n464), .A3(KEYINPUT35), .A4(new_n455), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n457), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT86), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n288), .A2(new_n291), .ZN(new_n468));
  XOR2_X1   g267(.A(KEYINPUT85), .B(KEYINPUT37), .Z(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n470), .B1(new_n471), .B2(new_n468), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT38), .B1(new_n472), .B2(new_n212), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT38), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n279), .A2(new_n280), .A3(new_n277), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n274), .B1(new_n257), .B2(new_n260), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(KEYINPUT37), .A3(new_n476), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n470), .A2(new_n474), .A3(new_n211), .A4(new_n477), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n473), .A2(new_n478), .A3(new_n282), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n463), .A2(new_n388), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n380), .A2(new_n297), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OR3_X1    g282(.A1(new_n340), .A2(new_n341), .A3(new_n297), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT39), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT39), .A4(new_n484), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n366), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT40), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n295), .B1(new_n387), .B2(new_n365), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n486), .A2(KEYINPUT40), .A3(new_n366), .A4(new_n487), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n455), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n467), .B1(new_n480), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(new_n458), .B2(new_n459), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n423), .A2(KEYINPUT36), .A3(new_n428), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n463), .A2(new_n388), .A3(new_n479), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n500), .A2(KEYINPUT86), .A3(new_n455), .A4(new_n493), .ZN(new_n501));
  INV_X1    g300(.A(new_n455), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n390), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n495), .A2(new_n499), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n466), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G230gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(new_n438), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n206), .A2(G57gat), .ZN(new_n508));
  INV_X1    g307(.A(G57gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(G64gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT9), .ZN(new_n512));
  XOR2_X1   g311(.A(G71gat), .B(G78gat), .Z(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G71gat), .ZN(new_n515));
  INV_X1    g314(.A(G78gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT9), .ZN(new_n517));
  NAND2_X1  g316(.A1(G71gat), .A2(G78gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n519), .A2(KEYINPUT93), .A3(new_n511), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT93), .B1(new_n519), .B2(new_n511), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n514), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT8), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT97), .ZN(new_n527));
  OR2_X1    g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n524), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G99gat), .B(G106gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n532), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n534), .B(new_n524), .C1(new_n529), .C2(new_n530), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n522), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT100), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n522), .ZN(new_n539));
  OAI211_X1 g338(.A(KEYINPUT98), .B(new_n524), .C1(new_n529), .C2(new_n530), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n532), .B1(new_n540), .B2(KEYINPUT99), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n528), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT97), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n528), .A3(new_n527), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n532), .A2(KEYINPUT99), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n545), .A2(new_n524), .B1(KEYINPUT98), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n539), .B1(new_n541), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n538), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT10), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n539), .B(new_n537), .C1(new_n541), .C2(new_n547), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n533), .A2(new_n535), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(new_n539), .A3(KEYINPUT10), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n507), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G120gat), .B(G148gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(new_n214), .ZN(new_n558));
  INV_X1    g357(.A(G204gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n507), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n549), .A2(new_n551), .ZN(new_n563));
  OAI211_X1 g362(.A(new_n556), .B(new_n561), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT101), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n563), .A2(new_n562), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n560), .B1(new_n566), .B2(new_n555), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(KEYINPUT101), .B(new_n560), .C1(new_n566), .C2(new_n555), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G43gat), .B(G50gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT89), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT89), .ZN(new_n574));
  INV_X1    g373(.A(G43gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(G50gat), .ZN(new_n576));
  INV_X1    g375(.A(G50gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(G43gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n574), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n573), .A2(new_n579), .A3(KEYINPUT15), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n572), .A2(KEYINPUT15), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G29gat), .ZN(new_n583));
  INV_X1    g382(.A(G36gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n584), .A3(KEYINPUT90), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT90), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(G29gat), .B2(G36gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n587), .A3(KEYINPUT14), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT14), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n586), .B(new_n589), .C1(G29gat), .C2(G36gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(G29gat), .A2(G36gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n582), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n580), .A2(new_n592), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G15gat), .B(G22gat), .ZN(new_n597));
  INV_X1    g396(.A(G1gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT16), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n597), .A2(G1gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(G8gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n600), .A2(new_n601), .A3(G8gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n596), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT91), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT17), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(KEYINPUT17), .ZN(new_n610));
  INV_X1    g409(.A(new_n595), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n592), .B1(new_n580), .B2(new_n581), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n594), .A2(new_n608), .A3(KEYINPUT17), .A4(new_n595), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n607), .B1(new_n615), .B2(new_n606), .ZN(new_n616));
  NAND2_X1  g415(.A1(G229gat), .A2(G233gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(KEYINPUT18), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT92), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n596), .B(new_n606), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n617), .B(KEYINPUT13), .Z(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT87), .B(G197gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(G113gat), .B(G141gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(KEYINPUT11), .B(G169gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n618), .A2(new_n622), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n604), .A2(new_n605), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(new_n613), .B2(new_n614), .ZN(new_n634));
  INV_X1    g433(.A(new_n617), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n634), .A2(new_n607), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(KEYINPUT18), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n623), .B(new_n631), .C1(new_n632), .C2(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n636), .A2(KEYINPUT18), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n636), .A2(KEYINPUT18), .B1(new_n620), .B2(new_n621), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n639), .B(new_n640), .C1(new_n619), .C2(new_n630), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n571), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT96), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G162gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n615), .A2(new_n533), .A3(new_n535), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n553), .A2(new_n594), .A3(new_n595), .ZN(new_n650));
  NAND3_X1  g449(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G190gat), .B(G218gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n306), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n652), .A2(new_n654), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n648), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(new_n655), .A3(new_n647), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n539), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(G183gat), .B(G211gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G231gat), .A2(G233gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT21), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n606), .B1(new_n670), .B2(new_n522), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT95), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g472(.A(G127gat), .B(G155gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n673), .A2(new_n676), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n669), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n673), .A2(new_n676), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(new_n677), .A3(new_n668), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n662), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n505), .A2(new_n644), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n386), .A2(new_n389), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT102), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g487(.A1(new_n684), .A2(new_n461), .ZN(new_n689));
  NOR2_X1   g488(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n690));
  AND2_X1   g489(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT42), .Z(new_n693));
  NAND2_X1  g492(.A1(new_n689), .A2(G8gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT103), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(G1325gat));
  AOI21_X1  g495(.A(G15gat), .B1(new_n684), .B2(new_n460), .ZN(new_n697));
  INV_X1    g496(.A(new_n499), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(G15gat), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n684), .B2(new_n699), .ZN(G1326gat));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n502), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT43), .B(G22gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  NAND2_X1  g502(.A1(new_n505), .A2(new_n662), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n680), .A2(new_n682), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n644), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(new_n583), .A3(new_n686), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n704), .A2(KEYINPUT44), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n661), .B1(new_n466), .B2(new_n504), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n707), .B1(new_n711), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n686), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G29gat), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT104), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n710), .A2(KEYINPUT104), .A3(new_n717), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1328gat));
  NAND3_X1  g521(.A1(new_n708), .A2(new_n584), .A3(new_n461), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT46), .Z(new_n724));
  NAND2_X1  g523(.A1(new_n715), .A2(new_n461), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n726), .B2(new_n584), .ZN(G1329gat));
  AOI21_X1  g526(.A(new_n575), .B1(new_n715), .B2(new_n698), .ZN(new_n728));
  INV_X1    g527(.A(new_n460), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(G43gat), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n728), .B1(new_n708), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n502), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(G50gat), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT48), .B1(new_n734), .B2(KEYINPUT105), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n708), .A2(new_n577), .A3(new_n502), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n734), .B(new_n736), .C1(KEYINPUT105), .C2(KEYINPUT48), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1331gat));
  NAND2_X1  g539(.A1(new_n683), .A2(new_n643), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n505), .A2(new_n571), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n505), .A2(KEYINPUT106), .A3(new_n571), .A4(new_n742), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n686), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(new_n509), .ZN(G1332gat));
  NOR2_X1   g549(.A1(new_n747), .A2(new_n295), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  AND2_X1   g551(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n751), .B2(new_n752), .ZN(G1333gat));
  OAI21_X1  g554(.A(new_n515), .B1(new_n747), .B2(new_n729), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n745), .A2(G71gat), .A3(new_n698), .A4(new_n746), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n757), .A2(KEYINPUT107), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n757), .A2(KEYINPUT107), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g560(.A1(new_n747), .A2(new_n455), .ZN(new_n762));
  XNOR2_X1  g561(.A(KEYINPUT108), .B(G78gat), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1335gat));
  INV_X1    g563(.A(KEYINPUT110), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n705), .A2(new_n642), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n712), .A2(KEYINPUT51), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(KEYINPUT51), .B1(new_n712), .B2(new_n766), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n505), .A2(new_n662), .A3(new_n766), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT110), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(G85gat), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n774), .A2(new_n775), .A3(new_n686), .A4(new_n571), .ZN(new_n776));
  INV_X1    g575(.A(new_n766), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n711), .B2(new_n714), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT109), .B1(new_n778), .B2(new_n571), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n712), .A2(new_n713), .ZN(new_n781));
  AOI211_X1 g580(.A(KEYINPUT44), .B(new_n661), .C1(new_n466), .C2(new_n504), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n571), .B(new_n766), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n748), .B1(new_n780), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n776), .B1(new_n787), .B2(new_n775), .ZN(G1336gat));
  NOR2_X1   g587(.A1(new_n295), .A2(G92gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n571), .A3(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791));
  OAI21_X1  g590(.A(G92gat), .B1(new_n783), .B2(new_n295), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n571), .B(new_n789), .C1(new_n767), .C2(new_n768), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n712), .A2(KEYINPUT51), .A3(new_n766), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n772), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n798), .A2(KEYINPUT111), .A3(new_n571), .A4(new_n789), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n461), .B1(new_n779), .B2(new_n785), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(G92gat), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n793), .B1(new_n802), .B2(new_n791), .ZN(G1337gat));
  AOI21_X1  g602(.A(new_n499), .B1(new_n780), .B2(new_n786), .ZN(new_n804));
  INV_X1    g603(.A(new_n774), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n460), .A2(new_n400), .A3(new_n571), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n806), .B(KEYINPUT112), .Z(new_n807));
  OAI22_X1  g606(.A1(new_n804), .A2(new_n400), .B1(new_n805), .B2(new_n807), .ZN(G1338gat));
  NOR2_X1   g607(.A1(new_n455), .A2(G106gat), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT110), .B1(new_n772), .B2(new_n797), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n768), .A2(new_n765), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n571), .B(new_n809), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT113), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n774), .A2(new_n814), .A3(new_n571), .A4(new_n809), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816));
  OAI21_X1  g615(.A(G106gat), .B1(new_n783), .B2(new_n455), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n813), .A2(new_n815), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n798), .A2(new_n571), .A3(new_n809), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n502), .B1(new_n779), .B2(new_n785), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(G106gat), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n818), .B1(new_n821), .B2(new_n816), .ZN(G1339gat));
  NAND3_X1  g621(.A1(new_n639), .A2(new_n640), .A3(new_n630), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n616), .B2(new_n617), .ZN(new_n825));
  OAI211_X1 g624(.A(KEYINPUT115), .B(new_n635), .C1(new_n634), .C2(new_n607), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n825), .B(new_n826), .C1(new_n620), .C2(new_n621), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n628), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n568), .A2(new_n569), .A3(new_n823), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n552), .A2(new_n554), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(new_n831), .A3(new_n562), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n552), .A2(new_n507), .A3(new_n554), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT54), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n560), .B(new_n832), .C1(new_n834), .C2(new_n555), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  OAI21_X1  g635(.A(KEYINPUT114), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n556), .A2(KEYINPUT54), .A3(new_n833), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n561), .B1(new_n555), .B2(new_n831), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(KEYINPUT55), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n837), .A2(new_n564), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n835), .A2(new_n836), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n642), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n829), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n661), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n662), .A2(new_n837), .A3(new_n564), .A4(new_n841), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n823), .A3(new_n828), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n842), .A2(new_n661), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851));
  INV_X1    g650(.A(new_n848), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n846), .A2(new_n849), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n706), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n683), .A2(new_n643), .A3(new_n570), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n456), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n686), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT117), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n860), .A2(new_n295), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n302), .A3(new_n642), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n859), .A2(new_n461), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(G113gat), .B1(new_n864), .B2(new_n643), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n862), .A2(new_n865), .ZN(G1340gat));
  NAND3_X1  g665(.A1(new_n861), .A2(new_n300), .A3(new_n571), .ZN(new_n867));
  OAI21_X1  g666(.A(G120gat), .B1(new_n864), .B2(new_n570), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1341gat));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n861), .A2(new_n870), .A3(new_n705), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n860), .A2(new_n705), .A3(new_n295), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT118), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n871), .A2(new_n308), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n863), .A2(G127gat), .A3(new_n705), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(G1342gat));
  NOR2_X1   g675(.A1(new_n661), .A2(G134gat), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n877), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n661), .A2(new_n461), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(G134gat), .B1(new_n859), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(KEYINPUT56), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(G1343gat));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n748), .A2(new_n698), .A3(new_n461), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n455), .B1(new_n855), .B2(new_n856), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(KEYINPUT57), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  AOI211_X1 g688(.A(new_n889), .B(new_n455), .C1(new_n855), .C2(new_n856), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(G141gat), .B1(new_n891), .B2(new_n643), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT120), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n885), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n886), .ZN(new_n895));
  INV_X1    g694(.A(new_n887), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n643), .A2(G141gat), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT119), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n892), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n894), .B(new_n901), .ZN(G1344gat));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n571), .B(new_n886), .C1(new_n888), .C2(new_n890), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n904), .A2(new_n905), .A3(G148gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n850), .A2(new_n852), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n705), .B1(new_n846), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n856), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT121), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n638), .A2(new_n641), .B1(new_n835), .B2(new_n836), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n911), .A2(new_n564), .A3(new_n837), .A4(new_n841), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n662), .B1(new_n912), .B2(new_n829), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n847), .A2(new_n848), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n706), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n916), .A3(new_n856), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n910), .A2(new_n502), .A3(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT122), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n918), .A2(new_n919), .A3(new_n889), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n918), .B2(new_n889), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n920), .A2(new_n921), .A3(new_n890), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n895), .A2(new_n570), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(G148gat), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n906), .B1(new_n925), .B2(KEYINPUT59), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n924), .A2(G148gat), .A3(new_n896), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n903), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n927), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n918), .A2(new_n889), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT122), .ZN(new_n931));
  INV_X1    g730(.A(new_n890), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n918), .A2(new_n919), .A3(new_n889), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n923), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n905), .B1(new_n935), .B2(G148gat), .ZN(new_n936));
  OAI211_X1 g735(.A(KEYINPUT123), .B(new_n929), .C1(new_n936), .C2(new_n906), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n928), .A2(new_n937), .ZN(G1345gat));
  NOR3_X1   g737(.A1(new_n891), .A2(new_n330), .A3(new_n706), .ZN(new_n939));
  AOI21_X1  g738(.A(G155gat), .B1(new_n897), .B2(new_n705), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(G1346gat));
  NOR2_X1   g740(.A1(new_n881), .A2(G162gat), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n887), .A2(new_n686), .A3(new_n499), .A4(new_n942), .ZN(new_n943));
  XOR2_X1   g742(.A(new_n943), .B(KEYINPUT124), .Z(new_n944));
  OAI21_X1  g743(.A(G162gat), .B1(new_n891), .B2(new_n661), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1347gat));
  NAND4_X1  g745(.A1(new_n857), .A2(new_n748), .A3(new_n461), .A4(new_n858), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(new_n643), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n213), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n949), .B1(new_n242), .B2(new_n948), .ZN(G1348gat));
  NOR2_X1   g749(.A1(new_n947), .A2(new_n570), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n218), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n952), .B1(new_n214), .B2(new_n951), .ZN(G1349gat));
  NOR2_X1   g752(.A1(new_n947), .A2(new_n706), .ZN(new_n954));
  MUX2_X1   g753(.A(G183gat), .B(new_n238), .S(new_n954), .Z(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT60), .ZN(G1350gat));
  XNOR2_X1  g755(.A(KEYINPUT61), .B(G190gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n947), .A2(new_n661), .ZN(new_n959));
  MUX2_X1   g758(.A(new_n957), .B(new_n958), .S(new_n959), .Z(G1351gat));
  XOR2_X1   g759(.A(KEYINPUT125), .B(G197gat), .Z(new_n961));
  NOR3_X1   g760(.A1(new_n686), .A2(new_n698), .A3(new_n295), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT126), .Z(new_n963));
  NAND2_X1  g762(.A1(new_n934), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n964), .B2(new_n643), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n887), .A2(new_n962), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n643), .A2(new_n961), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(G1352gat));
  OAI21_X1  g767(.A(G204gat), .B1(new_n964), .B2(new_n570), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n966), .A2(G204gat), .A3(new_n570), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(G1353gat));
  OR3_X1    g771(.A1(new_n966), .A2(G211gat), .A3(new_n706), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n934), .A2(new_n705), .A3(new_n962), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n974), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  NOR2_X1   g776(.A1(new_n964), .A2(KEYINPUT127), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n979), .B1(new_n934), .B2(new_n963), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n978), .A2(new_n661), .A3(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(G218gat), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n662), .A2(new_n982), .ZN(new_n983));
  OAI22_X1  g782(.A1(new_n981), .A2(new_n982), .B1(new_n966), .B2(new_n983), .ZN(G1355gat));
endmodule


