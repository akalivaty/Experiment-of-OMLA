

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737;

  XOR2_X1 U371 ( .A(KEYINPUT41), .B(n551), .Z(n639) );
  NOR2_X1 U372 ( .A1(n527), .A2(n620), .ZN(n528) );
  NOR2_X1 U373 ( .A1(n538), .A2(n537), .ZN(n539) );
  BUF_X1 U374 ( .A(n694), .Z(n699) );
  INV_X1 U375 ( .A(G953), .ZN(n723) );
  AND2_X1 U376 ( .A1(n359), .A2(n358), .ZN(n351) );
  XNOR2_X1 U377 ( .A(n489), .B(n488), .ZN(n522) );
  NOR2_X2 U378 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X2 U379 ( .A1(n390), .A2(n387), .ZN(n530) );
  XNOR2_X2 U380 ( .A(n366), .B(n704), .ZN(n685) );
  INV_X1 U381 ( .A(n592), .ZN(n620) );
  NAND2_X1 U382 ( .A1(n646), .A2(n645), .ZN(n372) );
  AND2_X1 U383 ( .A1(n381), .A2(n383), .ZN(n360) );
  XNOR2_X1 U384 ( .A(n361), .B(KEYINPUT44), .ZN(n600) );
  XNOR2_X1 U385 ( .A(n395), .B(n393), .ZN(n735) );
  NAND2_X1 U386 ( .A1(n522), .A2(n605), .ZN(n531) );
  OR2_X1 U387 ( .A1(n594), .A2(n572), .ZN(n376) );
  NOR2_X2 U388 ( .A1(n610), .A2(n352), .ZN(n551) );
  XNOR2_X1 U389 ( .A(n497), .B(n401), .ZN(n718) );
  XNOR2_X1 U390 ( .A(n402), .B(n504), .ZN(n401) );
  XNOR2_X1 U391 ( .A(n439), .B(KEYINPUT74), .ZN(n402) );
  XNOR2_X1 U392 ( .A(KEYINPUT4), .B(G137), .ZN(n439) );
  NOR2_X1 U393 ( .A1(G953), .A2(G237), .ZN(n505) );
  XNOR2_X1 U394 ( .A(n718), .B(n442), .ZN(n462) );
  XNOR2_X1 U395 ( .A(n457), .B(n456), .ZN(n481) );
  XOR2_X1 U396 ( .A(KEYINPUT3), .B(G119), .Z(n456) );
  XNOR2_X1 U397 ( .A(n455), .B(n454), .ZN(n457) );
  INV_X1 U398 ( .A(KEYINPUT90), .ZN(n454) );
  XNOR2_X1 U399 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U400 ( .A(KEYINPUT70), .B(n438), .Z(n621) );
  OR2_X1 U401 ( .A1(n689), .A2(n388), .ZN(n387) );
  AND2_X1 U402 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U403 ( .A1(G469), .A2(n389), .ZN(n388) );
  XNOR2_X1 U404 ( .A(n404), .B(G131), .ZN(n504) );
  INV_X1 U405 ( .A(KEYINPUT73), .ZN(n404) );
  XNOR2_X1 U406 ( .A(n554), .B(n416), .ZN(n555) );
  INV_X1 U407 ( .A(KEYINPUT45), .ZN(n410) );
  AND2_X2 U408 ( .A1(n368), .A2(n373), .ZN(n647) );
  INV_X1 U409 ( .A(n721), .ZN(n369) );
  XNOR2_X1 U410 ( .A(n592), .B(n520), .ZN(n572) );
  INV_X1 U411 ( .A(KEYINPUT6), .ZN(n520) );
  XNOR2_X1 U412 ( .A(n463), .B(n462), .ZN(n649) );
  XNOR2_X1 U413 ( .A(n461), .B(n460), .ZN(n463) );
  XNOR2_X1 U414 ( .A(n481), .B(n459), .ZN(n461) );
  XNOR2_X1 U415 ( .A(n515), .B(n514), .ZN(n655) );
  XOR2_X1 U416 ( .A(G140), .B(KEYINPUT93), .Z(n444) );
  XNOR2_X1 U417 ( .A(n479), .B(n476), .ZN(n414) );
  XNOR2_X1 U418 ( .A(n479), .B(n476), .ZN(n415) );
  XNOR2_X1 U419 ( .A(n379), .B(n481), .ZN(n704) );
  INV_X1 U420 ( .A(KEYINPUT39), .ZN(n491) );
  NOR2_X1 U421 ( .A1(n537), .A2(n490), .ZN(n492) );
  XNOR2_X1 U422 ( .A(n588), .B(n356), .ZN(n397) );
  INV_X1 U423 ( .A(n589), .ZN(n396) );
  XNOR2_X1 U424 ( .A(n433), .B(KEYINPUT25), .ZN(n434) );
  XNOR2_X1 U425 ( .A(n524), .B(KEYINPUT68), .ZN(n525) );
  XNOR2_X1 U426 ( .A(G116), .B(G113), .ZN(n455) );
  OR2_X1 U427 ( .A1(G237), .A2(G902), .ZN(n485) );
  INV_X1 U428 ( .A(G902), .ZN(n389) );
  NAND2_X1 U429 ( .A1(n412), .A2(G902), .ZN(n391) );
  XOR2_X1 U430 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n458) );
  AND2_X1 U431 ( .A1(n410), .A2(n599), .ZN(n382) );
  INV_X1 U432 ( .A(G134), .ZN(n441) );
  XOR2_X1 U433 ( .A(KEYINPUT99), .B(KEYINPUT11), .Z(n508) );
  XNOR2_X1 U434 ( .A(KEYINPUT100), .B(KEYINPUT12), .ZN(n507) );
  XNOR2_X1 U435 ( .A(G113), .B(G143), .ZN(n511) );
  XOR2_X1 U436 ( .A(G122), .B(G104), .Z(n512) );
  INV_X1 U437 ( .A(n504), .ZN(n403) );
  XNOR2_X1 U438 ( .A(n506), .B(KEYINPUT98), .ZN(n405) );
  XNOR2_X1 U439 ( .A(KEYINPUT17), .B(KEYINPUT89), .ZN(n471) );
  XNOR2_X1 U440 ( .A(KEYINPUT82), .B(G110), .ZN(n445) );
  XOR2_X1 U441 ( .A(G104), .B(G107), .Z(n446) );
  XOR2_X1 U442 ( .A(KEYINPUT78), .B(KEYINPUT16), .Z(n483) );
  XOR2_X1 U443 ( .A(KEYINPUT15), .B(G902), .Z(n645) );
  INV_X1 U444 ( .A(KEYINPUT2), .ZN(n373) );
  XOR2_X1 U445 ( .A(n562), .B(KEYINPUT38), .Z(n606) );
  NAND2_X1 U446 ( .A1(n374), .A2(n567), .ZN(n409) );
  AND2_X1 U447 ( .A1(n731), .A2(n399), .ZN(n398) );
  INV_X1 U448 ( .A(n683), .ZN(n399) );
  XNOR2_X1 U449 ( .A(G137), .B(G110), .ZN(n423) );
  XNOR2_X1 U450 ( .A(G119), .B(G128), .ZN(n420) );
  XOR2_X1 U451 ( .A(KEYINPUT72), .B(KEYINPUT10), .Z(n419) );
  XNOR2_X1 U452 ( .A(n472), .B(G140), .ZN(n418) );
  XNOR2_X1 U453 ( .A(KEYINPUT71), .B(KEYINPUT8), .ZN(n426) );
  XNOR2_X1 U454 ( .A(G116), .B(G107), .ZN(n494) );
  XOR2_X1 U455 ( .A(KEYINPUT9), .B(G122), .Z(n495) );
  XNOR2_X1 U456 ( .A(n407), .B(n406), .ZN(n549) );
  XNOR2_X1 U457 ( .A(n516), .B(G475), .ZN(n406) );
  OR2_X1 U458 ( .A1(n655), .A2(G902), .ZN(n407) );
  BUF_X1 U459 ( .A(n522), .Z(n562) );
  NOR2_X1 U460 ( .A1(G902), .A2(n649), .ZN(n465) );
  XNOR2_X1 U461 ( .A(n656), .B(n357), .ZN(n359) );
  NOR2_X1 U462 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U463 ( .A(n548), .B(KEYINPUT40), .ZN(n736) );
  XNOR2_X1 U464 ( .A(n394), .B(KEYINPUT86), .ZN(n393) );
  NAND2_X1 U465 ( .A1(n397), .A2(n396), .ZN(n395) );
  INV_X1 U466 ( .A(KEYINPUT35), .ZN(n394) );
  XNOR2_X1 U467 ( .A(n375), .B(KEYINPUT32), .ZN(n732) );
  NOR2_X1 U468 ( .A1(n376), .A2(n353), .ZN(n375) );
  INV_X1 U469 ( .A(KEYINPUT106), .ZN(n408) );
  INV_X1 U470 ( .A(n376), .ZN(n598) );
  XNOR2_X1 U471 ( .A(n695), .B(n362), .ZN(n698) );
  XNOR2_X1 U472 ( .A(n697), .B(n696), .ZN(n362) );
  XNOR2_X1 U473 ( .A(n692), .B(n693), .ZN(n367) );
  OR2_X1 U474 ( .A1(n550), .A2(n549), .ZN(n352) );
  XOR2_X1 U475 ( .A(KEYINPUT69), .B(G101), .Z(n477) );
  XOR2_X1 U476 ( .A(KEYINPUT105), .B(n597), .Z(n353) );
  AND2_X1 U477 ( .A1(n591), .A2(n590), .ZN(n354) );
  INV_X1 U478 ( .A(G469), .ZN(n412) );
  AND2_X1 U479 ( .A1(n367), .A2(n358), .ZN(G54) );
  XOR2_X1 U480 ( .A(n587), .B(KEYINPUT34), .Z(n356) );
  XNOR2_X1 U481 ( .A(n655), .B(KEYINPUT59), .ZN(n357) );
  XNOR2_X1 U482 ( .A(n462), .B(n448), .ZN(n689) );
  NOR2_X1 U483 ( .A1(G952), .A2(n723), .ZN(n703) );
  INV_X1 U484 ( .A(n703), .ZN(n358) );
  XNOR2_X1 U485 ( .A(n480), .B(n484), .ZN(n379) );
  OR2_X1 U486 ( .A1(n478), .A2(n414), .ZN(n380) );
  AND2_X2 U487 ( .A1(n360), .A2(n384), .ZN(n371) );
  NAND2_X1 U488 ( .A1(n601), .A2(n735), .ZN(n361) );
  XNOR2_X1 U489 ( .A(n363), .B(KEYINPUT48), .ZN(n400) );
  NOR2_X2 U490 ( .A1(n555), .A2(n556), .ZN(n363) );
  XNOR2_X1 U491 ( .A(n364), .B(n654), .ZN(G57) );
  NOR2_X2 U492 ( .A1(n652), .A2(n703), .ZN(n364) );
  INV_X1 U493 ( .A(n371), .ZN(n712) );
  NAND2_X1 U494 ( .A1(n369), .A2(n371), .ZN(n368) );
  XNOR2_X1 U495 ( .A(n365), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U496 ( .A1(n688), .A2(n703), .ZN(n365) );
  NAND2_X1 U497 ( .A1(n380), .A2(n413), .ZN(n366) );
  NAND2_X1 U498 ( .A1(n601), .A2(KEYINPUT44), .ZN(n602) );
  NOR2_X2 U499 ( .A1(n734), .A2(n732), .ZN(n601) );
  NAND2_X1 U500 ( .A1(n371), .A2(n370), .ZN(n646) );
  NOR2_X1 U501 ( .A1(n721), .A2(n373), .ZN(n370) );
  NOR2_X4 U502 ( .A1(n372), .A2(n647), .ZN(n694) );
  NAND2_X1 U503 ( .A1(n552), .A2(n374), .ZN(n671) );
  XNOR2_X2 U504 ( .A(n531), .B(KEYINPUT19), .ZN(n374) );
  XNOR2_X2 U505 ( .A(n377), .B(n408), .ZN(n734) );
  NAND2_X1 U506 ( .A1(n378), .A2(n596), .ZN(n377) );
  XNOR2_X1 U507 ( .A(n595), .B(KEYINPUT66), .ZN(n378) );
  XNOR2_X1 U508 ( .A(n475), .B(n474), .ZN(n478) );
  NAND2_X1 U509 ( .A1(n600), .A2(n382), .ZN(n381) );
  NAND2_X1 U510 ( .A1(n411), .A2(n410), .ZN(n383) );
  NAND2_X1 U511 ( .A1(n386), .A2(n385), .ZN(n384) );
  NAND2_X1 U512 ( .A1(n600), .A2(n599), .ZN(n385) );
  NOR2_X1 U513 ( .A1(n411), .A2(n410), .ZN(n386) );
  NAND2_X1 U514 ( .A1(n689), .A2(n412), .ZN(n392) );
  XNOR2_X2 U515 ( .A(n530), .B(n525), .ZN(n622) );
  XNOR2_X2 U516 ( .A(n553), .B(KEYINPUT42), .ZN(n737) );
  NAND2_X1 U517 ( .A1(n400), .A2(n398), .ZN(n721) );
  XNOR2_X2 U518 ( .A(n469), .B(n441), .ZN(n497) );
  XNOR2_X2 U519 ( .A(n440), .B(G143), .ZN(n469) );
  XNOR2_X1 U520 ( .A(n405), .B(n403), .ZN(n510) );
  XNOR2_X2 U521 ( .A(n409), .B(KEYINPUT0), .ZN(n586) );
  NAND2_X1 U522 ( .A1(n603), .A2(n354), .ZN(n411) );
  NAND2_X1 U523 ( .A1(n478), .A2(n415), .ZN(n413) );
  XNOR2_X2 U524 ( .A(n419), .B(n418), .ZN(n719) );
  XNOR2_X1 U525 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n416) );
  AND2_X1 U526 ( .A1(n493), .A2(G221), .ZN(n417) );
  XNOR2_X1 U527 ( .A(n458), .B(KEYINPUT5), .ZN(n459) );
  XNOR2_X1 U528 ( .A(n447), .B(n480), .ZN(n448) );
  XNOR2_X1 U529 ( .A(n428), .B(n417), .ZN(n429) );
  XNOR2_X1 U530 ( .A(n653), .B(KEYINPUT63), .ZN(n654) );
  XNOR2_X1 U531 ( .A(KEYINPUT120), .B(KEYINPUT60), .ZN(n657) );
  XNOR2_X1 U532 ( .A(n644), .B(n643), .ZN(G75) );
  XOR2_X2 U533 ( .A(G146), .B(G125), .Z(n472) );
  XOR2_X1 U534 ( .A(KEYINPUT23), .B(KEYINPUT94), .Z(n421) );
  XNOR2_X1 U535 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U536 ( .A(n719), .B(n422), .ZN(n430) );
  XOR2_X1 U537 ( .A(KEYINPUT95), .B(KEYINPUT75), .Z(n424) );
  XNOR2_X1 U538 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U539 ( .A(n425), .B(KEYINPUT24), .Z(n428) );
  NAND2_X1 U540 ( .A1(n723), .A2(G234), .ZN(n427) );
  XNOR2_X1 U541 ( .A(n427), .B(n426), .ZN(n493) );
  XNOR2_X1 U542 ( .A(n430), .B(n429), .ZN(n701) );
  NOR2_X1 U543 ( .A1(G902), .A2(n701), .ZN(n435) );
  INV_X1 U544 ( .A(n645), .ZN(n431) );
  NAND2_X1 U545 ( .A1(G234), .A2(n431), .ZN(n432) );
  XNOR2_X1 U546 ( .A(KEYINPUT20), .B(n432), .ZN(n436) );
  NAND2_X1 U547 ( .A1(n436), .A2(G217), .ZN(n433) );
  XNOR2_X2 U548 ( .A(n435), .B(n434), .ZN(n616) );
  NAND2_X1 U549 ( .A1(n436), .A2(G221), .ZN(n437) );
  XOR2_X1 U550 ( .A(KEYINPUT21), .B(n437), .Z(n617) );
  NAND2_X1 U551 ( .A1(n616), .A2(n617), .ZN(n438) );
  INV_X1 U552 ( .A(n621), .ZN(n449) );
  XNOR2_X2 U553 ( .A(G128), .B(KEYINPUT65), .ZN(n440) );
  XNOR2_X1 U554 ( .A(n477), .B(G146), .ZN(n442) );
  NAND2_X1 U555 ( .A1(G227), .A2(n723), .ZN(n443) );
  XNOR2_X1 U556 ( .A(n444), .B(n443), .ZN(n447) );
  XNOR2_X1 U557 ( .A(n446), .B(n445), .ZN(n480) );
  NOR2_X1 U558 ( .A1(n449), .A2(n530), .ZN(n577) );
  NOR2_X1 U559 ( .A1(G900), .A2(n723), .ZN(n450) );
  NAND2_X1 U560 ( .A1(n450), .A2(G902), .ZN(n451) );
  NAND2_X1 U561 ( .A1(G952), .A2(n723), .ZN(n564) );
  NAND2_X1 U562 ( .A1(n451), .A2(n564), .ZN(n453) );
  NAND2_X1 U563 ( .A1(G234), .A2(G237), .ZN(n452) );
  XNOR2_X1 U564 ( .A(n452), .B(KEYINPUT14), .ZN(n633) );
  NAND2_X1 U565 ( .A1(n453), .A2(n633), .ZN(n518) );
  NAND2_X1 U566 ( .A1(n505), .A2(G210), .ZN(n460) );
  INV_X1 U567 ( .A(G472), .ZN(n464) );
  XNOR2_X2 U568 ( .A(n465), .B(n464), .ZN(n592) );
  NAND2_X1 U569 ( .A1(G214), .A2(n485), .ZN(n605) );
  NAND2_X1 U570 ( .A1(n592), .A2(n605), .ZN(n466) );
  XNOR2_X1 U571 ( .A(KEYINPUT30), .B(n466), .ZN(n467) );
  NOR2_X1 U572 ( .A1(n518), .A2(n467), .ZN(n468) );
  NAND2_X1 U573 ( .A1(n577), .A2(n468), .ZN(n537) );
  XNOR2_X1 U574 ( .A(n469), .B(KEYINPUT4), .ZN(n475) );
  INV_X1 U575 ( .A(KEYINPUT18), .ZN(n470) );
  XNOR2_X1 U576 ( .A(n471), .B(n470), .ZN(n473) );
  XNOR2_X1 U577 ( .A(n473), .B(n472), .ZN(n474) );
  INV_X1 U578 ( .A(n477), .ZN(n476) );
  NAND2_X1 U579 ( .A1(G224), .A2(n723), .ZN(n479) );
  XNOR2_X1 U580 ( .A(G122), .B(KEYINPUT77), .ZN(n482) );
  XNOR2_X1 U581 ( .A(n483), .B(n482), .ZN(n484) );
  NOR2_X2 U582 ( .A1(n685), .A2(n645), .ZN(n489) );
  NAND2_X1 U583 ( .A1(G210), .A2(n485), .ZN(n487) );
  INV_X1 U584 ( .A(KEYINPUT91), .ZN(n486) );
  INV_X1 U585 ( .A(n606), .ZN(n490) );
  XNOR2_X1 U586 ( .A(n492), .B(n491), .ZN(n547) );
  XNOR2_X1 U587 ( .A(KEYINPUT103), .B(G478), .ZN(n503) );
  NAND2_X1 U588 ( .A1(n493), .A2(G217), .ZN(n501) );
  XNOR2_X1 U589 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U590 ( .A(n496), .B(KEYINPUT7), .Z(n499) );
  XNOR2_X1 U591 ( .A(n497), .B(KEYINPUT102), .ZN(n498) );
  XNOR2_X1 U592 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U593 ( .A(n501), .B(n500), .ZN(n697) );
  NOR2_X1 U594 ( .A1(G902), .A2(n697), .ZN(n502) );
  XNOR2_X1 U595 ( .A(n503), .B(n502), .ZN(n550) );
  INV_X1 U596 ( .A(n550), .ZN(n517) );
  XNOR2_X1 U597 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n516) );
  NAND2_X1 U598 ( .A1(G214), .A2(n505), .ZN(n506) );
  XNOR2_X1 U599 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U600 ( .A(n510), .B(n509), .Z(n515) );
  XNOR2_X1 U601 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U602 ( .A(n719), .B(n513), .ZN(n514) );
  NOR2_X1 U603 ( .A1(n517), .A2(n549), .ZN(n677) );
  AND2_X1 U604 ( .A1(n547), .A2(n677), .ZN(n683) );
  NAND2_X1 U605 ( .A1(n517), .A2(n549), .ZN(n672) );
  INV_X1 U606 ( .A(n672), .ZN(n674) );
  INV_X1 U607 ( .A(n616), .ZN(n596) );
  INV_X1 U608 ( .A(n617), .ZN(n568) );
  NOR2_X1 U609 ( .A1(n568), .A2(n518), .ZN(n519) );
  NAND2_X1 U610 ( .A1(n596), .A2(n519), .ZN(n527) );
  INV_X1 U611 ( .A(n572), .ZN(n583) );
  NOR2_X1 U612 ( .A1(n527), .A2(n583), .ZN(n521) );
  NAND2_X1 U613 ( .A1(n674), .A2(n521), .ZN(n557) );
  NOR2_X1 U614 ( .A1(n557), .A2(n531), .ZN(n523) );
  XNOR2_X1 U615 ( .A(KEYINPUT36), .B(n523), .ZN(n526) );
  INV_X1 U616 ( .A(KEYINPUT1), .ZN(n524) );
  NAND2_X1 U617 ( .A1(n526), .A2(n622), .ZN(n682) );
  XOR2_X1 U618 ( .A(KEYINPUT28), .B(n528), .Z(n529) );
  NOR2_X1 U619 ( .A1(n530), .A2(n529), .ZN(n552) );
  NAND2_X1 U620 ( .A1(KEYINPUT47), .A2(n671), .ZN(n532) );
  NAND2_X1 U621 ( .A1(n682), .A2(n532), .ZN(n536) );
  NOR2_X1 U622 ( .A1(KEYINPUT47), .A2(n671), .ZN(n533) );
  INV_X1 U623 ( .A(n677), .ZN(n665) );
  NAND2_X1 U624 ( .A1(n672), .A2(n665), .ZN(n541) );
  NAND2_X1 U625 ( .A1(n533), .A2(n541), .ZN(n534) );
  XNOR2_X1 U626 ( .A(KEYINPUT79), .B(n534), .ZN(n535) );
  NOR2_X1 U627 ( .A1(n536), .A2(n535), .ZN(n546) );
  NAND2_X1 U628 ( .A1(n550), .A2(n549), .ZN(n589) );
  INV_X1 U629 ( .A(n562), .ZN(n538) );
  XOR2_X1 U630 ( .A(KEYINPUT108), .B(n539), .Z(n540) );
  NOR2_X1 U631 ( .A1(n589), .A2(n540), .ZN(n669) );
  INV_X1 U632 ( .A(n541), .ZN(n609) );
  NAND2_X1 U633 ( .A1(n609), .A2(KEYINPUT47), .ZN(n542) );
  XNOR2_X1 U634 ( .A(KEYINPUT85), .B(n542), .ZN(n543) );
  NOR2_X1 U635 ( .A1(n669), .A2(n543), .ZN(n544) );
  XNOR2_X1 U636 ( .A(n544), .B(KEYINPUT84), .ZN(n545) );
  NAND2_X1 U637 ( .A1(n546), .A2(n545), .ZN(n556) );
  NAND2_X1 U638 ( .A1(n547), .A2(n674), .ZN(n548) );
  NAND2_X1 U639 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U640 ( .A1(n552), .A2(n639), .ZN(n553) );
  NAND2_X1 U641 ( .A1(n736), .A2(n737), .ZN(n554) );
  INV_X1 U642 ( .A(n557), .ZN(n558) );
  NAND2_X1 U643 ( .A1(n558), .A2(n605), .ZN(n559) );
  NOR2_X1 U644 ( .A1(n622), .A2(n559), .ZN(n560) );
  XNOR2_X1 U645 ( .A(n560), .B(KEYINPUT43), .ZN(n561) );
  NOR2_X1 U646 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U647 ( .A(KEYINPUT107), .B(n563), .ZN(n731) );
  XNOR2_X1 U648 ( .A(KEYINPUT92), .B(G898), .ZN(n709) );
  NOR2_X1 U649 ( .A1(n723), .A2(n709), .ZN(n707) );
  NAND2_X1 U650 ( .A1(n707), .A2(G902), .ZN(n565) );
  NAND2_X1 U651 ( .A1(n565), .A2(n564), .ZN(n566) );
  AND2_X1 U652 ( .A1(n566), .A2(n633), .ZN(n567) );
  OR2_X1 U653 ( .A1(n352), .A2(n568), .ZN(n569) );
  NOR2_X1 U654 ( .A1(n586), .A2(n569), .ZN(n571) );
  XNOR2_X1 U655 ( .A(KEYINPUT67), .B(KEYINPUT22), .ZN(n570) );
  XNOR2_X1 U656 ( .A(n571), .B(n570), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n598), .A2(n616), .ZN(n573) );
  NOR2_X1 U658 ( .A1(n622), .A2(n573), .ZN(n658) );
  XOR2_X1 U659 ( .A(KEYINPUT31), .B(KEYINPUT97), .Z(n575) );
  NAND2_X1 U660 ( .A1(n622), .A2(n621), .ZN(n584) );
  NOR2_X1 U661 ( .A1(n620), .A2(n584), .ZN(n627) );
  INV_X1 U662 ( .A(n586), .ZN(n576) );
  NAND2_X1 U663 ( .A1(n627), .A2(n576), .ZN(n574) );
  XNOR2_X1 U664 ( .A(n575), .B(n574), .ZN(n678) );
  NAND2_X1 U665 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U666 ( .A1(n578), .A2(n592), .ZN(n579) );
  XNOR2_X1 U667 ( .A(n579), .B(KEYINPUT96), .ZN(n660) );
  NOR2_X1 U668 ( .A1(n678), .A2(n660), .ZN(n580) );
  NOR2_X1 U669 ( .A1(n609), .A2(n580), .ZN(n581) );
  XNOR2_X1 U670 ( .A(n581), .B(KEYINPUT104), .ZN(n582) );
  NOR2_X1 U671 ( .A1(n658), .A2(n582), .ZN(n591) );
  XNOR2_X1 U672 ( .A(n585), .B(KEYINPUT33), .ZN(n613) );
  NOR2_X1 U673 ( .A1(n613), .A2(n586), .ZN(n588) );
  INV_X1 U674 ( .A(KEYINPUT76), .ZN(n587) );
  NAND2_X1 U675 ( .A1(n735), .A2(KEYINPUT87), .ZN(n590) );
  OR2_X1 U676 ( .A1(n622), .A2(n592), .ZN(n593) );
  NAND2_X1 U677 ( .A1(n622), .A2(n596), .ZN(n597) );
  INV_X1 U678 ( .A(KEYINPUT87), .ZN(n599) );
  NAND2_X1 U679 ( .A1(n602), .A2(KEYINPUT87), .ZN(n603) );
  XNOR2_X1 U680 ( .A(n647), .B(KEYINPUT83), .ZN(n604) );
  NAND2_X1 U681 ( .A1(n604), .A2(n646), .ZN(n638) );
  NOR2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U683 ( .A1(n352), .A2(n607), .ZN(n608) );
  XNOR2_X1 U684 ( .A(n608), .B(KEYINPUT116), .ZN(n612) );
  NOR2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n614) );
  NOR2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n615), .B(KEYINPUT117), .ZN(n631) );
  NOR2_X1 U689 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n618), .B(KEYINPUT49), .ZN(n619) );
  NAND2_X1 U691 ( .A1(n620), .A2(n619), .ZN(n625) );
  NOR2_X1 U692 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U693 ( .A(n623), .B(KEYINPUT50), .ZN(n624) );
  NOR2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U695 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U696 ( .A(KEYINPUT51), .B(n628), .ZN(n629) );
  NAND2_X1 U697 ( .A1(n629), .A2(n639), .ZN(n630) );
  NAND2_X1 U698 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U699 ( .A(KEYINPUT52), .B(n632), .Z(n635) );
  NAND2_X1 U700 ( .A1(G952), .A2(n633), .ZN(n634) );
  NOR2_X1 U701 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U702 ( .A1(G953), .A2(n636), .ZN(n637) );
  NAND2_X1 U703 ( .A1(n638), .A2(n637), .ZN(n642) );
  INV_X1 U704 ( .A(n639), .ZN(n640) );
  NOR2_X1 U705 ( .A1(n640), .A2(n613), .ZN(n641) );
  NOR2_X1 U706 ( .A1(n642), .A2(n641), .ZN(n644) );
  XNOR2_X1 U707 ( .A(KEYINPUT53), .B(KEYINPUT118), .ZN(n643) );
  NAND2_X1 U708 ( .A1(n694), .A2(G472), .ZN(n651) );
  XOR2_X1 U709 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n648) );
  XNOR2_X1 U710 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U711 ( .A(n651), .B(n650), .ZN(n652) );
  INV_X1 U712 ( .A(KEYINPUT88), .ZN(n653) );
  NAND2_X1 U713 ( .A1(n694), .A2(G475), .ZN(n656) );
  XNOR2_X1 U714 ( .A(n351), .B(n657), .ZN(G60) );
  XOR2_X1 U715 ( .A(G101), .B(n658), .Z(G3) );
  NAND2_X1 U716 ( .A1(n660), .A2(n674), .ZN(n659) );
  XNOR2_X1 U717 ( .A(n659), .B(G104), .ZN(G6) );
  XNOR2_X1 U718 ( .A(KEYINPUT110), .B(KEYINPUT26), .ZN(n664) );
  XOR2_X1 U719 ( .A(G107), .B(KEYINPUT27), .Z(n662) );
  NAND2_X1 U720 ( .A1(n677), .A2(n660), .ZN(n661) );
  XNOR2_X1 U721 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U722 ( .A(n664), .B(n663), .ZN(G9) );
  NOR2_X1 U723 ( .A1(n665), .A2(n671), .ZN(n667) );
  XNOR2_X1 U724 ( .A(KEYINPUT111), .B(KEYINPUT29), .ZN(n666) );
  XNOR2_X1 U725 ( .A(n667), .B(n666), .ZN(n668) );
  XOR2_X1 U726 ( .A(G128), .B(n668), .Z(G30) );
  XOR2_X1 U727 ( .A(G143), .B(n669), .Z(n670) );
  XNOR2_X1 U728 ( .A(KEYINPUT112), .B(n670), .ZN(G45) );
  NOR2_X1 U729 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U730 ( .A(G146), .B(n673), .Z(G48) );
  XOR2_X1 U731 ( .A(G113), .B(KEYINPUT113), .Z(n676) );
  NAND2_X1 U732 ( .A1(n678), .A2(n674), .ZN(n675) );
  XNOR2_X1 U733 ( .A(n676), .B(n675), .ZN(G15) );
  NAND2_X1 U734 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U735 ( .A(n679), .B(KEYINPUT114), .ZN(n680) );
  XNOR2_X1 U736 ( .A(G116), .B(n680), .ZN(G18) );
  XOR2_X1 U737 ( .A(G125), .B(KEYINPUT37), .Z(n681) );
  XNOR2_X1 U738 ( .A(n682), .B(n681), .ZN(G27) );
  XOR2_X1 U739 ( .A(G134), .B(n683), .Z(G36) );
  NAND2_X1 U740 ( .A1(n694), .A2(G210), .ZN(n687) );
  XOR2_X1 U741 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n684) );
  XNOR2_X1 U742 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U743 ( .A(n687), .B(n686), .ZN(n688) );
  XOR2_X1 U744 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n691) );
  XNOR2_X1 U745 ( .A(n689), .B(KEYINPUT119), .ZN(n690) );
  XNOR2_X1 U746 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U747 ( .A1(n699), .A2(G469), .ZN(n692) );
  XOR2_X1 U748 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n696) );
  NAND2_X1 U749 ( .A1(n699), .A2(G478), .ZN(n695) );
  NOR2_X1 U750 ( .A1(n703), .A2(n698), .ZN(G63) );
  NAND2_X1 U751 ( .A1(G217), .A2(n699), .ZN(n700) );
  XNOR2_X1 U752 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U753 ( .A1(n703), .A2(n702), .ZN(G66) );
  XNOR2_X1 U754 ( .A(G101), .B(n704), .ZN(n705) );
  XNOR2_X1 U755 ( .A(n705), .B(KEYINPUT125), .ZN(n706) );
  NOR2_X1 U756 ( .A1(n707), .A2(n706), .ZN(n717) );
  NAND2_X1 U757 ( .A1(G953), .A2(G224), .ZN(n708) );
  XNOR2_X1 U758 ( .A(n708), .B(KEYINPUT61), .ZN(n710) );
  NAND2_X1 U759 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U760 ( .A(KEYINPUT123), .B(n711), .ZN(n715) );
  NOR2_X1 U761 ( .A1(G953), .A2(n712), .ZN(n713) );
  XNOR2_X1 U762 ( .A(KEYINPUT124), .B(n713), .ZN(n714) );
  NOR2_X1 U763 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U764 ( .A(n717), .B(n716), .Z(G69) );
  XNOR2_X1 U765 ( .A(n718), .B(KEYINPUT93), .ZN(n720) );
  XNOR2_X1 U766 ( .A(n720), .B(n719), .ZN(n725) );
  XNOR2_X1 U767 ( .A(n725), .B(KEYINPUT126), .ZN(n722) );
  XNOR2_X1 U768 ( .A(n722), .B(n721), .ZN(n724) );
  NAND2_X1 U769 ( .A1(n724), .A2(n723), .ZN(n729) );
  XNOR2_X1 U770 ( .A(G227), .B(n725), .ZN(n726) );
  NAND2_X1 U771 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U772 ( .A1(n727), .A2(G953), .ZN(n728) );
  NAND2_X1 U773 ( .A1(n729), .A2(n728), .ZN(G72) );
  XOR2_X1 U774 ( .A(G140), .B(KEYINPUT115), .Z(n730) );
  XNOR2_X1 U775 ( .A(n731), .B(n730), .ZN(G42) );
  XNOR2_X1 U776 ( .A(G119), .B(KEYINPUT127), .ZN(n733) );
  XNOR2_X1 U777 ( .A(n733), .B(n732), .ZN(G21) );
  XOR2_X1 U778 ( .A(n734), .B(G110), .Z(G12) );
  XNOR2_X1 U779 ( .A(n735), .B(G122), .ZN(G24) );
  XNOR2_X1 U780 ( .A(G131), .B(n736), .ZN(G33) );
  XNOR2_X1 U781 ( .A(G137), .B(n737), .ZN(G39) );
endmodule

