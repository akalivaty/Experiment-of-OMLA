//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n441, new_n445, new_n448, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n570, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT67), .B(G57), .Z(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT68), .Z(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT69), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT70), .Z(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g029(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT2), .ZN(new_n456));
  NAND4_X1  g031(.A1(new_n441), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT71), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  NAND2_X1  g035(.A1(new_n458), .A2(G567), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT72), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n462), .B1(G2106), .B2(new_n456), .ZN(G319));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT73), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n467), .A2(new_n469), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OR3_X1    g054(.A1(new_n473), .A2(KEYINPUT74), .A3(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT74), .B1(new_n473), .B2(G2105), .ZN(new_n481));
  AND2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n473), .A2(new_n476), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  OAI21_X1  g063(.A(KEYINPUT75), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OR3_X1    g064(.A1(new_n487), .A2(KEYINPUT75), .A3(new_n488), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n483), .A2(new_n485), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND4_X1  g067(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n476), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT3), .B(G2104), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .A3(G138), .A4(new_n476), .ZN(new_n497));
  OR2_X1    g072(.A1(KEYINPUT76), .A2(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT76), .A2(G114), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n498), .A2(G2105), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n496), .A2(G126), .A3(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n495), .A2(new_n497), .A3(new_n503), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n508), .B(new_n510), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(G543), .B1(new_n511), .B2(new_n512), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n508), .A2(new_n510), .A3(G62), .ZN(new_n519));
  NAND2_X1  g094(.A1(G75), .A2(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n517), .A2(new_n521), .ZN(G166));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT77), .B(G89), .Z(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n513), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT78), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n524), .B(new_n528), .C1(new_n513), .C2(new_n525), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT5), .B(G543), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n531), .A2(G63), .A3(G651), .ZN(new_n532));
  INV_X1    g107(.A(new_n515), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G51), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n530), .A2(new_n532), .A3(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n531), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n518), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT80), .B(G90), .Z(new_n539));
  XOR2_X1   g114(.A(KEYINPUT79), .B(G52), .Z(new_n540));
  OAI22_X1  g115(.A1(new_n513), .A2(new_n539), .B1(new_n540), .B2(new_n515), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n531), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n518), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n513), .A2(new_n545), .B1(new_n515), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND3_X1  g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT8), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n552), .A2(KEYINPUT8), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT81), .Z(G188));
  NAND3_X1  g131(.A1(new_n508), .A2(new_n510), .A3(G65), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n557), .A2(KEYINPUT82), .A3(new_n558), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(G651), .A3(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n513), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G91), .ZN(new_n565));
  OAI211_X1 g140(.A(G53), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n563), .A2(new_n565), .A3(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  OR2_X1    g144(.A1(new_n511), .A2(new_n512), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n570), .A2(G88), .A3(new_n531), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n570), .A2(G50), .A3(G543), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n531), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n518), .ZN(G303));
  OAI211_X1 g149(.A(G49), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT83), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n508), .A2(new_n510), .ZN(new_n578));
  INV_X1    g153(.A(G74), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n564), .A2(G87), .B1(new_n580), .B2(G651), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(G288));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(new_n533), .B2(G48), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT84), .ZN(new_n587));
  INV_X1    g162(.A(G86), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n513), .B2(new_n588), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n570), .A2(KEYINPUT84), .A3(G86), .A4(new_n531), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n586), .A2(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n531), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n518), .ZN(new_n594));
  INV_X1    g169(.A(G85), .ZN(new_n595));
  INV_X1    g170(.A(G47), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n513), .A2(new_n595), .B1(new_n515), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n533), .A2(KEYINPUT86), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT86), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n515), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n601), .A2(G54), .A3(new_n603), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n531), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n605));
  OR2_X1    g180(.A1(new_n605), .A2(new_n518), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n513), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g184(.A(KEYINPUT85), .B(KEYINPUT10), .Z(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n600), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n600), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(G868), .B2(new_n616), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(G868), .B2(new_n616), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  INV_X1    g195(.A(new_n612), .ZN(new_n621));
  OAI21_X1  g196(.A(G868), .B1(new_n621), .B2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n486), .A2(G123), .ZN(new_n625));
  NOR2_X1   g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(new_n476), .B2(G111), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n480), .A2(new_n481), .ZN(new_n628));
  INV_X1    g203(.A(G135), .ZN(new_n629));
  OAI221_X1 g204(.A(new_n625), .B1(new_n626), .B2(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2096), .Z(new_n631));
  NAND3_X1  g206(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT88), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2427), .B(G2430), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT89), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2443), .B(G2446), .Z(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(G14), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(G401));
  XNOR2_X1  g228(.A(G2084), .B(G2090), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2072), .B(G2078), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT90), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT91), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n656), .B(KEYINPUT17), .Z(new_n660));
  INV_X1    g235(.A(new_n657), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n654), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n656), .A2(new_n657), .A3(new_n663), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT18), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G2096), .ZN(new_n668));
  INV_X1    g243(.A(G2100), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT92), .Z(new_n676));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n673), .A2(new_n674), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(new_n678), .B2(new_n675), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT93), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n682), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1981), .B(G1986), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT94), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n690), .B(new_n692), .ZN(G229));
  INV_X1    g268(.A(KEYINPUT101), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G5), .B2(G16), .ZN(new_n695));
  OR3_X1    g270(.A1(new_n694), .A2(G5), .A3(G16), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n695), .B(new_n696), .C1(G301), .C2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G1961), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g275(.A1(KEYINPUT95), .A2(G29), .ZN(new_n701));
  NOR2_X1   g276(.A1(KEYINPUT95), .A2(G29), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT24), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(G34), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(G34), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n708), .B1(new_n478), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G2084), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(G29), .A2(G32), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n482), .A2(G141), .ZN(new_n714));
  NAND3_X1  g289(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT26), .Z(new_n716));
  NAND3_X1  g291(.A1(new_n476), .A2(G105), .A3(G2104), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n486), .A2(G129), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n714), .A2(new_n716), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n713), .B1(new_n719), .B2(new_n709), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT27), .B(G1996), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n700), .B(new_n712), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT102), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n697), .A2(KEYINPUT23), .A3(G20), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT23), .ZN(new_n725));
  INV_X1    g300(.A(G20), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G16), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n724), .B(new_n727), .C1(new_n616), .C2(new_n697), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1956), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT30), .B(G28), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n720), .A2(new_n721), .B1(new_n709), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n704), .A2(G27), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G164), .B2(new_n704), .ZN(new_n734));
  INV_X1    g309(.A(G2078), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT31), .B(G11), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n732), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n697), .A2(G21), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G168), .B2(new_n697), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1966), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n630), .A2(new_n704), .ZN(new_n742));
  NOR2_X1   g317(.A1(G16), .A2(G19), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n548), .B2(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G1341), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n698), .B2(new_n699), .ZN(new_n746));
  NOR4_X1   g321(.A1(new_n738), .A2(new_n741), .A3(new_n742), .A4(new_n746), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n710), .A2(new_n711), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT99), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G4), .B2(G16), .ZN(new_n750));
  OR3_X1    g325(.A1(new_n749), .A2(G4), .A3(G16), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n750), .B(new_n751), .C1(new_n621), .C2(new_n697), .ZN(new_n752));
  INV_X1    g327(.A(G1348), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(KEYINPUT28), .B1(new_n704), .B2(G26), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n704), .A2(KEYINPUT28), .A3(G26), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n486), .A2(G128), .ZN(new_n758));
  NOR2_X1   g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(new_n476), .B2(G116), .ZN(new_n760));
  INV_X1    g335(.A(G140), .ZN(new_n761));
  OAI221_X1 g336(.A(new_n758), .B1(new_n759), .B2(new_n760), .C1(new_n628), .C2(new_n761), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n755), .B(new_n757), .C1(new_n762), .C2(G29), .ZN(new_n763));
  INV_X1    g338(.A(G2067), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n754), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n730), .A2(new_n747), .A3(new_n748), .A4(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(G16), .A2(G22), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G166), .B2(G16), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT97), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n772), .A2(G1971), .A3(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G1971), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n769), .A2(new_n770), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n771), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  OR2_X1    g353(.A1(G16), .A2(G23), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(G288), .B2(new_n697), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT33), .B(G1976), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n697), .A2(G6), .ZN(new_n783));
  INV_X1    g358(.A(G305), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(new_n697), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT32), .B(G1981), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n778), .A2(KEYINPUT34), .A3(new_n782), .A4(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT34), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n782), .A2(new_n774), .A3(new_n777), .ZN(new_n790));
  INV_X1    g365(.A(new_n786), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n785), .B(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n789), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n482), .A2(G131), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n486), .A2(G119), .ZN(new_n796));
  OR2_X1    g371(.A1(G95), .A2(G2105), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n797), .B(G2104), .C1(G107), .C2(new_n476), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n795), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(new_n703), .ZN(new_n800));
  INV_X1    g375(.A(G25), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n703), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT35), .B(G1991), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n803), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n800), .B(new_n805), .C1(new_n801), .C2(new_n703), .ZN(new_n806));
  INV_X1    g381(.A(G24), .ZN(new_n807));
  OAI21_X1  g382(.A(KEYINPUT96), .B1(new_n807), .B2(G16), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n807), .A2(KEYINPUT96), .A3(G16), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n808), .B(new_n809), .C1(new_n598), .C2(new_n697), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(G1986), .Z(new_n811));
  NAND3_X1  g386(.A1(new_n804), .A2(new_n806), .A3(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n794), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT98), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT98), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n794), .A2(new_n816), .A3(new_n813), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n815), .A2(KEYINPUT36), .A3(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT36), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n816), .B1(new_n794), .B2(new_n813), .ZN(new_n820));
  AOI211_X1 g395(.A(KEYINPUT98), .B(new_n812), .C1(new_n788), .C2(new_n793), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n767), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(G29), .A2(G33), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT25), .Z(new_n826));
  AOI22_X1  g401(.A1(new_n496), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n827));
  INV_X1    g402(.A(G139), .ZN(new_n828));
  OAI221_X1 g403(.A(new_n826), .B1(new_n476), .B2(new_n827), .C1(new_n628), .C2(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT100), .Z(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n824), .B1(new_n831), .B2(G29), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(G2072), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n704), .A2(G35), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(G162), .B2(new_n704), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT29), .B(G2090), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n744), .A2(G1341), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n823), .A2(new_n833), .A3(new_n837), .A4(new_n839), .ZN(G150));
  INV_X1    g415(.A(KEYINPUT103), .ZN(new_n841));
  NAND2_X1  g416(.A1(G150), .A2(new_n841), .ZN(new_n842));
  AOI211_X1 g417(.A(new_n838), .B(new_n767), .C1(new_n818), .C2(new_n822), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n843), .A2(KEYINPUT103), .A3(new_n833), .A4(new_n837), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(G311));
  AOI22_X1  g420(.A1(new_n531), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n518), .ZN(new_n847));
  INV_X1    g422(.A(G93), .ZN(new_n848));
  INV_X1    g423(.A(G55), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n513), .A2(new_n848), .B1(new_n515), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n548), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n851), .B1(new_n544), .B2(new_n547), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g432(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n621), .A2(new_n619), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n854), .B1(new_n861), .B2(G860), .ZN(G145));
  XNOR2_X1  g437(.A(new_n630), .B(KEYINPUT104), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(G160), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(G160), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n491), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n866), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n868), .A2(G162), .A3(new_n864), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n867), .A2(new_n799), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n799), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI22_X1  g447(.A1(new_n482), .A2(G142), .B1(G130), .B2(new_n486), .ZN(new_n873));
  NOR2_X1   g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(new_n476), .B2(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n633), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n762), .B(G164), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n878), .A2(new_n719), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n719), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n830), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n879), .A2(new_n880), .A3(new_n829), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  INV_X1    g460(.A(new_n877), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n885), .A2(new_n881), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n872), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(G37), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n884), .B(new_n887), .C1(new_n870), .C2(new_n871), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g468(.A1(new_n852), .A2(G868), .ZN(new_n894));
  XNOR2_X1  g469(.A(G305), .B(G288), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n598), .B(G303), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT42), .Z(new_n898));
  NAND4_X1  g473(.A1(new_n563), .A2(KEYINPUT105), .A3(new_n565), .A4(new_n567), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n612), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT105), .ZN(new_n901));
  NAND2_X1  g476(.A1(G299), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n612), .A2(new_n902), .A3(new_n899), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT41), .ZN(new_n907));
  INV_X1    g482(.A(new_n905), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n902), .B1(new_n612), .B2(new_n899), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n904), .A2(KEYINPUT41), .A3(new_n905), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n612), .A2(new_n619), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n857), .ZN(new_n914));
  MUX2_X1   g489(.A(new_n906), .B(new_n912), .S(new_n914), .Z(new_n915));
  AOI21_X1  g490(.A(new_n898), .B1(new_n915), .B2(KEYINPUT106), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(KEYINPUT106), .ZN(new_n917));
  MUX2_X1   g492(.A(new_n916), .B(new_n898), .S(new_n917), .Z(new_n918));
  AOI21_X1  g493(.A(new_n894), .B1(new_n918), .B2(G868), .ZN(G295));
  AOI21_X1  g494(.A(new_n894), .B1(new_n918), .B2(G868), .ZN(G331));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n922));
  NOR2_X1   g497(.A1(G286), .A2(G171), .ZN(new_n923));
  AOI22_X1  g498(.A1(new_n527), .A2(new_n529), .B1(G51), .B2(new_n533), .ZN(new_n924));
  AOI21_X1  g499(.A(G301), .B1(new_n924), .B2(new_n532), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n857), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(G286), .A2(G171), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n532), .A3(G301), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n927), .A2(new_n928), .A3(new_n855), .A4(new_n856), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n926), .A2(KEYINPUT107), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n931), .B(new_n857), .C1(new_n923), .C2(new_n925), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n930), .A2(new_n910), .A3(new_n911), .A4(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n926), .A2(new_n929), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n934), .B1(new_n935), .B2(new_n906), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n908), .A2(new_n909), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n937), .A2(KEYINPUT108), .A3(new_n926), .A4(new_n929), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n933), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n939), .A2(new_n897), .ZN(new_n940));
  INV_X1    g515(.A(new_n897), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n933), .A2(new_n936), .A3(new_n941), .A4(new_n938), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n890), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n922), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n942), .A2(new_n890), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n935), .A2(new_n910), .A3(new_n911), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n906), .B1(new_n930), .B2(new_n932), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n897), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n945), .A2(KEYINPUT43), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n921), .B1(new_n944), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n940), .B2(new_n943), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n922), .A3(new_n948), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT44), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n950), .A2(new_n953), .A3(KEYINPUT109), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n944), .A2(new_n949), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n939), .A2(new_n897), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n922), .B1(new_n945), .B2(new_n958), .ZN(new_n959));
  AND4_X1   g534(.A1(new_n922), .A2(new_n948), .A3(new_n890), .A4(new_n942), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n921), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n955), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n954), .A2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n495), .A2(new_n497), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n503), .A2(new_n504), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n471), .A2(new_n477), .A3(G40), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1996), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n719), .B(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n762), .B(new_n764), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n799), .A2(new_n803), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n799), .A2(new_n803), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G1986), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n979), .B1(new_n980), .B2(new_n598), .ZN(new_n981));
  NOR2_X1   g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n972), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n971), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n968), .B1(new_n505), .B2(new_n964), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n986), .A2(G1996), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n967), .A2(new_n971), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT58), .B(G1341), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n548), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT59), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT59), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n994), .B(new_n548), .C1(new_n988), .C2(new_n991), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT56), .B(G2072), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT118), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n970), .A2(new_n984), .A3(new_n985), .A4(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n967), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n505), .A2(KEYINPUT50), .A3(new_n964), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n971), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n999), .B1(new_n1003), .B2(G1956), .ZN(new_n1004));
  XNOR2_X1  g579(.A(G299), .B(KEYINPUT57), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT61), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n505), .A2(KEYINPUT50), .A3(new_n964), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT50), .B1(new_n505), .B2(new_n964), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n984), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1956), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT57), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G299), .B(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1014), .A3(new_n999), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1006), .A2(new_n1007), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1007), .B1(new_n1006), .B2(new_n1015), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n996), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n1010), .A2(new_n753), .B1(new_n764), .B2(new_n989), .ZN(new_n1021));
  AND3_X1   g596(.A1(new_n1021), .A2(KEYINPUT60), .A3(new_n621), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n621), .B1(new_n1021), .B2(KEYINPUT60), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n1022), .A2(new_n1023), .B1(KEYINPUT60), .B2(new_n1021), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n996), .B(KEYINPUT119), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1020), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1021), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1015), .A2(new_n1027), .A3(new_n612), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1026), .A2(new_n1006), .A3(new_n1028), .ZN(new_n1029));
  XOR2_X1   g604(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1030));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n970), .A2(new_n735), .A3(new_n984), .A4(new_n985), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n1031), .A2(new_n1032), .B1(new_n1010), .B2(new_n699), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1034));
  OR2_X1    g609(.A1(new_n1034), .A2(G171), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n967), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(KEYINPUT115), .A3(new_n984), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT45), .B1(new_n505), .B2(new_n964), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1039), .B1(new_n1040), .B2(new_n971), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n505), .A2(new_n964), .A3(new_n968), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1031), .A2(G2078), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1038), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1033), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(G171), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1030), .B1(new_n1035), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n775), .B1(new_n986), .B2(new_n987), .ZN(new_n1048));
  INV_X1    g623(.A(G2090), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1049), .B(new_n984), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT55), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(G303), .B2(G8), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1052), .B(G8), .C1(new_n517), .C2(new_n521), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1053), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G8), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1057), .A2(KEYINPUT114), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1051), .A2(G8), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n1057), .B(new_n1060), .C1(new_n1048), .C2(new_n1050), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT111), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n967), .B2(new_n971), .ZN(new_n1064));
  INV_X1    g639(.A(G1976), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G288), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1063), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(G288), .A2(new_n1065), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n585), .A2(G651), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n533), .A2(G48), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n513), .A2(new_n588), .ZN(new_n1076));
  OAI21_X1  g651(.A(G1981), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  XOR2_X1   g652(.A(KEYINPUT112), .B(G1981), .Z(new_n1078));
  NAND3_X1  g653(.A1(new_n586), .A2(new_n591), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT113), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT49), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1064), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT49), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1080), .A2(new_n1081), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1067), .A2(new_n1063), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1072), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT123), .B1(new_n1062), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1089), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1051), .A2(G8), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1060), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1051), .A2(KEYINPUT114), .A3(G8), .A4(new_n1056), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1091), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1047), .B1(new_n1090), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1034), .B2(G171), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1101), .B1(new_n1045), .B2(G171), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1033), .A2(KEYINPUT124), .A3(G301), .A4(new_n1044), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT125), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT125), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1100), .A2(new_n1106), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n711), .B(new_n984), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1110), .A2(new_n1111), .A3(new_n711), .A4(new_n984), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1038), .A2(new_n1042), .A3(new_n1041), .ZN(new_n1114));
  INV_X1    g689(.A(G1966), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1113), .A2(new_n1116), .ZN(new_n1117));
  AND4_X1   g692(.A1(KEYINPUT120), .A2(new_n1117), .A3(G8), .A4(G286), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1057), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT120), .B1(new_n1119), .B2(G286), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1113), .A2(new_n1116), .A3(G168), .ZN(new_n1122));
  AND2_X1   g697(.A1(KEYINPUT121), .A2(G8), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1122), .A2(KEYINPUT51), .A3(new_n1123), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1105), .A2(new_n1107), .B1(new_n1121), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1029), .A2(new_n1098), .A3(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1089), .A2(new_n1092), .A3(new_n1056), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1087), .A2(new_n1065), .ZN(new_n1132));
  INV_X1    g707(.A(G288), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1064), .B1(new_n1134), .B2(new_n1079), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1119), .A2(G168), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(new_n1091), .A3(new_n1095), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1056), .A2(KEYINPUT117), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1051), .A2(G8), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1140), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1138), .B1(new_n1092), .B2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1136), .A2(new_n1091), .A3(new_n1141), .A4(new_n1143), .ZN(new_n1144));
  AOI211_X1 g719(.A(new_n1131), .B(new_n1135), .C1(new_n1139), .C2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1130), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1121), .A2(new_n1128), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1046), .B1(new_n1097), .B2(new_n1090), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1149), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1147), .B1(new_n1121), .B2(new_n1128), .ZN(new_n1153));
  NOR3_X1   g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n983), .B1(new_n1146), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n972), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n974), .A2(new_n977), .A3(new_n975), .ZN(new_n1157));
  OR2_X1    g732(.A1(new_n762), .A2(G2067), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n975), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n972), .B1(new_n1160), .B2(new_n719), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT46), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1156), .B2(G1996), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n972), .A2(KEYINPUT46), .A3(new_n973), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  XOR2_X1   g740(.A(new_n1165), .B(KEYINPUT47), .Z(new_n1166));
  OR2_X1    g741(.A1(new_n979), .A2(new_n1156), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n972), .A2(new_n982), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT48), .ZN(new_n1169));
  AOI211_X1 g744(.A(new_n1159), .B(new_n1166), .C1(new_n1167), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1155), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g746(.A(G229), .B1(new_n951), .B2(new_n952), .ZN(new_n1173));
  NAND3_X1  g747(.A1(new_n670), .A2(G319), .A3(new_n671), .ZN(new_n1174));
  NOR2_X1   g748(.A1(G401), .A2(new_n1174), .ZN(new_n1175));
  AND2_X1   g749(.A1(new_n892), .A2(new_n1175), .ZN(new_n1176));
  AND2_X1   g750(.A1(new_n1173), .A2(new_n1176), .ZN(G308));
  NAND2_X1  g751(.A1(new_n1173), .A2(new_n1176), .ZN(G225));
endmodule


