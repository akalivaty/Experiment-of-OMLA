

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592;

  XOR2_X1 U323 ( .A(G22GAT), .B(G155GAT), .Z(n385) );
  AND2_X1 U324 ( .A1(G231GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U325 ( .A(n385), .B(n291), .ZN(n386) );
  XNOR2_X1 U326 ( .A(n387), .B(n386), .ZN(n388) );
  INV_X1 U327 ( .A(G64GAT), .ZN(n393) );
  XNOR2_X1 U328 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U329 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U330 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U331 ( .A(n396), .B(n395), .ZN(n400) );
  XNOR2_X1 U332 ( .A(n353), .B(KEYINPUT26), .ZN(n578) );
  INV_X1 U333 ( .A(n578), .ZN(n551) );
  XOR2_X1 U334 ( .A(n330), .B(n364), .Z(n479) );
  NOR2_X1 U335 ( .A1(n539), .A2(n481), .ZN(n571) );
  XNOR2_X1 U336 ( .A(n482), .B(G190GAT), .ZN(n483) );
  XNOR2_X1 U337 ( .A(n460), .B(KEYINPUT108), .ZN(n461) );
  XNOR2_X1 U338 ( .A(n484), .B(n483), .ZN(G1351GAT) );
  XNOR2_X1 U339 ( .A(n462), .B(n461), .ZN(G1329GAT) );
  NAND2_X1 U340 ( .A1(G226GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U341 ( .A(G36GAT), .B(G190GAT), .Z(n404) );
  XNOR2_X1 U342 ( .A(n292), .B(n404), .ZN(n306) );
  XOR2_X1 U343 ( .A(KEYINPUT80), .B(G211GAT), .Z(n294) );
  XNOR2_X1 U344 ( .A(G8GAT), .B(G183GAT), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n387) );
  XOR2_X1 U346 ( .A(G64GAT), .B(G92GAT), .Z(n296) );
  XNOR2_X1 U347 ( .A(G176GAT), .B(G204GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n454) );
  XNOR2_X1 U349 ( .A(n387), .B(n454), .ZN(n301) );
  XOR2_X1 U350 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n298) );
  XNOR2_X1 U351 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n344) );
  XNOR2_X1 U353 ( .A(n344), .B(KEYINPUT97), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n299), .B(KEYINPUT96), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U356 ( .A(n302), .B(KEYINPUT98), .Z(n304) );
  XOR2_X1 U357 ( .A(G197GAT), .B(KEYINPUT21), .Z(n309) );
  XNOR2_X1 U358 ( .A(G218GAT), .B(n309), .ZN(n303) );
  XNOR2_X1 U359 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U360 ( .A(n306), .B(n305), .Z(n526) );
  INV_X1 U361 ( .A(n526), .ZN(n513) );
  XOR2_X1 U362 ( .A(G78GAT), .B(G148GAT), .Z(n308) );
  XNOR2_X1 U363 ( .A(G106GAT), .B(KEYINPUT72), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n455) );
  XNOR2_X1 U365 ( .A(n385), .B(n309), .ZN(n311) );
  XOR2_X1 U366 ( .A(KEYINPUT22), .B(KEYINPUT90), .Z(n310) );
  XNOR2_X1 U367 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U368 ( .A(KEYINPUT89), .B(KEYINPUT91), .Z(n313) );
  XNOR2_X1 U369 ( .A(G211GAT), .B(G204GAT), .ZN(n312) );
  XOR2_X1 U370 ( .A(n313), .B(n312), .Z(n314) );
  XNOR2_X1 U371 ( .A(n315), .B(n314), .ZN(n319) );
  INV_X1 U372 ( .A(n319), .ZN(n317) );
  NAND2_X1 U373 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  INV_X1 U374 ( .A(n318), .ZN(n316) );
  NAND2_X1 U375 ( .A1(n317), .A2(n316), .ZN(n321) );
  NAND2_X1 U376 ( .A1(n319), .A2(n318), .ZN(n320) );
  NAND2_X1 U377 ( .A1(n321), .A2(n320), .ZN(n327) );
  XOR2_X1 U378 ( .A(G162GAT), .B(KEYINPUT77), .Z(n323) );
  XNOR2_X1 U379 ( .A(G50GAT), .B(G218GAT), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n323), .B(n322), .ZN(n414) );
  XNOR2_X1 U381 ( .A(n414), .B(KEYINPUT24), .ZN(n325) );
  INV_X1 U382 ( .A(KEYINPUT23), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n455), .B(n328), .ZN(n330) );
  XOR2_X1 U384 ( .A(G141GAT), .B(KEYINPUT3), .Z(n329) );
  XOR2_X1 U385 ( .A(KEYINPUT2), .B(n329), .Z(n364) );
  XOR2_X1 U386 ( .A(G15GAT), .B(G127GAT), .Z(n392) );
  XOR2_X1 U387 ( .A(KEYINPUT88), .B(G99GAT), .Z(n332) );
  XNOR2_X1 U388 ( .A(G43GAT), .B(G190GAT), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U390 ( .A(n392), .B(n333), .Z(n335) );
  NAND2_X1 U391 ( .A1(G227GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n348) );
  XOR2_X1 U393 ( .A(G176GAT), .B(G71GAT), .Z(n337) );
  XNOR2_X1 U394 ( .A(G113GAT), .B(KEYINPUT20), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U396 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n339) );
  XNOR2_X1 U397 ( .A(KEYINPUT87), .B(G183GAT), .ZN(n338) );
  XNOR2_X1 U398 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U399 ( .A(n341), .B(n340), .Z(n346) );
  XOR2_X1 U400 ( .A(G120GAT), .B(KEYINPUT84), .Z(n343) );
  XNOR2_X1 U401 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n368) );
  XNOR2_X1 U403 ( .A(n368), .B(n344), .ZN(n345) );
  XNOR2_X1 U404 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U405 ( .A(n348), .B(n347), .Z(n528) );
  INV_X1 U406 ( .A(n528), .ZN(n539) );
  NOR2_X1 U407 ( .A1(n539), .A2(n513), .ZN(n349) );
  NOR2_X1 U408 ( .A1(n479), .A2(n349), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n350), .B(KEYINPUT101), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n351), .B(KEYINPUT25), .ZN(n355) );
  NAND2_X1 U411 ( .A1(n479), .A2(n539), .ZN(n352) );
  XNOR2_X1 U412 ( .A(n352), .B(KEYINPUT100), .ZN(n353) );
  XOR2_X1 U413 ( .A(KEYINPUT27), .B(n526), .Z(n378) );
  NOR2_X1 U414 ( .A1(n578), .A2(n378), .ZN(n354) );
  NOR2_X1 U415 ( .A1(n355), .A2(n354), .ZN(n377) );
  XOR2_X1 U416 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n357) );
  XNOR2_X1 U417 ( .A(KEYINPUT92), .B(KEYINPUT1), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n376) );
  XOR2_X1 U419 ( .A(G85GAT), .B(G155GAT), .Z(n359) );
  XNOR2_X1 U420 ( .A(G127GAT), .B(G148GAT), .ZN(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U422 ( .A(KEYINPUT4), .B(KEYINPUT95), .Z(n361) );
  XNOR2_X1 U423 ( .A(G57GAT), .B(KEYINPUT94), .ZN(n360) );
  XNOR2_X1 U424 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U425 ( .A(n363), .B(n362), .Z(n374) );
  INV_X1 U426 ( .A(n364), .ZN(n365) );
  XNOR2_X1 U427 ( .A(n365), .B(KEYINPUT93), .ZN(n367) );
  NAND2_X1 U428 ( .A1(G225GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n372) );
  XOR2_X1 U430 ( .A(G162GAT), .B(n368), .Z(n370) );
  XOR2_X1 U431 ( .A(G113GAT), .B(G1GAT), .Z(n434) );
  XNOR2_X1 U432 ( .A(G29GAT), .B(n434), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U436 ( .A(n376), .B(n375), .ZN(n524) );
  NOR2_X1 U437 ( .A1(n377), .A2(n524), .ZN(n382) );
  XOR2_X1 U438 ( .A(KEYINPUT28), .B(n479), .Z(n537) );
  INV_X1 U439 ( .A(n537), .ZN(n531) );
  INV_X1 U440 ( .A(n524), .ZN(n509) );
  NOR2_X1 U441 ( .A1(n509), .A2(n378), .ZN(n379) );
  XNOR2_X1 U442 ( .A(KEYINPUT99), .B(n379), .ZN(n535) );
  OR2_X1 U443 ( .A1(n528), .A2(n535), .ZN(n380) );
  NOR2_X1 U444 ( .A1(n531), .A2(n380), .ZN(n381) );
  NOR2_X1 U445 ( .A1(n382), .A2(n381), .ZN(n384) );
  INV_X1 U446 ( .A(KEYINPUT102), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n487) );
  XOR2_X1 U448 ( .A(n388), .B(KEYINPUT14), .Z(n391) );
  XNOR2_X1 U449 ( .A(G71GAT), .B(G57GAT), .ZN(n389) );
  XNOR2_X1 U450 ( .A(n389), .B(KEYINPUT13), .ZN(n451) );
  XNOR2_X1 U451 ( .A(n451), .B(KEYINPUT15), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n396) );
  XNOR2_X1 U453 ( .A(n392), .B(G78GAT), .ZN(n394) );
  XOR2_X1 U454 ( .A(KEYINPUT12), .B(KEYINPUT81), .Z(n398) );
  XNOR2_X1 U455 ( .A(G1GAT), .B(KEYINPUT82), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n468) );
  INV_X1 U458 ( .A(n468), .ZN(n586) );
  XOR2_X1 U459 ( .A(G92GAT), .B(KEYINPUT10), .Z(n402) );
  XNOR2_X1 U460 ( .A(G134GAT), .B(G106GAT), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U462 ( .A(n404), .B(n403), .Z(n406) );
  NAND2_X1 U463 ( .A1(G232GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n419) );
  XOR2_X1 U465 ( .A(KEYINPUT11), .B(KEYINPUT78), .Z(n408) );
  XNOR2_X1 U466 ( .A(KEYINPUT9), .B(KEYINPUT79), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X1 U468 ( .A(G99GAT), .B(G85GAT), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n409), .B(KEYINPUT73), .ZN(n443) );
  XOR2_X1 U470 ( .A(n410), .B(n443), .Z(n417) );
  XOR2_X1 U471 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n412) );
  XNOR2_X1 U472 ( .A(G43GAT), .B(G29GAT), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U474 ( .A(KEYINPUT7), .B(n413), .Z(n440) );
  INV_X1 U475 ( .A(n440), .ZN(n415) );
  XOR2_X1 U476 ( .A(n415), .B(n414), .Z(n416) );
  XNOR2_X1 U477 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U478 ( .A(n419), .B(n418), .ZN(n546) );
  XOR2_X1 U479 ( .A(n546), .B(KEYINPUT36), .Z(n590) );
  NOR2_X1 U480 ( .A1(n586), .A2(n590), .ZN(n420) );
  NAND2_X1 U481 ( .A1(n487), .A2(n420), .ZN(n422) );
  XOR2_X1 U482 ( .A(KEYINPUT105), .B(KEYINPUT37), .Z(n421) );
  XNOR2_X1 U483 ( .A(n422), .B(n421), .ZN(n521) );
  XOR2_X1 U484 ( .A(KEYINPUT66), .B(KEYINPUT65), .Z(n424) );
  XNOR2_X1 U485 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n423) );
  XNOR2_X1 U486 ( .A(n424), .B(n423), .ZN(n438) );
  XOR2_X1 U487 ( .A(G197GAT), .B(G22GAT), .Z(n426) );
  XNOR2_X1 U488 ( .A(G36GAT), .B(G50GAT), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U490 ( .A(KEYINPUT30), .B(G15GAT), .Z(n428) );
  XNOR2_X1 U491 ( .A(G169GAT), .B(G141GAT), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U493 ( .A(n430), .B(n429), .Z(n436) );
  XOR2_X1 U494 ( .A(KEYINPUT29), .B(G8GAT), .Z(n432) );
  NAND2_X1 U495 ( .A1(G229GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U496 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U497 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U499 ( .A(n438), .B(n437), .Z(n439) );
  XOR2_X1 U500 ( .A(n440), .B(n439), .Z(n580) );
  INV_X1 U501 ( .A(n580), .ZN(n552) );
  XOR2_X1 U502 ( .A(KEYINPUT71), .B(KEYINPUT74), .Z(n442) );
  XNOR2_X1 U503 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n441) );
  XNOR2_X1 U504 ( .A(n442), .B(n441), .ZN(n447) );
  XOR2_X1 U505 ( .A(n443), .B(KEYINPUT76), .Z(n445) );
  NAND2_X1 U506 ( .A1(G230GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U507 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U508 ( .A(n447), .B(n446), .Z(n453) );
  XOR2_X1 U509 ( .A(KEYINPUT75), .B(KEYINPUT31), .Z(n449) );
  XNOR2_X1 U510 ( .A(KEYINPUT70), .B(KEYINPUT32), .ZN(n448) );
  XNOR2_X1 U511 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U512 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n453), .B(n452), .ZN(n457) );
  XOR2_X1 U514 ( .A(n455), .B(n454), .Z(n456) );
  XNOR2_X1 U515 ( .A(n457), .B(n456), .ZN(n583) );
  NOR2_X1 U516 ( .A1(n552), .A2(n583), .ZN(n489) );
  NAND2_X1 U517 ( .A1(n521), .A2(n489), .ZN(n458) );
  XNOR2_X1 U518 ( .A(n458), .B(KEYINPUT38), .ZN(n459) );
  XNOR2_X1 U519 ( .A(KEYINPUT106), .B(n459), .ZN(n506) );
  NOR2_X1 U520 ( .A1(n513), .A2(n506), .ZN(n462) );
  INV_X1 U521 ( .A(G36GAT), .ZN(n460) );
  XNOR2_X1 U522 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n476) );
  XOR2_X1 U523 ( .A(KEYINPUT117), .B(KEYINPUT47), .Z(n467) );
  XOR2_X1 U524 ( .A(KEYINPUT116), .B(n468), .Z(n572) );
  XOR2_X1 U525 ( .A(KEYINPUT41), .B(n583), .Z(n566) );
  INV_X1 U526 ( .A(n566), .ZN(n555) );
  NOR2_X1 U527 ( .A1(n555), .A2(n552), .ZN(n463) );
  XNOR2_X1 U528 ( .A(n463), .B(KEYINPUT46), .ZN(n464) );
  NOR2_X1 U529 ( .A1(n572), .A2(n464), .ZN(n465) );
  INV_X1 U530 ( .A(n546), .ZN(n561) );
  NAND2_X1 U531 ( .A1(n465), .A2(n561), .ZN(n466) );
  XNOR2_X1 U532 ( .A(n467), .B(n466), .ZN(n474) );
  NOR2_X1 U533 ( .A1(n468), .A2(n590), .ZN(n469) );
  XOR2_X1 U534 ( .A(KEYINPUT45), .B(n469), .Z(n470) );
  NOR2_X1 U535 ( .A1(n583), .A2(n470), .ZN(n471) );
  XOR2_X1 U536 ( .A(KEYINPUT118), .B(n471), .Z(n472) );
  NOR2_X1 U537 ( .A1(n580), .A2(n472), .ZN(n473) );
  NOR2_X1 U538 ( .A1(n474), .A2(n473), .ZN(n475) );
  XNOR2_X1 U539 ( .A(n476), .B(n475), .ZN(n536) );
  NOR2_X1 U540 ( .A1(n536), .A2(n513), .ZN(n477) );
  XNOR2_X1 U541 ( .A(n477), .B(KEYINPUT54), .ZN(n478) );
  NAND2_X1 U542 ( .A1(n478), .A2(n509), .ZN(n579) );
  NOR2_X1 U543 ( .A1(n479), .A2(n579), .ZN(n480) );
  XNOR2_X1 U544 ( .A(n480), .B(KEYINPUT55), .ZN(n481) );
  NAND2_X1 U545 ( .A1(n571), .A2(n546), .ZN(n484) );
  XOR2_X1 U546 ( .A(KEYINPUT58), .B(KEYINPUT125), .Z(n482) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n492) );
  NAND2_X1 U548 ( .A1(n586), .A2(n561), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n485), .B(KEYINPUT83), .ZN(n486) );
  XNOR2_X1 U550 ( .A(KEYINPUT16), .B(n486), .ZN(n488) );
  AND2_X1 U551 ( .A1(n488), .A2(n487), .ZN(n508) );
  NAND2_X1 U552 ( .A1(n489), .A2(n508), .ZN(n490) );
  XNOR2_X1 U553 ( .A(KEYINPUT103), .B(n490), .ZN(n496) );
  NAND2_X1 U554 ( .A1(n496), .A2(n524), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(G1324GAT) );
  NAND2_X1 U556 ( .A1(n496), .A2(n526), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n493), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U558 ( .A(G15GAT), .B(KEYINPUT35), .Z(n495) );
  NAND2_X1 U559 ( .A1(n496), .A2(n528), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n495), .B(n494), .ZN(G1326GAT) );
  NAND2_X1 U561 ( .A1(n496), .A2(n531), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n497), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U563 ( .A1(n506), .A2(n509), .ZN(n501) );
  XOR2_X1 U564 ( .A(KEYINPUT104), .B(KEYINPUT107), .Z(n499) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U566 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n503) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(n505) );
  NOR2_X1 U571 ( .A1(n539), .A2(n506), .ZN(n504) );
  XOR2_X1 U572 ( .A(n505), .B(n504), .Z(G1330GAT) );
  NOR2_X1 U573 ( .A1(n537), .A2(n506), .ZN(n507) );
  XOR2_X1 U574 ( .A(G50GAT), .B(n507), .Z(G1331GAT) );
  NOR2_X1 U575 ( .A1(n580), .A2(n555), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n522), .A2(n508), .ZN(n517) );
  NOR2_X1 U577 ( .A1(n509), .A2(n517), .ZN(n511) );
  XNOR2_X1 U578 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n510) );
  XNOR2_X1 U579 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U580 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n513), .A2(n517), .ZN(n514) );
  XOR2_X1 U582 ( .A(KEYINPUT112), .B(n514), .Z(n515) );
  XNOR2_X1 U583 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NOR2_X1 U584 ( .A1(n539), .A2(n517), .ZN(n516) );
  XOR2_X1 U585 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U586 ( .A1(n537), .A2(n517), .ZN(n519) );
  XNOR2_X1 U587 ( .A(KEYINPUT43), .B(KEYINPUT113), .ZN(n518) );
  XNOR2_X1 U588 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U589 ( .A(G78GAT), .B(n520), .Z(G1335GAT) );
  NAND2_X1 U590 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U591 ( .A(KEYINPUT114), .B(n523), .Z(n532) );
  NAND2_X1 U592 ( .A1(n524), .A2(n532), .ZN(n525) );
  XNOR2_X1 U593 ( .A(G85GAT), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U594 ( .A1(n526), .A2(n532), .ZN(n527) );
  XNOR2_X1 U595 ( .A(G92GAT), .B(n527), .ZN(G1337GAT) );
  XOR2_X1 U596 ( .A(G99GAT), .B(KEYINPUT115), .Z(n530) );
  NAND2_X1 U597 ( .A1(n528), .A2(n532), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(G1338GAT) );
  NAND2_X1 U599 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n533), .B(KEYINPUT44), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(n534), .ZN(G1339GAT) );
  XOR2_X1 U602 ( .A(G113GAT), .B(KEYINPUT119), .Z(n541) );
  NOR2_X1 U603 ( .A1(n536), .A2(n535), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n550), .A2(n537), .ZN(n538) );
  NOR2_X1 U605 ( .A1(n539), .A2(n538), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n547), .A2(n580), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U609 ( .A1(n547), .A2(n566), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  NAND2_X1 U611 ( .A1(n572), .A2(n547), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n544), .B(KEYINPUT50), .ZN(n545) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n560) );
  NOR2_X1 U618 ( .A1(n552), .A2(n560), .ZN(n553) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n553), .Z(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT120), .B(n554), .ZN(G1344GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n560), .ZN(n557) );
  XNOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n468), .A2(n560), .ZN(n559) );
  XOR2_X1 U626 ( .A(G155GAT), .B(n559), .Z(G1346GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n563) );
  XNOR2_X1 U628 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G162GAT), .B(n564), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n571), .A2(n580), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT56), .Z(n568) );
  NAND2_X1 U634 ( .A1(n571), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(KEYINPUT124), .ZN(n574) );
  XNOR2_X1 U640 ( .A(G183GAT), .B(n574), .ZN(G1350GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n576) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT126), .B(n577), .Z(n582) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n588) );
  NAND2_X1 U646 ( .A1(n588), .A2(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U649 ( .A1(n588), .A2(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n588), .A2(n586), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U653 ( .A(n588), .ZN(n589) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

