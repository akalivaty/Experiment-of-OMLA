//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(new_n204), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n209), .B1(new_n212), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G87), .B(G97), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT64), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(KEYINPUT76), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT9), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n210), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G50), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n252), .B1(new_n203), .B2(G20), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n251), .A2(new_n253), .B1(new_n252), .B2(new_n248), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT66), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT8), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G58), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(KEYINPUT66), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n256), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G68), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n252), .A2(new_n221), .A3(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(G20), .A2(G33), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n265), .A2(G20), .B1(G150), .B2(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n250), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n246), .B(new_n254), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n269), .B1(new_n263), .B2(new_n267), .ZN(new_n271));
  INV_X1    g0071(.A(new_n254), .ZN(new_n272));
  OAI21_X1  g0072(.A(KEYINPUT9), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G222), .A2(G1698), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G223), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  OAI211_X1 g0083(.A(G1), .B(G13), .C1(new_n261), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n275), .A2(new_n277), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(new_n215), .ZN(new_n286));
  AND2_X1   g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n210), .ZN(new_n288));
  INV_X1    g0088(.A(G45), .ZN(new_n289));
  AOI21_X1  g0089(.A(G1), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n282), .A2(new_n286), .B1(G226), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT65), .ZN(new_n293));
  INV_X1    g0093(.A(new_n290), .ZN(new_n294));
  OAI21_X1  g0094(.A(G274), .B1(new_n287), .B2(new_n210), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n284), .A2(KEYINPUT65), .A3(new_n290), .A4(G274), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G200), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n292), .A2(G190), .A3(new_n298), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n274), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT69), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT10), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n300), .A2(new_n305), .A3(new_n301), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT68), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n274), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n270), .A2(new_n273), .A3(KEYINPUT68), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n304), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n274), .A2(new_n307), .ZN(new_n311));
  INV_X1    g0111(.A(new_n306), .ZN(new_n312));
  AND4_X1   g0112(.A1(new_n304), .A2(new_n311), .A3(new_n312), .A4(new_n309), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n303), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n271), .A2(new_n272), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n299), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n292), .A2(new_n318), .A3(new_n298), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n203), .A2(G20), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n251), .A2(G77), .A3(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(G77), .B2(new_n247), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(new_n262), .B1(G20), .B2(G77), .ZN(new_n327));
  INV_X1    g0127(.A(new_n266), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n255), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n324), .B1(new_n329), .B2(new_n250), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n278), .A2(G238), .A3(G1698), .ZN(new_n331));
  OR2_X1    g0131(.A1(KEYINPUT67), .A2(G107), .ZN(new_n332));
  NAND2_X1  g0132(.A1(KEYINPUT67), .A2(G107), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n331), .B1(new_n278), .B2(new_n335), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n285), .A2(new_n222), .A3(G1698), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n288), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n291), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n338), .B(new_n298), .C1(new_n216), .C2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n330), .B1(new_n340), .B2(new_n316), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(G179), .B2(new_n340), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(G200), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n330), .C1(new_n344), .C2(new_n340), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n314), .A2(new_n321), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n248), .A2(new_n264), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT12), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n262), .A2(G77), .B1(G20), .B2(new_n264), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n252), .B2(new_n328), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n351), .A2(KEYINPUT11), .A3(new_n250), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n251), .A2(G68), .A3(new_n322), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n349), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT11), .B1(new_n351), .B2(new_n250), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n298), .A2(KEYINPUT70), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT70), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n296), .A2(new_n359), .A3(new_n297), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G97), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n222), .A2(G1698), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(G226), .B2(G1698), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n361), .B1(new_n363), .B2(new_n285), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n288), .B1(new_n291), .B2(G238), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n358), .A2(new_n360), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT13), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT13), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n358), .A2(new_n365), .A3(new_n368), .A4(new_n360), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT14), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(G169), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n367), .A2(G179), .A3(new_n369), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n371), .B1(new_n370), .B2(G169), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n357), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n356), .B1(new_n370), .B2(new_n344), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n367), .B2(new_n369), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n347), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n259), .B1(new_n255), .B2(KEYINPUT66), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n322), .ZN(new_n385));
  OR2_X1    g0185(.A1(new_n385), .A2(KEYINPUT74), .ZN(new_n386));
  INV_X1    g0186(.A(new_n251), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n385), .B2(KEYINPUT74), .ZN(new_n388));
  INV_X1    g0188(.A(new_n384), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n386), .A2(new_n388), .B1(new_n248), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT71), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n276), .B2(G33), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n261), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT72), .B1(new_n261), .B2(KEYINPUT3), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT72), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(new_n276), .A3(G33), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(G20), .B1(new_n395), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI211_X1 g0202(.A(KEYINPUT7), .B(G20), .C1(new_n395), .C2(new_n399), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT73), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n396), .A2(new_n398), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n393), .A2(new_n394), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n204), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n264), .B1(new_n407), .B2(KEYINPUT7), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT73), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n400), .A2(new_n401), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n221), .A2(new_n264), .ZN(new_n413));
  NOR2_X1   g0213(.A1(G58), .A2(G68), .ZN(new_n414));
  OAI21_X1  g0214(.A(G20), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n266), .A2(G159), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT16), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n269), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n401), .B1(new_n278), .B2(G20), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n264), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n418), .B1(new_n423), .B2(new_n417), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n391), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  AND2_X1   g0225(.A1(G226), .A2(G1698), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n395), .A2(new_n399), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT75), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n395), .A2(KEYINPUT75), .A3(new_n399), .A4(new_n426), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n405), .A2(new_n406), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n280), .A2(G223), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n432), .A2(new_n434), .B1(G33), .B2(G87), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n284), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n298), .B1(new_n222), .B2(new_n339), .ZN(new_n437));
  OAI21_X1  g0237(.A(G169), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n437), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n395), .A2(new_n399), .ZN(new_n440));
  INV_X1    g0240(.A(G87), .ZN(new_n441));
  OAI22_X1  g0241(.A1(new_n440), .A2(new_n433), .B1(new_n261), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n429), .B2(new_n430), .ZN(new_n443));
  OAI211_X1 g0243(.A(G179), .B(new_n439), .C1(new_n443), .C2(new_n284), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n438), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT18), .B1(new_n425), .B2(new_n446), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n402), .A2(KEYINPUT73), .A3(new_n403), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n409), .B1(new_n408), .B2(new_n410), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n419), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(new_n250), .A3(new_n424), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n378), .B1(new_n436), .B2(new_n437), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n344), .B(new_n439), .C1(new_n443), .C2(new_n284), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n451), .A2(new_n454), .A3(new_n390), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT17), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n451), .A2(new_n390), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT18), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n458), .A2(new_n459), .A3(new_n445), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n425), .A2(KEYINPUT17), .A3(new_n454), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n447), .A2(new_n457), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n245), .B1(new_n383), .B2(new_n463), .ZN(new_n464));
  NOR4_X1   g0264(.A1(new_n347), .A2(new_n462), .A3(KEYINPUT76), .A4(new_n382), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OR3_X1    g0266(.A1(new_n247), .A2(KEYINPUT25), .A3(G107), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT25), .B1(new_n247), .B2(G107), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n203), .A2(G33), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n247), .A2(new_n469), .A3(new_n210), .A4(new_n249), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n467), .B(new_n468), .C1(new_n217), .C2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n471), .B(KEYINPUT84), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT24), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT22), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(new_n441), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n399), .A2(new_n393), .A3(new_n394), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G116), .ZN(new_n477));
  AOI21_X1  g0277(.A(G20), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT23), .B1(new_n334), .B2(new_n204), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n204), .A2(G87), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n474), .B1(new_n285), .B2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT23), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n217), .A3(G20), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT83), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n482), .A2(new_n217), .A3(KEYINPUT83), .A4(G20), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n479), .A2(new_n481), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n473), .B1(new_n478), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n250), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n478), .A2(new_n488), .A3(new_n473), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n472), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT85), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n476), .A2(new_n477), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n204), .ZN(new_n495));
  INV_X1    g0295(.A(new_n488), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(KEYINPUT24), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(new_n250), .A3(new_n489), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT85), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n498), .A2(new_n499), .A3(new_n472), .ZN(new_n500));
  NOR2_X1   g0300(.A1(G250), .A2(G1698), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(new_n224), .B2(G1698), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n399), .A2(new_n502), .A3(new_n393), .A4(new_n394), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G294), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n288), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT86), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT5), .B(G41), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n289), .A2(G1), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n510), .A2(G264), .A3(new_n284), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n508), .A2(new_n284), .A3(G274), .A4(new_n509), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n506), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n284), .B1(new_n503), .B2(new_n504), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n511), .A2(new_n512), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT86), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(G169), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n515), .A2(new_n516), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(G179), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n518), .A2(KEYINPUT87), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT87), .B1(new_n518), .B2(new_n520), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n493), .B(new_n500), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT88), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n518), .A2(new_n520), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n518), .A2(KEYINPUT87), .A3(new_n520), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n498), .A2(new_n499), .A3(new_n472), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n499), .B1(new_n498), .B2(new_n472), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n533), .A3(KEYINPUT88), .ZN(new_n534));
  AOI21_X1  g0334(.A(G190), .B1(new_n514), .B2(new_n517), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n519), .A2(G200), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n472), .B(new_n498), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n525), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n247), .A2(G116), .ZN(new_n539));
  INV_X1    g0339(.A(new_n470), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n540), .B2(G116), .ZN(new_n541));
  AOI21_X1  g0341(.A(G20), .B1(new_n261), .B2(G97), .ZN(new_n542));
  NAND3_X1  g0342(.A1(KEYINPUT77), .A2(G33), .A3(G283), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT77), .B1(G33), .B2(G283), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(G116), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n249), .A2(new_n210), .B1(G20), .B2(new_n547), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n546), .A2(KEYINPUT20), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT20), .B1(new_n546), .B2(new_n548), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n541), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n552), .A2(new_n318), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n288), .B1(new_n509), .B2(new_n508), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G270), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n512), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(G257), .A2(G1698), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n218), .B2(G1698), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n395), .A2(new_n399), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n285), .A2(G303), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n284), .B1(new_n562), .B2(KEYINPUT81), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT81), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n564), .A3(new_n561), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n557), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n553), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n551), .A2(G169), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n563), .A2(new_n565), .ZN(new_n569));
  INV_X1    g0369(.A(new_n557), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n567), .B1(new_n571), .B2(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n570), .ZN(new_n573));
  INV_X1    g0373(.A(new_n568), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(KEYINPUT21), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT82), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT82), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n571), .A2(new_n577), .A3(KEYINPUT21), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n572), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n566), .A2(G190), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n580), .B(new_n552), .C1(new_n378), .C2(new_n566), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n284), .B1(G250), .B2(new_n509), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n289), .A2(G1), .A3(G274), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n280), .A2(G238), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n399), .A2(new_n393), .A3(new_n394), .A4(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT79), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n395), .A2(G244), .A3(G1698), .A4(new_n399), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n395), .A2(KEYINPUT79), .A3(new_n399), .A4(new_n585), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n588), .A2(new_n477), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n584), .B1(new_n591), .B2(new_n288), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G190), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n326), .A2(new_n247), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n470), .A2(new_n441), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT19), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n204), .B1(new_n361), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT80), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n332), .A2(new_n441), .A3(new_n223), .A4(new_n333), .ZN(new_n600));
  OAI211_X1 g0400(.A(KEYINPUT80), .B(new_n204), .C1(new_n361), .C2(new_n596), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n262), .A2(G97), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n596), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n204), .A2(G68), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n602), .B(new_n604), .C1(new_n440), .C2(new_n605), .ZN(new_n606));
  AOI211_X1 g0406(.A(new_n594), .B(new_n595), .C1(new_n606), .C2(new_n250), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n593), .B(new_n607), .C1(new_n378), .C2(new_n592), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n591), .A2(new_n288), .ZN(new_n609));
  INV_X1    g0409(.A(new_n584), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n318), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n594), .B1(new_n606), .B2(new_n250), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n325), .B2(new_n470), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n611), .B(new_n613), .C1(G169), .C2(new_n592), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n512), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(G257), .B2(new_n554), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT4), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n618), .A2(new_n216), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n619), .A2(new_n280), .A3(new_n275), .A4(new_n277), .ZN(new_n620));
  INV_X1    g0420(.A(new_n545), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n543), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n275), .A2(new_n277), .A3(G250), .A4(G1698), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n620), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n395), .A2(G244), .A3(new_n280), .A4(new_n399), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n624), .B1(new_n625), .B2(new_n618), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n617), .B1(new_n626), .B2(new_n284), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n316), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n335), .B1(new_n421), .B2(new_n422), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT6), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n630), .A2(new_n223), .A3(G107), .ZN(new_n631));
  XNOR2_X1  g0431(.A(G97), .B(G107), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n631), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  OAI22_X1  g0433(.A1(new_n633), .A2(new_n204), .B1(new_n215), .B2(new_n328), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n250), .B1(new_n629), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n247), .A2(G97), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n540), .B2(G97), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n617), .B(new_n318), .C1(new_n626), .C2(new_n284), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n628), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT78), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n378), .B1(new_n627), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n642), .B1(new_n641), .B2(new_n627), .ZN(new_n643));
  INV_X1    g0443(.A(new_n627), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n638), .B1(new_n644), .B2(G190), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n640), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n579), .A2(new_n581), .A3(new_n615), .A4(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n466), .A2(new_n538), .A3(new_n647), .ZN(G372));
  AND2_X1   g0448(.A1(new_n376), .A2(new_n342), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n457), .A2(new_n381), .A3(new_n461), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n447), .B(new_n460), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n320), .B1(new_n651), .B2(new_n314), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n607), .B1(new_n592), .B2(new_n378), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT89), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n607), .B(KEYINPUT89), .C1(new_n592), .C2(new_n378), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n593), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n640), .A3(new_n614), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT90), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT90), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n658), .A2(new_n662), .A3(new_n659), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n615), .A2(KEYINPUT26), .A3(new_n640), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n614), .ZN(new_n666));
  AND4_X1   g0466(.A1(new_n537), .A2(new_n646), .A3(new_n614), .A4(new_n657), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n526), .A2(new_n492), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n579), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n666), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n665), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n652), .B1(new_n466), .B2(new_n672), .ZN(G369));
  INV_X1    g0473(.A(new_n579), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n552), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n674), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n572), .ZN(new_n684));
  INV_X1    g0484(.A(new_n578), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n577), .B1(new_n571), .B2(KEYINPUT21), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n684), .B(new_n581), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n683), .B1(new_n687), .B2(new_n682), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT91), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT91), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n691), .A3(G330), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g0493(.A1(new_n531), .A2(new_n532), .A3(new_n681), .ZN(new_n694));
  OAI22_X1  g0494(.A1(new_n538), .A2(new_n694), .B1(new_n523), .B2(new_n681), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n525), .A2(new_n534), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n579), .A2(new_n680), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n537), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n526), .A2(new_n492), .A3(new_n681), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT92), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n699), .A2(KEYINPUT92), .A3(new_n700), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n696), .B1(new_n701), .B2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n207), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n600), .A2(G116), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n213), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT94), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n658), .A2(KEYINPUT26), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n608), .A2(new_n614), .A3(new_n640), .A4(new_n659), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT93), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n614), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n592), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n316), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(KEYINPUT93), .A3(new_n611), .A4(new_n613), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n714), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n525), .A2(new_n534), .A3(new_n579), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n667), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n712), .B1(new_n724), .B2(new_n681), .ZN(new_n725));
  AOI211_X1 g0525(.A(KEYINPUT94), .B(new_n680), .C1(new_n721), .C2(new_n723), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT29), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n680), .B1(new_n665), .B2(new_n670), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n643), .A2(new_n645), .ZN(new_n731));
  INV_X1    g0531(.A(new_n640), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(new_n608), .A4(new_n614), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n687), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n697), .A2(new_n537), .A3(new_n734), .A4(new_n681), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n506), .A2(G179), .A3(new_n511), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n627), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n566), .A3(new_n592), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT30), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n737), .A2(KEYINPUT30), .A3(new_n566), .A4(new_n592), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n519), .A2(G179), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n573), .A2(new_n717), .A3(new_n627), .A4(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n680), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n735), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G330), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n730), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n711), .B1(new_n754), .B2(G1), .ZN(G364));
  INV_X1    g0555(.A(G13), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n203), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n706), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n207), .A2(new_n278), .ZN(new_n761));
  INV_X1    g0561(.A(G355), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n762), .B1(G116), .B2(new_n207), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n440), .A2(new_n207), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT95), .Z(new_n765));
  NOR2_X1   g0565(.A1(new_n213), .A2(G45), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n243), .B2(G45), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n763), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT96), .Z(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n210), .B1(G20), .B2(new_n316), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n760), .B1(new_n768), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n204), .A2(G179), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(G190), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n441), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n318), .A2(new_n378), .A3(G190), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n778), .A2(new_n344), .A3(G200), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n783), .A2(new_n223), .B1(new_n784), .B2(new_n217), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n204), .A2(new_n318), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n344), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n780), .B(new_n785), .C1(G50), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G190), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n786), .A2(G190), .A3(new_n378), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n278), .B1(new_n791), .B2(new_n215), .C1(new_n221), .C2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT32), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n778), .A2(new_n790), .ZN(new_n795));
  INV_X1    g0595(.A(G159), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n795), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(KEYINPUT32), .A3(G159), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n793), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n787), .A2(G190), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n801), .A2(KEYINPUT97), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(KEYINPUT97), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n789), .B(new_n800), .C1(new_n264), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n804), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT99), .B(KEYINPUT33), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(G317), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n779), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n788), .A2(G326), .B1(new_n810), .B2(G303), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  INV_X1    g0612(.A(G294), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n811), .B1(new_n812), .B2(new_n784), .C1(new_n813), .C2(new_n783), .ZN(new_n814));
  INV_X1    g0614(.A(new_n792), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(G322), .B1(new_n798), .B2(G329), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n816), .B(new_n285), .C1(new_n817), .C2(new_n791), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n805), .A2(KEYINPUT98), .B1(new_n809), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(KEYINPUT98), .B2(new_n805), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n777), .B1(new_n821), .B2(new_n774), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n688), .B2(new_n772), .ZN(new_n823));
  INV_X1    g0623(.A(new_n760), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n688), .B2(G330), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n823), .B1(new_n693), .B2(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT100), .Z(G396));
  INV_X1    g0627(.A(new_n791), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n815), .A2(G143), .B1(new_n828), .B2(G159), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  INV_X1    g0630(.A(new_n788), .ZN(new_n831));
  INV_X1    g0631(.A(G150), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n829), .B1(new_n830), .B2(new_n831), .C1(new_n804), .C2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n834), .A2(KEYINPUT34), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n834), .A2(KEYINPUT34), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n432), .B1(new_n837), .B2(new_n795), .ZN(new_n838));
  INV_X1    g0638(.A(new_n784), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n839), .A2(G68), .B1(new_n782), .B2(G58), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n252), .B2(new_n779), .ZN(new_n841));
  NOR4_X1   g0641(.A1(new_n835), .A2(new_n836), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n784), .A2(new_n441), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n783), .A2(new_n223), .B1(new_n779), .B2(new_n217), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n843), .B(new_n844), .C1(G303), .C2(new_n788), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n791), .A2(new_n547), .B1(new_n795), .B2(new_n817), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n278), .B(new_n846), .C1(G294), .C2(new_n815), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n845), .B(new_n847), .C1(new_n812), .C2(new_n804), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT102), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n774), .B1(new_n842), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n774), .A2(new_n769), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT101), .Z(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n824), .B1(new_n853), .B2(new_n215), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n345), .B1(new_n330), .B2(new_n681), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n342), .ZN(new_n856));
  OR2_X1    g0656(.A1(new_n342), .A2(new_n680), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n850), .B(new_n854), .C1(new_n859), .C2(new_n770), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT103), .B1(new_n728), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n728), .B2(new_n859), .ZN(new_n862));
  INV_X1    g0662(.A(new_n728), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(KEYINPUT103), .A3(new_n858), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n752), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n824), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n752), .B1(new_n862), .B2(new_n864), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n860), .B1(new_n866), .B2(new_n867), .ZN(G384));
  NAND2_X1  g0668(.A1(new_n458), .A2(new_n445), .ZN(new_n869));
  INV_X1    g0669(.A(new_n678), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n458), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n871), .A3(new_n455), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT37), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n869), .A2(new_n871), .A3(new_n874), .A4(new_n455), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n462), .A2(new_n458), .A3(new_n870), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT105), .ZN(new_n880));
  INV_X1    g0680(.A(new_n417), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n448), .B2(new_n449), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n418), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n391), .B1(new_n883), .B2(new_n420), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n455), .B1(new_n884), .B2(new_n678), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n446), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n884), .A2(new_n678), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n875), .A2(new_n887), .B1(new_n462), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n880), .B1(new_n889), .B2(KEYINPUT38), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n887), .A2(new_n875), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n462), .A2(new_n888), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n891), .A2(new_n892), .A3(new_n880), .A4(KEYINPUT38), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n879), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n375), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n373), .A3(new_n372), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n357), .B(new_n680), .C1(new_n897), .C2(new_n380), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n357), .A2(new_n680), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n376), .A2(new_n381), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n858), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n751), .A2(KEYINPUT40), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n895), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n538), .A2(new_n647), .A3(new_n680), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n901), .B1(new_n905), .B2(new_n749), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n891), .A2(new_n892), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT38), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n904), .B1(KEYINPUT40), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n314), .A2(new_n321), .ZN(new_n913));
  INV_X1    g0713(.A(new_n382), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(new_n914), .A3(new_n346), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT76), .B1(new_n915), .B2(new_n462), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n383), .A2(new_n245), .A3(new_n463), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n751), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n912), .A2(new_n919), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n920), .A2(G330), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n870), .B1(new_n447), .B2(new_n460), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n898), .A2(new_n900), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n671), .A2(new_n681), .A3(new_n859), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n925), .B1(new_n926), .B2(new_n857), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n909), .A2(new_n910), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n897), .A2(new_n357), .A3(new_n681), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n909), .A2(KEYINPUT39), .A3(new_n910), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n910), .A2(KEYINPUT105), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n878), .B1(new_n933), .B2(new_n893), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n931), .B(new_n932), .C1(new_n934), .C2(KEYINPUT39), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n727), .A2(new_n729), .A3(new_n918), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n652), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n936), .B(new_n938), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n922), .A2(new_n939), .B1(new_n203), .B2(new_n757), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT106), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n922), .A2(new_n939), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n633), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n547), .B(new_n212), .C1(new_n946), .C2(KEYINPUT35), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(KEYINPUT35), .B2(new_n946), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT36), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n413), .A2(new_n213), .A3(new_n215), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n950), .A2(KEYINPUT104), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n950), .A2(KEYINPUT104), .B1(G50), .B2(new_n264), .ZN(new_n952));
  OAI211_X1 g0752(.A(G1), .B(new_n756), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n945), .A2(new_n949), .A3(new_n953), .ZN(G367));
  INV_X1    g0754(.A(new_n765), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n235), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n775), .B1(new_n207), .B2(new_n325), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n760), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n806), .A2(G159), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n791), .A2(new_n252), .B1(new_n795), .B2(new_n830), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n285), .B(new_n960), .C1(G150), .C2(new_n815), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n839), .A2(G77), .B1(new_n782), .B2(G68), .ZN(new_n962));
  AOI22_X1  g0762(.A1(new_n788), .A2(G143), .B1(new_n810), .B2(G58), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n959), .A2(new_n961), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n806), .A2(G294), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n782), .A2(new_n334), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n788), .A2(G311), .B1(new_n839), .B2(G97), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n965), .A2(new_n440), .A3(new_n966), .A4(new_n967), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n815), .A2(G303), .B1(new_n828), .B2(G283), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n810), .A2(KEYINPUT46), .A3(G116), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT46), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n779), .B2(new_n547), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n798), .A2(G317), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n969), .A2(new_n970), .A3(new_n972), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n964), .B1(new_n968), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n958), .B1(new_n976), .B2(new_n774), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n657), .B(new_n614), .C1(new_n607), .C2(new_n681), .ZN(new_n978));
  OR3_X1    g0778(.A1(new_n614), .A2(new_n607), .A3(new_n681), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n977), .B1(new_n980), .B2(new_n772), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT109), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n699), .A2(new_n700), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT92), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n638), .A2(new_n680), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n646), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n640), .A2(new_n680), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n985), .A2(new_n702), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n993));
  INV_X1    g0793(.A(new_n991), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n985), .A2(new_n702), .A3(new_n989), .A4(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n989), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n703), .B2(new_n701), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT45), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g0800(.A(KEYINPUT45), .B(new_n997), .C1(new_n703), .C2(new_n701), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n996), .A2(new_n1002), .A3(new_n696), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n696), .B1(new_n996), .B2(new_n1002), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n699), .B1(new_n695), .B2(new_n698), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n693), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n693), .A2(new_n1007), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n753), .B1(new_n1006), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n706), .B(KEYINPUT41), .Z(new_n1012));
  OAI21_X1  g0812(.A(new_n758), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n525), .A2(new_n534), .B1(new_n643), .B2(new_n645), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n681), .B1(new_n1014), .B2(new_n640), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n699), .A2(new_n989), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT42), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1015), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT107), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1018), .A2(new_n1019), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n1020), .A2(new_n1021), .B1(KEYINPUT43), .B2(new_n980), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(KEYINPUT43), .B2(new_n980), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n693), .A2(new_n695), .A3(new_n997), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT43), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n980), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1020), .A2(new_n1021), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1023), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1025), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n982), .B1(new_n1013), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1005), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n753), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n1034), .A3(new_n1003), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1012), .B1(new_n1035), .B2(new_n754), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1031), .B(new_n982), .C1(new_n1036), .C2(new_n759), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n981), .B1(new_n1032), .B2(new_n1038), .ZN(G387));
  NAND2_X1  g0839(.A1(new_n1010), .A2(new_n759), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n695), .A2(new_n772), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n765), .B1(new_n289), .B2(new_n232), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n708), .B2(new_n761), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n255), .A2(G50), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT50), .ZN(new_n1045));
  AOI21_X1  g0845(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1045), .A2(new_n708), .A3(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1043), .A2(new_n1047), .B1(new_n217), .B2(new_n705), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n760), .B1(new_n1048), .B2(new_n776), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n806), .A2(new_n384), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n779), .A2(new_n215), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n783), .A2(new_n325), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(G159), .C2(new_n788), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n791), .A2(new_n264), .B1(new_n795), .B2(new_n832), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G50), .B2(new_n815), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n440), .B1(G97), .B2(new_n839), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1050), .A2(new_n1053), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n432), .B1(G326), .B2(new_n798), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n815), .A2(G317), .B1(new_n828), .B2(G303), .ZN(new_n1059));
  INV_X1    g0859(.A(G322), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1059), .B1(new_n1060), .B2(new_n831), .C1(new_n804), .C2(new_n817), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n810), .A2(G294), .B1(new_n782), .B2(G283), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT49), .Z(new_n1067));
  INV_X1    g0867(.A(KEYINPUT110), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1058), .B1(new_n547), .B2(new_n784), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1057), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1049), .B1(new_n1071), .B2(new_n774), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT111), .Z(new_n1073));
  INV_X1    g0873(.A(new_n1034), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n706), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n754), .A2(new_n1010), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1040), .B1(new_n1041), .B2(new_n1073), .C1(new_n1075), .C2(new_n1076), .ZN(G393));
  OAI21_X1  g0877(.A(new_n1074), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1078), .A2(new_n1035), .A3(new_n706), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1006), .A2(new_n759), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n774), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G317), .A2(new_n788), .B1(new_n815), .B2(G311), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT52), .Z(new_n1083));
  OAI22_X1  g0883(.A1(new_n779), .A2(new_n812), .B1(new_n795), .B2(new_n1060), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT112), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n806), .A2(G303), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n285), .B1(new_n791), .B2(new_n813), .C1(new_n217), .C2(new_n784), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(G116), .B2(new_n782), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n831), .A2(new_n832), .B1(new_n796), .B2(new_n792), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT51), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n806), .A2(G50), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n791), .A2(new_n255), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n1093), .B(new_n440), .C1(G143), .C2(new_n798), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n779), .A2(new_n264), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n843), .B(new_n1095), .C1(G77), .C2(new_n782), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1081), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n765), .A2(new_n240), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n776), .B1(G97), .B2(new_n705), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n824), .B(new_n1098), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n997), .B2(new_n772), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1079), .A2(new_n1080), .A3(new_n1102), .ZN(G390));
  OAI21_X1  g0903(.A(new_n932), .B1(new_n934), .B2(KEYINPUT39), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n769), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n810), .A2(G150), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT53), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n285), .B1(new_n798), .B2(G125), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT54), .B(G143), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1108), .B1(new_n791), .B2(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n783), .A2(new_n796), .B1(new_n784), .B2(new_n252), .ZN(new_n1111));
  OR3_X1    g0911(.A1(new_n1107), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(G128), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n831), .A2(new_n1113), .B1(new_n837), .B2(new_n792), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT116), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1112), .B(new_n1115), .C1(G137), .C2(new_n806), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(KEYINPUT117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n806), .A2(new_n334), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n791), .A2(new_n223), .B1(new_n795), .B2(new_n813), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n278), .B(new_n1120), .C1(G116), .C2(new_n815), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n780), .B1(G68), .B2(new_n839), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n788), .A2(G283), .B1(G77), .B2(new_n782), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1119), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT117), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1124), .B1(new_n1116), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n774), .B1(new_n1118), .B2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n824), .B1(new_n853), .B2(new_n389), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1105), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n857), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n728), .B2(new_n859), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n930), .B1(new_n1131), .B2(new_n925), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1104), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n713), .A2(new_n720), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n667), .B2(new_n722), .ZN(new_n1135));
  OAI21_X1  g0935(.A(KEYINPUT94), .B1(new_n1135), .B2(new_n680), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n724), .A2(new_n712), .A3(new_n681), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n1137), .A3(new_n857), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1138), .A2(new_n856), .A3(new_n924), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n934), .A2(new_n931), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1133), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(G330), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n735), .B2(new_n750), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n1144), .A2(new_n859), .A3(new_n924), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1144), .A2(new_n859), .A3(new_n924), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1133), .A2(new_n1141), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1129), .B1(new_n1149), .B2(new_n758), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT115), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1148), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1147), .B1(new_n1133), .B2(new_n1141), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT113), .B1(new_n466), .B2(new_n752), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT113), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n918), .A2(new_n1156), .A3(new_n1144), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1158), .A2(new_n652), .A3(new_n937), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n924), .B1(new_n1144), .B2(new_n859), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1145), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1138), .A2(new_n856), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT114), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1131), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n925), .B1(new_n752), .B2(new_n858), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n1147), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1163), .A2(new_n1164), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1161), .A2(new_n1162), .A3(KEYINPUT114), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1159), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1151), .B1(new_n1154), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n725), .A2(new_n726), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1172), .A2(new_n857), .B1(new_n342), .B2(new_n855), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1164), .B1(new_n1173), .B2(new_n1167), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1167), .A2(new_n1165), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1174), .A2(new_n1169), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1159), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1149), .A2(new_n1178), .A3(KEYINPUT115), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1171), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n707), .B1(new_n1154), .B2(new_n1170), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1150), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(G378));
  OAI21_X1  g0983(.A(G330), .B1(new_n911), .B2(KEYINPUT40), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n933), .A2(new_n893), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n902), .B1(new_n1185), .B2(new_n879), .ZN(new_n1186));
  OAI21_X1  g0986(.A(KEYINPUT120), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n891), .A2(new_n892), .A3(KEYINPUT38), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT38), .B1(new_n891), .B2(new_n892), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n751), .B(new_n901), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT40), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1143), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT120), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1192), .A2(new_n904), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n913), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n315), .A2(new_n678), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT55), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1195), .B(new_n1198), .ZN(new_n1199));
  XOR2_X1   g0999(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1200));
  AND2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1187), .A2(new_n1194), .A3(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1203), .A2(new_n1193), .A3(new_n904), .A4(new_n1192), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(KEYINPUT121), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT122), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n929), .B2(new_n935), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n929), .A2(new_n1208), .A3(new_n935), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1207), .A2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1207), .A2(new_n1212), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n759), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1203), .A2(new_n769), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n760), .B1(new_n852), .B2(G50), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n791), .A2(new_n325), .B1(new_n795), .B2(new_n812), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n440), .A2(new_n283), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(G107), .C2(new_n815), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n784), .A2(new_n221), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n783), .A2(new_n264), .B1(new_n779), .B2(new_n215), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(G116), .C2(new_n788), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1220), .B(new_n1223), .C1(new_n223), .C2(new_n804), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT58), .ZN(new_n1225));
  AOI21_X1  g1025(.A(G50), .B1(new_n261), .B2(new_n283), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1224), .A2(new_n1225), .B1(new_n1219), .B2(new_n1226), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n792), .A2(new_n1113), .B1(new_n791), .B2(new_n830), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1109), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1228), .B1(new_n810), .B2(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n788), .A2(G125), .B1(G150), .B2(new_n782), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n804), .C2(new_n837), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(KEYINPUT59), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n839), .A2(G159), .ZN(new_n1235));
  AOI211_X1 g1035(.A(G33), .B(G41), .C1(new_n798), .C2(G124), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1227), .B1(new_n1225), .B2(new_n1224), .C1(new_n1233), .C2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1217), .B1(new_n1238), .B2(new_n774), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1216), .A2(new_n1239), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT119), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1215), .A2(KEYINPUT123), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT123), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n929), .A2(new_n1208), .A3(new_n935), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1245), .A2(new_n1209), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1246), .A2(KEYINPUT121), .A3(new_n1206), .A4(new_n1205), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1207), .A2(new_n1212), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n758), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1244), .B1(new_n1249), .B2(new_n1241), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1243), .A2(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1146), .A2(new_n1176), .A3(new_n1148), .A4(new_n1177), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1177), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT57), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n936), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1205), .A2(new_n1257), .A3(new_n1206), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1257), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n1255), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n707), .B1(new_n1260), .B2(new_n1253), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1256), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1251), .A2(new_n1262), .ZN(G375));
  AOI21_X1  g1063(.A(new_n758), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n925), .A2(new_n769), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n760), .B1(new_n852), .B2(G68), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n831), .A2(new_n813), .B1(new_n779), .B2(new_n223), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1052), .B(new_n1267), .C1(G77), .C2(new_n839), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n335), .A2(new_n791), .B1(new_n792), .B2(new_n812), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n278), .B(new_n1269), .C1(G303), .C2(new_n798), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1268), .B(new_n1270), .C1(new_n547), .C2(new_n804), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n779), .A2(new_n796), .B1(new_n795), .B2(new_n1113), .ZN(new_n1272));
  XOR2_X1   g1072(.A(new_n1272), .B(KEYINPUT124), .Z(new_n1273));
  NOR2_X1   g1073(.A1(new_n783), .A2(new_n252), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1221), .B(new_n1274), .C1(G132), .C2(new_n788), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n792), .A2(new_n830), .B1(new_n791), .B2(new_n832), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(new_n440), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1275), .B(new_n1277), .C1(new_n804), .C2(new_n1109), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1271), .B1(new_n1273), .B2(new_n1278), .ZN(new_n1279));
  OR2_X1    g1079(.A1(new_n1279), .A2(KEYINPUT125), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1081), .B1(new_n1279), .B2(KEYINPUT125), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1266), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1265), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT126), .B1(new_n1264), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1176), .A2(new_n759), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT126), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n1287), .A3(new_n1283), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1012), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1159), .A2(new_n1174), .A3(new_n1169), .A4(new_n1175), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1178), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1292), .ZN(G381));
  AOI22_X1  g1093(.A1(new_n1243), .A2(new_n1250), .B1(new_n1256), .B2(new_n1261), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1182), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1031), .B1(new_n1036), .B2(new_n759), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT109), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1037), .ZN(new_n1298));
  INV_X1    g1098(.A(G390), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1298), .A2(new_n981), .A3(new_n1299), .ZN(new_n1300));
  OR4_X1    g1100(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1301));
  OR3_X1    g1101(.A1(new_n1295), .A2(new_n1300), .A3(new_n1301), .ZN(G407));
  OAI211_X1 g1102(.A(G407), .B(G213), .C1(G343), .C2(new_n1295), .ZN(G409));
  AND2_X1   g1103(.A1(new_n679), .A2(G213), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n936), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1205), .A2(new_n1257), .A3(new_n1206), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(new_n759), .A3(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1242), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1247), .A2(new_n1248), .B1(new_n1252), .B2(new_n1177), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1309), .B1(new_n1290), .B2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1304), .B1(new_n1311), .B2(new_n1182), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1312), .B1(new_n1294), .B2(new_n1182), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1291), .A2(KEYINPUT60), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT60), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1168), .A2(new_n1315), .A3(new_n1159), .A4(new_n1169), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1317), .A2(new_n706), .A3(new_n1178), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1318), .A2(new_n1289), .A3(G384), .ZN(new_n1319));
  AOI21_X1  g1119(.A(G384), .B1(new_n1318), .B2(new_n1289), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1304), .A2(G2897), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1319), .A2(new_n1320), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(G384), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1287), .B1(new_n1286), .B2(new_n1283), .ZN(new_n1325));
  AOI211_X1 g1125(.A(KEYINPUT126), .B(new_n1284), .C1(new_n1176), .C2(new_n759), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1178), .A2(new_n706), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1328), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1324), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1318), .A2(new_n1289), .A3(G384), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1321), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1323), .A2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT61), .B1(new_n1313), .B2(new_n1333), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1312), .B(new_n1335), .C1(new_n1294), .C2(new_n1182), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(KEYINPUT62), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(G375), .A2(G378), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT62), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1338), .A2(new_n1339), .A3(new_n1312), .A4(new_n1335), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1334), .A2(new_n1337), .A3(new_n1340), .ZN(new_n1341));
  XOR2_X1   g1141(.A(G393), .B(G396), .Z(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1299), .B1(new_n1298), .B2(new_n981), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n981), .ZN(new_n1345));
  AOI211_X1 g1145(.A(new_n1345), .B(G390), .C1(new_n1297), .C2(new_n1037), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1343), .B1(new_n1344), .B2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(G387), .A2(G390), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1348), .A2(new_n1300), .A3(new_n1342), .ZN(new_n1349));
  AND2_X1   g1149(.A1(new_n1347), .A2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1341), .A2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1347), .A2(new_n1349), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT63), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1336), .A2(new_n1353), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1338), .A2(KEYINPUT63), .A3(new_n1312), .A4(new_n1335), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1352), .A2(new_n1334), .A3(new_n1354), .A4(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1351), .A2(new_n1356), .ZN(G405));
  NAND2_X1  g1157(.A1(new_n1338), .A2(new_n1295), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1335), .ZN(new_n1359));
  OAI211_X1 g1159(.A(new_n1338), .B(new_n1295), .C1(new_n1320), .C2(new_n1319), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1352), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1350), .A2(new_n1359), .A3(new_n1360), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1362), .A2(new_n1363), .ZN(G402));
endmodule


