//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n188));
  INV_X1    g002(.A(G137), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT66), .B1(new_n189), .B2(G134), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT66), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G137), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G134), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT1), .B1(new_n199), .B2(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G128), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n201), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n203), .A2(new_n204), .A3(new_n207), .A4(G128), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n198), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  AOI22_X1  g025(.A1(KEYINPUT65), .A2(new_n211), .B1(new_n192), .B2(G137), .ZN(new_n212));
  OAI22_X1  g026(.A1(KEYINPUT65), .A2(new_n211), .B1(new_n192), .B2(G137), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n215), .A2(new_n189), .A3(KEYINPUT11), .A4(G134), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n197), .B1(new_n196), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n188), .B1(new_n210), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n196), .A2(new_n217), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n196), .A2(new_n197), .B1(new_n206), .B2(new_n208), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(KEYINPUT69), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(KEYINPUT2), .A2(G113), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n224), .B(KEYINPUT68), .ZN(new_n225));
  OR2_X1    g039(.A1(KEYINPUT2), .A2(G113), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G116), .B(G119), .ZN(new_n228));
  XNOR2_X1  g042(.A(new_n227), .B(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n212), .A2(new_n213), .A3(new_n216), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G131), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n217), .ZN(new_n232));
  XNOR2_X1  g046(.A(G143), .B(G146), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT0), .ZN(new_n234));
  INV_X1    g048(.A(G128), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT0), .B(G128), .Z(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n219), .A2(new_n223), .A3(new_n229), .A4(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G237), .ZN(new_n241));
  INV_X1    g055(.A(G953), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n241), .A2(new_n242), .A3(G210), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n243), .B(KEYINPUT71), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT26), .B(G101), .Z(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n221), .A2(new_n222), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n237), .A2(new_n233), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n234), .A2(new_n235), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n205), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n236), .B(KEYINPUT64), .C1(new_n233), .C2(new_n237), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n232), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT30), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n250), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n219), .A2(new_n239), .A3(new_n223), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n259), .B1(KEYINPUT30), .B2(new_n260), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n240), .B(new_n249), .C1(new_n261), .C2(new_n229), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n187), .B1(new_n262), .B2(KEYINPUT31), .ZN(new_n263));
  INV_X1    g077(.A(new_n240), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(KEYINPUT30), .ZN(new_n265));
  INV_X1    g079(.A(new_n259), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n227), .B(new_n228), .Z(new_n268));
  AOI21_X1  g082(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT31), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n269), .A2(KEYINPUT72), .A3(new_n270), .A4(new_n249), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n263), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n250), .A2(new_n257), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n268), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n275), .B2(new_n240), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n250), .A2(new_n229), .A3(new_n239), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n277), .A2(new_n273), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AOI22_X1  g093(.A1(new_n279), .A2(new_n248), .B1(new_n262), .B2(KEYINPUT31), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(G472), .A2(G902), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT32), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(KEYINPUT73), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT73), .ZN(new_n286));
  INV_X1    g100(.A(new_n282), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n272), .B2(new_n280), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n286), .B1(new_n288), .B2(KEYINPUT32), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n260), .A2(new_n268), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n240), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n278), .B1(new_n292), .B2(KEYINPUT28), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n248), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(G902), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n269), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n248), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n294), .B1(new_n279), .B2(new_n248), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G472), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n288), .A2(KEYINPUT32), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT74), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n288), .A2(new_n305), .A3(KEYINPUT32), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n290), .A2(new_n302), .A3(new_n304), .A4(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT22), .B(G137), .Z(new_n309));
  NAND3_X1  g123(.A1(new_n242), .A2(G221), .A3(G234), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n235), .A2(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(KEYINPUT75), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n235), .A2(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(KEYINPUT23), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n312), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT24), .B(G110), .Z(new_n320));
  OAI22_X1  g134(.A1(new_n317), .A2(G110), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n322), .A2(KEYINPUT16), .A3(G140), .ZN(new_n323));
  XNOR2_X1  g137(.A(G125), .B(G140), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(KEYINPUT16), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G146), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n202), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n325), .B(G146), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n317), .A2(G110), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n319), .A2(new_n320), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n311), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n335), .B1(new_n334), .B2(new_n333), .ZN(new_n336));
  AOI211_X1 g150(.A(KEYINPUT76), .B(new_n311), .C1(new_n328), .C2(new_n332), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n308), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT25), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G217), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(G234), .B2(new_n308), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n336), .A2(new_n337), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n342), .A2(G902), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(G125), .B1(new_n206), .B2(new_n208), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(G125), .B2(new_n238), .ZN(new_n350));
  INV_X1    g164(.A(G224), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(G953), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n350), .B(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n354));
  INV_X1    g168(.A(G107), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n355), .A3(G104), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(KEYINPUT3), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n355), .A2(G104), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n354), .A2(new_n360), .A3(new_n355), .A4(G104), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT79), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT4), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n362), .A2(G101), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(G101), .ZN(new_n366));
  INV_X1    g180(.A(G101), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n357), .A2(new_n367), .A3(new_n359), .A4(new_n361), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n366), .A2(new_n363), .A3(KEYINPUT4), .A4(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n268), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n225), .A2(new_n226), .A3(new_n228), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n228), .A2(KEYINPUT5), .ZN(new_n372));
  INV_X1    g186(.A(G116), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n373), .A2(KEYINPUT5), .A3(G119), .ZN(new_n374));
  INV_X1    g188(.A(G113), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n371), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n355), .A2(G104), .ZN(new_n378));
  OAI21_X1  g192(.A(G101), .B1(new_n378), .B2(new_n358), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n368), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n370), .A2(new_n382), .ZN(new_n383));
  XOR2_X1   g197(.A(G110), .B(G122), .Z(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n384), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n370), .A2(new_n382), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(KEYINPUT6), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n386), .B1(new_n370), .B2(new_n382), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n391));
  AND3_X1   g205(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n390), .B1(new_n389), .B2(new_n391), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n353), .B(new_n388), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n377), .A2(new_n380), .ZN(new_n395));
  XOR2_X1   g209(.A(new_n384), .B(KEYINPUT8), .Z(new_n396));
  OR2_X1    g210(.A1(new_n376), .A2(KEYINPUT88), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n376), .A2(KEYINPUT88), .B1(KEYINPUT5), .B2(new_n228), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n371), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n395), .B(new_n396), .C1(new_n380), .C2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT7), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n352), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT89), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n403), .ZN(new_n405));
  OR3_X1    g219(.A1(new_n350), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n405), .B1(new_n350), .B2(new_n404), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n387), .A2(new_n400), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n394), .A2(new_n308), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G210), .B1(G237), .B2(G902), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n394), .A2(new_n308), .A3(new_n410), .A4(new_n408), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G214), .B1(G237), .B2(G902), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(G128), .B(G143), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT13), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n199), .A2(G128), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n418), .B(G134), .C1(KEYINPUT13), .C2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G116), .B(G122), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(new_n355), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n417), .A2(new_n192), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n417), .B(new_n192), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n373), .A2(KEYINPUT14), .A3(G122), .ZN(new_n426));
  INV_X1    g240(.A(new_n421), .ZN(new_n427));
  OAI211_X1 g241(.A(G107), .B(new_n426), .C1(new_n427), .C2(KEYINPUT14), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n421), .A2(new_n355), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n425), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT9), .B(G234), .Z(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(G217), .A3(new_n242), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n431), .A2(new_n433), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n308), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G478), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(KEYINPUT15), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n438), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT93), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(KEYINPUT93), .B(new_n308), .C1(new_n434), .C2(new_n435), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT94), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT94), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  AND2_X1   g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n242), .A2(G952), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(G234), .B2(G237), .ZN(new_n453));
  XOR2_X1   g267(.A(KEYINPUT21), .B(G898), .Z(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  AOI211_X1 g269(.A(new_n308), .B(new_n242), .C1(G234), .C2(G237), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G113), .B(G122), .ZN(new_n458));
  XNOR2_X1  g272(.A(KEYINPUT91), .B(G104), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n329), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n241), .A2(new_n242), .A3(G214), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT90), .B(G143), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n462), .B1(KEYINPUT90), .B2(new_n199), .ZN(new_n466));
  OAI21_X1  g280(.A(G131), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT17), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n465), .A2(new_n466), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n214), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n467), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n461), .B(new_n469), .C1(new_n472), .C2(KEYINPUT17), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n468), .A2(KEYINPUT18), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT18), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n324), .B(new_n202), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n474), .A2(new_n476), .A3(new_n477), .A4(new_n471), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n460), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  XOR2_X1   g293(.A(new_n324), .B(KEYINPUT19), .Z(new_n480));
  OAI211_X1 g294(.A(new_n472), .B(new_n326), .C1(G146), .C2(new_n480), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n481), .A2(new_n478), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n479), .B1(new_n460), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT20), .ZN(new_n484));
  INV_X1    g298(.A(G475), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .A4(new_n308), .ZN(new_n486));
  INV_X1    g300(.A(new_n479), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n481), .A2(new_n478), .A3(new_n460), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n487), .A2(new_n485), .A3(new_n308), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT20), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n473), .A2(new_n478), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n460), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n494), .B1(new_n491), .B2(new_n493), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n486), .A2(new_n490), .B1(G475), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NOR4_X1   g311(.A1(new_n416), .A2(new_n451), .A3(new_n457), .A4(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(G221), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n499), .B1(new_n432), .B2(new_n308), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n242), .A2(G227), .ZN(new_n501));
  XOR2_X1   g315(.A(new_n501), .B(G140), .Z(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT77), .B(G110), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n232), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT80), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n208), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n233), .A2(KEYINPUT80), .A3(new_n207), .A4(G128), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT81), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n235), .B1(new_n200), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n203), .A2(KEYINPUT81), .A3(KEYINPUT1), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n233), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT82), .B1(new_n514), .B2(new_n380), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n200), .A2(new_n510), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(G128), .A3(new_n512), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n205), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n507), .A3(new_n508), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT82), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n520), .A3(new_n381), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n381), .A2(new_n209), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n505), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT84), .B1(new_n525), .B2(KEYINPUT12), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n523), .B1(new_n515), .B2(new_n521), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT84), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n529));
  NOR4_X1   g343(.A1(new_n527), .A2(new_n528), .A3(new_n529), .A4(new_n505), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n514), .A2(KEYINPUT82), .A3(new_n380), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n520), .B1(new_n519), .B2(new_n381), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n524), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT12), .B1(new_n533), .B2(new_n232), .ZN(new_n534));
  NOR3_X1   g348(.A1(new_n526), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n522), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n369), .A2(new_n238), .A3(new_n365), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n381), .A2(KEYINPUT10), .A3(new_n209), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n537), .A2(new_n505), .A3(new_n538), .A4(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n504), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n543), .A2(new_n232), .ZN(new_n544));
  INV_X1    g358(.A(new_n504), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n540), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n542), .A2(KEYINPUT85), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT85), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n533), .A2(KEYINPUT12), .A3(new_n232), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n528), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n529), .B1(new_n527), .B2(new_n505), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n525), .A2(KEYINPUT84), .A3(KEYINPUT12), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n545), .B1(new_n555), .B2(new_n540), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n550), .B1(new_n556), .B2(new_n547), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n549), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G469), .B1(new_n558), .B2(G902), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT86), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n546), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n540), .A2(KEYINPUT86), .A3(new_n545), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n555), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n504), .B1(new_n544), .B2(new_n541), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G469), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n308), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n500), .B1(new_n559), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n307), .A2(new_n348), .A3(new_n498), .A4(new_n568), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT95), .B(G101), .Z(new_n570));
  XNOR2_X1  g384(.A(new_n569), .B(new_n570), .ZN(G3));
  AOI21_X1  g385(.A(G902), .B1(new_n272), .B2(new_n280), .ZN(new_n572));
  INV_X1    g386(.A(G472), .ZN(new_n573));
  OAI22_X1  g387(.A1(KEYINPUT96), .A2(new_n288), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n281), .A2(new_n308), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT96), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(G472), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n559), .A2(new_n567), .ZN(new_n580));
  INV_X1    g394(.A(new_n500), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n348), .A4(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT33), .ZN(new_n583));
  OR3_X1    g397(.A1(new_n434), .A2(new_n435), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n583), .B1(new_n434), .B2(new_n435), .ZN(new_n585));
  AND4_X1   g399(.A1(G478), .A2(new_n584), .A3(new_n308), .A4(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(G478), .B1(new_n443), .B2(new_n444), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n496), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n416), .A2(new_n457), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n582), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT97), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT34), .B(G104), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(G6));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n486), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n487), .A2(new_n485), .A3(new_n488), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n599), .A2(KEYINPUT98), .A3(new_n484), .A4(new_n308), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n598), .A2(new_n600), .A3(new_n490), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n448), .A2(new_n601), .A3(new_n450), .ZN(new_n602));
  INV_X1    g416(.A(new_n457), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n495), .A2(G475), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n602), .A2(KEYINPUT99), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n415), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n412), .B2(new_n413), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n448), .A2(new_n601), .A3(new_n604), .A4(new_n450), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n608), .B1(new_n609), .B2(new_n457), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n605), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n582), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT100), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT35), .B(G107), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  NOR2_X1   g430(.A1(new_n311), .A2(KEYINPUT36), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n333), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n345), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n343), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n498), .A2(new_n568), .A3(new_n579), .A4(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT37), .B(G110), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G12));
  INV_X1    g437(.A(G900), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n456), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n453), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n495), .B2(G475), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n602), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n416), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n307), .A2(new_n631), .A3(new_n568), .A4(new_n620), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G128), .ZN(G30));
  XOR2_X1   g447(.A(new_n627), .B(KEYINPUT39), .Z(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n568), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT40), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n412), .A2(new_n413), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n638), .B1(new_n412), .B2(new_n413), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n451), .A2(new_n497), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n568), .A2(new_n644), .A3(new_n635), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n637), .A2(new_n641), .A3(new_n643), .A4(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n269), .A2(new_n248), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n308), .B1(new_n292), .B2(new_n249), .ZN(new_n648));
  OAI21_X1  g462(.A(G472), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n290), .A2(new_n304), .A3(new_n306), .A4(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n620), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(new_n415), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n199), .ZN(G45));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n496), .A2(new_n588), .A3(new_n628), .ZN(new_n656));
  AND3_X1   g470(.A1(new_n607), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n655), .B1(new_n607), .B2(new_n656), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n307), .A2(new_n659), .A3(new_n568), .A4(new_n620), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G146), .ZN(G48));
  NAND2_X1  g475(.A1(new_n565), .A2(new_n308), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(G469), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n567), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n500), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n307), .A2(new_n348), .A3(new_n591), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT41), .B(G113), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G15));
  NAND4_X1  g482(.A1(new_n611), .A2(new_n307), .A3(new_n348), .A4(new_n665), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT103), .B(G116), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G18));
  NAND4_X1  g485(.A1(new_n307), .A2(new_n498), .A3(new_n620), .A4(new_n665), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G119), .ZN(G21));
  INV_X1    g487(.A(new_n262), .ZN(new_n674));
  OAI221_X1 g488(.A(new_n272), .B1(new_n270), .B2(new_n674), .C1(new_n249), .C2(new_n293), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT104), .B(G472), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n282), .A2(new_n675), .B1(new_n575), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n348), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n416), .A2(new_n457), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n679), .A3(new_n643), .A4(new_n665), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G122), .ZN(G24));
  AND2_X1   g495(.A1(new_n677), .A2(new_n620), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n682), .A2(new_n607), .A3(new_n656), .A4(new_n665), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G125), .ZN(G27));
  AND2_X1   g498(.A1(new_n303), .A2(new_n302), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n283), .A2(new_n284), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n347), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n556), .A2(new_n547), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(G469), .ZN(new_n689));
  NAND2_X1  g503(.A1(G469), .A2(G902), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT105), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n689), .A2(new_n567), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n581), .ZN(new_n693));
  INV_X1    g507(.A(new_n656), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n414), .A2(new_n606), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n687), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n698));
  INV_X1    g512(.A(new_n693), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n307), .A2(new_n348), .A3(new_n696), .A4(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n694), .A2(KEYINPUT42), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n698), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n214), .ZN(G33));
  XNOR2_X1  g518(.A(new_n630), .B(KEYINPUT106), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n192), .ZN(G36));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n549), .A2(new_n557), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n566), .B1(new_n688), .B2(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(KEYINPUT46), .A3(new_n691), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n567), .ZN(new_n713));
  INV_X1    g527(.A(new_n691), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n709), .B2(new_n710), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(KEYINPUT46), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n581), .B(new_n635), .C1(new_n713), .C2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n711), .A2(new_n691), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n567), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n715), .B2(KEYINPUT46), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(KEYINPUT107), .A3(new_n581), .A4(new_n635), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n719), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n696), .B(KEYINPUT109), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n586), .A2(new_n587), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n496), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT43), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n496), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n578), .A2(new_n620), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n728), .B1(new_n735), .B2(KEYINPUT44), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n578), .A2(KEYINPUT44), .A3(new_n620), .A4(new_n734), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n731), .A2(new_n733), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n574), .B2(new_n577), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(KEYINPUT108), .A3(KEYINPUT44), .A4(new_n620), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n727), .A2(new_n737), .A3(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT110), .B(G137), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G39));
  NAND2_X1  g562(.A1(new_n725), .A2(new_n581), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n500), .B1(new_n722), .B2(new_n724), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT47), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n694), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n696), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n307), .A2(new_n348), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT111), .B(G140), .Z(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G42));
  XOR2_X1   g573(.A(new_n664), .B(KEYINPUT49), .Z(new_n760));
  INV_X1    g574(.A(new_n650), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n641), .A2(new_n347), .A3(new_n500), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n730), .A2(new_n606), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n760), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT112), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n663), .A2(new_n500), .A3(new_n567), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n751), .A2(new_n753), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n348), .A2(new_n453), .A3(new_n677), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n741), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n728), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n665), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n606), .B1(new_n639), .B2(new_n640), .ZN(new_n772));
  NOR4_X1   g586(.A1(new_n768), .A2(new_n771), .A3(new_n772), .A4(new_n741), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT50), .B1(new_n773), .B2(KEYINPUT114), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT114), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n769), .A2(new_n665), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n775), .B(new_n776), .C1(new_n777), .C2(new_n772), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n696), .A2(new_n663), .A3(new_n581), .A4(new_n567), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n626), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n665), .A2(KEYINPUT115), .A3(new_n696), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n682), .A4(new_n734), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT116), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n497), .A2(new_n729), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n348), .A3(new_n761), .A4(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n770), .A2(new_n779), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n791), .A2(new_n792), .A3(new_n452), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n769), .A2(new_n607), .A3(new_n665), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n589), .B1(new_n496), .B2(new_n447), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n679), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n569), .B(new_n621), .C1(new_n582), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n706), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n666), .A2(new_n669), .A3(new_n672), .A4(new_n680), .ZN(new_n801));
  INV_X1    g615(.A(new_n703), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n601), .A2(new_n629), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n307), .A2(new_n568), .A3(new_n446), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n695), .A2(new_n677), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(new_n620), .A3(new_n696), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n800), .A2(new_n801), .A3(new_n802), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n642), .A2(new_n416), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n620), .A2(new_n628), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n650), .A2(new_n699), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n632), .A2(new_n660), .A3(new_n811), .A4(new_n683), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT52), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n795), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n812), .B(new_n815), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n651), .B(new_n755), .C1(new_n804), .C2(new_n805), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n817), .A2(new_n799), .A3(new_n706), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n669), .A2(new_n672), .A3(new_n680), .A4(new_n666), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n703), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n816), .A2(KEYINPUT53), .A3(new_n818), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n814), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT54), .ZN(new_n823));
  XOR2_X1   g637(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n814), .A2(new_n821), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n793), .A2(new_n794), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n348), .A2(new_n786), .A3(new_n589), .A4(new_n761), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n786), .A2(new_n687), .A3(new_n734), .ZN(new_n829));
  XOR2_X1   g643(.A(new_n829), .B(KEYINPUT48), .Z(new_n830));
  NOR3_X1   g644(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(G952), .A2(G953), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n765), .B1(new_n831), .B2(new_n832), .ZN(G75));
  OAI21_X1  g647(.A(new_n388), .B1(new_n392), .B2(new_n393), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(new_n353), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT55), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n836), .B1(KEYINPUT117), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n308), .B1(new_n814), .B2(new_n821), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(G210), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n839), .B1(new_n841), .B2(new_n837), .ZN(new_n842));
  AOI211_X1 g656(.A(KEYINPUT56), .B(new_n838), .C1(new_n840), .C2(G210), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n242), .A2(G952), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(G51));
  XOR2_X1   g659(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n846));
  NAND2_X1  g660(.A1(new_n714), .A2(new_n846), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n714), .A2(new_n846), .ZN(new_n848));
  INV_X1    g662(.A(new_n826), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n825), .B1(new_n814), .B2(new_n821), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n565), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n840), .A2(new_n709), .A3(new_n710), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n844), .B1(new_n852), .B2(new_n853), .ZN(G54));
  NAND3_X1  g668(.A1(new_n840), .A2(KEYINPUT58), .A3(G475), .ZN(new_n855));
  INV_X1    g669(.A(new_n483), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n857), .A2(new_n858), .A3(new_n844), .ZN(G60));
  AND2_X1   g673(.A1(new_n584), .A2(new_n585), .ZN(new_n860));
  NAND2_X1  g674(.A1(G478), .A2(G902), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(KEYINPUT59), .Z(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n860), .B(new_n863), .C1(new_n849), .C2(new_n850), .ZN(new_n864));
  INV_X1    g678(.A(new_n844), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n862), .B1(new_n823), .B2(new_n826), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(new_n860), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(G63));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n869));
  NAND2_X1  g683(.A1(G217), .A2(G902), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT60), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n344), .B1(new_n822), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n869), .B1(new_n873), .B2(new_n844), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n871), .B1(new_n814), .B2(new_n821), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n618), .ZN(new_n876));
  OAI211_X1 g690(.A(KEYINPUT120), .B(new_n865), .C1(new_n875), .C2(new_n344), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g692(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n873), .A2(new_n844), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(KEYINPUT61), .A3(new_n876), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n882), .ZN(G66));
  NOR2_X1   g697(.A1(new_n819), .A2(new_n799), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n242), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT121), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n242), .B1(new_n454), .B2(G224), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n888), .B(KEYINPUT122), .Z(new_n889));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n834), .B1(G898), .B2(new_n242), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n890), .B(new_n891), .ZN(G69));
  AOI211_X1 g706(.A(new_n736), .B(new_n744), .C1(new_n719), .C2(new_n726), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n754), .B2(new_n756), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n307), .A2(new_n348), .A3(new_n696), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n895), .A2(new_n636), .A3(new_n796), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT123), .Z(new_n897));
  NAND3_X1  g711(.A1(new_n632), .A2(new_n660), .A3(new_n683), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n653), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(KEYINPUT62), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n653), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n894), .B(new_n897), .C1(new_n900), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n242), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n267), .B(new_n480), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n242), .A2(G900), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT125), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n893), .B2(new_n898), .ZN(new_n910));
  INV_X1    g724(.A(new_n898), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n746), .A2(KEYINPUT126), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n703), .B1(new_n754), .B2(new_n756), .ZN(new_n914));
  INV_X1    g728(.A(new_n726), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT107), .B1(new_n752), .B2(new_n635), .ZN(new_n916));
  OAI211_X1 g730(.A(new_n687), .B(new_n809), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n727), .A2(KEYINPUT127), .A3(new_n687), .A4(new_n809), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n706), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n913), .A2(new_n914), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n908), .B1(new_n922), .B2(new_n242), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n906), .B1(new_n923), .B2(new_n905), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT124), .B1(new_n923), .B2(new_n905), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n242), .B1(G227), .B2(G900), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  OAI221_X1 g742(.A(new_n906), .B1(KEYINPUT124), .B2(new_n926), .C1(new_n923), .C2(new_n905), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(G72));
  NAND2_X1  g744(.A1(G472), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT63), .Z(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n903), .B2(new_n885), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n647), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n822), .B(new_n932), .C1(new_n299), .C2(new_n674), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n865), .A3(new_n935), .ZN(new_n936));
  OR2_X1    g750(.A1(new_n922), .A2(new_n885), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n297), .B1(new_n937), .B2(new_n932), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n936), .B1(new_n248), .B2(new_n938), .ZN(G57));
endmodule


