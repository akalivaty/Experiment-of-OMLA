

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768;

  AND2_X1 U373 ( .A1(n768), .A2(n645), .ZN(n552) );
  NOR2_X1 U374 ( .A1(n681), .A2(n679), .ZN(n596) );
  XNOR2_X1 U375 ( .A(n586), .B(n587), .ZN(n676) );
  NOR2_X2 U376 ( .A1(G953), .A2(G237), .ZN(n376) );
  NAND2_X2 U377 ( .A1(n399), .A2(n414), .ZN(n608) );
  NOR2_X2 U378 ( .A1(n589), .A2(n582), .ZN(n583) );
  NOR2_X2 U379 ( .A1(n765), .A2(n767), .ZN(n598) );
  NOR2_X2 U380 ( .A1(n558), .A2(n607), .ZN(n486) );
  INV_X2 U381 ( .A(n562), .ZN(n594) );
  XNOR2_X1 U382 ( .A(n452), .B(n451), .ZN(n488) );
  XNOR2_X1 U383 ( .A(G113), .B(G119), .ZN(n440) );
  NOR2_X1 U384 ( .A1(n552), .A2(KEYINPUT44), .ZN(n424) );
  XNOR2_X1 U385 ( .A(n548), .B(KEYINPUT32), .ZN(n768) );
  XNOR2_X1 U386 ( .A(n397), .B(n364), .ZN(n544) );
  OR2_X1 U387 ( .A1(n734), .A2(G902), .ZN(n397) );
  AND2_X1 U388 ( .A1(n422), .A2(KEYINPUT87), .ZN(n415) );
  XNOR2_X1 U389 ( .A(n488), .B(n487), .ZN(n744) );
  XNOR2_X1 U390 ( .A(n388), .B(n453), .ZN(n387) );
  XNOR2_X1 U391 ( .A(n440), .B(KEYINPUT72), .ZN(n452) );
  INV_X2 U392 ( .A(G953), .ZN(n758) );
  NOR2_X1 U393 ( .A1(n561), .A2(n540), .ZN(n350) );
  BUF_X1 U394 ( .A(n768), .Z(n351) );
  XNOR2_X1 U395 ( .A(n352), .B(KEYINPUT34), .ZN(n534) );
  NOR2_X1 U396 ( .A1(n372), .A2(n708), .ZN(n352) );
  NAND2_X1 U397 ( .A1(n688), .A2(n687), .ZN(n558) );
  BUF_X1 U398 ( .A(n380), .Z(n353) );
  NAND2_X1 U399 ( .A1(KEYINPUT24), .A2(n355), .ZN(n356) );
  NAND2_X1 U400 ( .A1(n354), .A2(G110), .ZN(n357) );
  NAND2_X1 U401 ( .A1(n356), .A2(n357), .ZN(n472) );
  INV_X1 U402 ( .A(KEYINPUT24), .ZN(n354) );
  INV_X1 U403 ( .A(G110), .ZN(n355) );
  XNOR2_X1 U404 ( .A(n350), .B(n369), .ZN(n358) );
  BUF_X1 U405 ( .A(n632), .Z(n359) );
  XNOR2_X1 U406 ( .A(n541), .B(n369), .ZN(n554) );
  XNOR2_X1 U407 ( .A(n375), .B(n377), .ZN(n632) );
  XNOR2_X2 U408 ( .A(n360), .B(n361), .ZN(n562) );
  NOR2_X1 U409 ( .A1(n722), .A2(G902), .ZN(n360) );
  XOR2_X1 U410 ( .A(KEYINPUT71), .B(G469), .Z(n361) );
  NAND2_X1 U411 ( .A1(n418), .A2(KEYINPUT87), .ZN(n417) );
  AND2_X1 U412 ( .A1(n386), .A2(n420), .ZN(n398) );
  INV_X1 U413 ( .A(n714), .ZN(n410) );
  INV_X1 U414 ( .A(KEYINPUT39), .ZN(n434) );
  NAND2_X1 U415 ( .A1(n413), .A2(n420), .ZN(n412) );
  INV_X1 U416 ( .A(n445), .ZN(n413) );
  NAND2_X1 U417 ( .A1(n629), .A2(KEYINPUT65), .ZN(n409) );
  INV_X1 U418 ( .A(G237), .ZN(n497) );
  XNOR2_X1 U419 ( .A(n385), .B(KEYINPUT45), .ZN(n630) );
  XNOR2_X1 U420 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n449) );
  XNOR2_X1 U421 ( .A(G137), .B(KEYINPUT69), .ZN(n476) );
  XOR2_X1 U422 ( .A(KEYINPUT79), .B(KEYINPUT74), .Z(n473) );
  XNOR2_X1 U423 ( .A(n493), .B(n470), .ZN(n754) );
  XNOR2_X1 U424 ( .A(G140), .B(KEYINPUT10), .ZN(n470) );
  XNOR2_X1 U425 ( .A(n443), .B(n442), .ZN(n527) );
  INV_X1 U426 ( .A(KEYINPUT8), .ZN(n442) );
  NAND2_X1 U427 ( .A1(n758), .A2(G234), .ZN(n443) );
  XNOR2_X1 U428 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n489) );
  XNOR2_X1 U429 ( .A(n469), .B(G125), .ZN(n493) );
  INV_X1 U430 ( .A(G146), .ZN(n469) );
  INV_X1 U431 ( .A(KEYINPUT83), .ZN(n379) );
  INV_X1 U432 ( .A(KEYINPUT1), .ZN(n400) );
  XNOR2_X1 U433 ( .A(n437), .B(n436), .ZN(n584) );
  INV_X1 U434 ( .A(KEYINPUT30), .ZN(n436) );
  AND2_X1 U435 ( .A1(n366), .A2(n390), .ZN(n593) );
  INV_X1 U436 ( .A(KEYINPUT87), .ZN(n421) );
  XOR2_X1 U437 ( .A(G131), .B(G134), .Z(n464) );
  INV_X1 U438 ( .A(n409), .ZN(n392) );
  NAND2_X1 U439 ( .A1(n446), .A2(n496), .ZN(n445) );
  NAND2_X1 U440 ( .A1(n499), .A2(n628), .ZN(n447) );
  XNOR2_X1 U441 ( .A(G113), .B(G131), .ZN(n509) );
  NAND2_X1 U442 ( .A1(G234), .A2(G237), .ZN(n501) );
  XNOR2_X1 U443 ( .A(G116), .B(G134), .ZN(n521) );
  AND2_X1 U444 ( .A1(n737), .A2(n367), .ZN(n714) );
  XNOR2_X1 U445 ( .A(n381), .B(KEYINPUT107), .ZN(n619) );
  INV_X1 U446 ( .A(KEYINPUT19), .ZN(n401) );
  INV_X1 U447 ( .A(n591), .ZN(n389) );
  INV_X1 U448 ( .A(KEYINPUT105), .ZN(n391) );
  INV_X1 U449 ( .A(n760), .ZN(n393) );
  XNOR2_X1 U450 ( .A(n477), .B(n448), .ZN(n478) );
  XOR2_X1 U451 ( .A(n638), .B(KEYINPUT59), .Z(n639) );
  XNOR2_X1 U452 ( .A(n744), .B(n495), .ZN(n377) );
  XNOR2_X1 U453 ( .A(n433), .B(n588), .ZN(n765) );
  NAND2_X1 U454 ( .A1(n557), .A2(n556), .ZN(n427) );
  AND2_X1 U455 ( .A1(n402), .A2(n374), .ZN(n362) );
  AND2_X1 U456 ( .A1(n432), .A2(n447), .ZN(n363) );
  XOR2_X1 U457 ( .A(n482), .B(KEYINPUT25), .Z(n364) );
  OR2_X1 U458 ( .A1(n506), .A2(n581), .ZN(n365) );
  INV_X1 U459 ( .A(n496), .ZN(n628) );
  XNOR2_X1 U460 ( .A(G902), .B(KEYINPUT15), .ZN(n496) );
  AND2_X1 U461 ( .A1(n592), .A2(n591), .ZN(n366) );
  INV_X1 U462 ( .A(n675), .ZN(n418) );
  AND2_X1 U463 ( .A1(n378), .A2(KEYINPUT2), .ZN(n367) );
  AND2_X1 U464 ( .A1(n674), .A2(n644), .ZN(n368) );
  AND2_X1 U465 ( .A1(n675), .A2(n421), .ZN(n420) );
  XOR2_X1 U466 ( .A(KEYINPUT75), .B(KEYINPUT22), .Z(n369) );
  OR2_X1 U467 ( .A1(n629), .A2(KEYINPUT65), .ZN(n370) );
  XOR2_X1 U468 ( .A(KEYINPUT84), .B(KEYINPUT48), .Z(n371) );
  XNOR2_X1 U469 ( .A(n508), .B(KEYINPUT0), .ZN(n372) );
  XNOR2_X1 U470 ( .A(n508), .B(KEYINPUT0), .ZN(n561) );
  XNOR2_X1 U471 ( .A(n694), .B(n391), .ZN(n390) );
  BUF_X1 U472 ( .A(n694), .Z(n384) );
  XNOR2_X1 U473 ( .A(n486), .B(n485), .ZN(n708) );
  NAND2_X1 U474 ( .A1(n407), .A2(n370), .ZN(n406) );
  BUF_X1 U475 ( .A(n608), .Z(n373) );
  XNOR2_X1 U476 ( .A(n373), .B(n401), .ZN(n374) );
  XNOR2_X1 U477 ( .A(n608), .B(n401), .ZN(n507) );
  INV_X1 U478 ( .A(n603), .ZN(n402) );
  NAND2_X1 U479 ( .A1(n419), .A2(n417), .ZN(n416) );
  OR2_X1 U480 ( .A1(n632), .A2(n412), .ZN(n419) );
  BUF_X1 U481 ( .A(n721), .Z(n732) );
  NAND2_X1 U482 ( .A1(n432), .A2(n447), .ZN(n386) );
  XOR2_X1 U483 ( .A(KEYINPUT62), .B(n648), .Z(n649) );
  NAND2_X1 U484 ( .A1(n394), .A2(n368), .ZN(n380) );
  OR2_X1 U485 ( .A1(n618), .A2(n670), .ZN(n674) );
  XNOR2_X1 U486 ( .A(n462), .B(n746), .ZN(n375) );
  XNOR2_X1 U487 ( .A(n462), .B(n746), .ZN(n383) );
  INV_X1 U488 ( .A(n737), .ZN(n711) );
  BUF_X1 U489 ( .A(n630), .Z(n737) );
  NAND2_X1 U490 ( .A1(n376), .A2(G210), .ZN(n388) );
  NAND2_X1 U491 ( .A1(n376), .A2(G214), .ZN(n512) );
  XNOR2_X2 U492 ( .A(n757), .B(G101), .ZN(n462) );
  XNOR2_X2 U493 ( .A(n530), .B(n449), .ZN(n757) );
  INV_X1 U494 ( .A(n353), .ZN(n378) );
  XNOR2_X2 U495 ( .A(n380), .B(n379), .ZN(n712) );
  INV_X1 U496 ( .A(n542), .ZN(n607) );
  NAND2_X1 U497 ( .A1(n382), .A2(n542), .ZN(n381) );
  AND2_X1 U498 ( .A1(n664), .A2(n366), .ZN(n382) );
  XNOR2_X1 U499 ( .A(n383), .B(n468), .ZN(n722) );
  NOR2_X2 U500 ( .A1(n627), .A2(n409), .ZN(n408) );
  XNOR2_X2 U501 ( .A(n576), .B(n575), .ZN(n627) );
  NAND2_X1 U502 ( .A1(n429), .A2(n425), .ZN(n385) );
  NAND2_X1 U503 ( .A1(n428), .A2(n427), .ZN(n426) );
  NOR2_X1 U504 ( .A1(n408), .A2(n406), .ZN(n405) );
  NOR2_X1 U505 ( .A1(n574), .A2(n426), .ZN(n425) );
  AND2_X2 U506 ( .A1(n411), .A2(n410), .ZN(n721) );
  NOR2_X1 U507 ( .A1(n712), .A2(KEYINPUT65), .ZN(n404) );
  XNOR2_X1 U508 ( .A(n387), .B(n464), .ZN(n457) );
  NOR2_X1 U509 ( .A1(n390), .A2(n389), .ZN(n549) );
  NAND2_X1 U510 ( .A1(n390), .A2(n675), .ZN(n437) );
  NAND2_X1 U511 ( .A1(n712), .A2(n392), .ZN(n407) );
  XNOR2_X1 U512 ( .A(n712), .B(n393), .ZN(n759) );
  XNOR2_X1 U513 ( .A(n395), .B(n371), .ZN(n394) );
  NAND2_X1 U514 ( .A1(n617), .A2(n616), .ZN(n395) );
  XNOR2_X2 U515 ( .A(n396), .B(KEYINPUT67), .ZN(n687) );
  NAND2_X1 U516 ( .A1(n544), .A2(n441), .ZN(n396) );
  NOR2_X1 U517 ( .A1(n398), .A2(n416), .ZN(n399) );
  INV_X1 U518 ( .A(n688), .ZN(n621) );
  XNOR2_X2 U519 ( .A(n562), .B(n400), .ZN(n688) );
  NAND2_X1 U520 ( .A1(n405), .A2(n403), .ZN(n411) );
  NAND2_X1 U521 ( .A1(n627), .A2(n404), .ZN(n403) );
  OR2_X1 U522 ( .A1(n632), .A2(n445), .ZN(n422) );
  XNOR2_X1 U523 ( .A(n479), .B(n478), .ZN(n734) );
  XNOR2_X1 U524 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U525 ( .A1(n599), .A2(n676), .ZN(n435) );
  NAND2_X1 U526 ( .A1(n363), .A2(n422), .ZN(n586) );
  NAND2_X1 U527 ( .A1(n415), .A2(n363), .ZN(n414) );
  NAND2_X1 U528 ( .A1(n423), .A2(n552), .ZN(n430) );
  NAND2_X1 U529 ( .A1(n573), .A2(n551), .ZN(n423) );
  NAND2_X1 U530 ( .A1(n424), .A2(n538), .ZN(n431) );
  INV_X1 U531 ( .A(n571), .ZN(n428) );
  INV_X1 U532 ( .A(n427), .ZN(n654) );
  NAND2_X1 U533 ( .A1(n431), .A2(n430), .ZN(n429) );
  NAND2_X1 U534 ( .A1(n632), .A2(n499), .ZN(n432) );
  NOR2_X2 U535 ( .A1(n618), .A2(n667), .ZN(n433) );
  XNOR2_X2 U536 ( .A(n435), .B(n434), .ZN(n618) );
  XNOR2_X2 U537 ( .A(n438), .B(G472), .ZN(n694) );
  NAND2_X1 U538 ( .A1(n648), .A2(n498), .ZN(n438) );
  XNOR2_X1 U539 ( .A(n462), .B(n439), .ZN(n648) );
  XNOR2_X1 U540 ( .A(n458), .B(n488), .ZN(n439) );
  INV_X1 U541 ( .A(n544), .ZN(n591) );
  NAND2_X1 U542 ( .A1(n594), .A2(n687), .ZN(n582) );
  INV_X1 U543 ( .A(n691), .ZN(n441) );
  XNOR2_X2 U544 ( .A(n444), .B(G143), .ZN(n530) );
  XNOR2_X2 U545 ( .A(G128), .B(KEYINPUT64), .ZN(n444) );
  INV_X1 U546 ( .A(n499), .ZN(n446) );
  NOR2_X2 U547 ( .A1(n641), .A2(n736), .ZN(n643) );
  XOR2_X1 U548 ( .A(n476), .B(KEYINPUT23), .Z(n448) );
  INV_X1 U549 ( .A(KEYINPUT82), .ZN(n575) );
  INV_X1 U550 ( .A(KEYINPUT77), .ZN(n453) );
  NAND2_X1 U551 ( .A1(n507), .A2(n365), .ZN(n508) );
  XNOR2_X1 U552 ( .A(KEYINPUT60), .B(KEYINPUT66), .ZN(n642) );
  XNOR2_X1 U553 ( .A(G116), .B(KEYINPUT73), .ZN(n450) );
  XNOR2_X1 U554 ( .A(n450), .B(KEYINPUT3), .ZN(n451) );
  XOR2_X1 U555 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n455) );
  XNOR2_X1 U556 ( .A(G146), .B(G137), .ZN(n454) );
  XNOR2_X1 U557 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U558 ( .A(n457), .B(n456), .ZN(n458) );
  INV_X1 U559 ( .A(G902), .ZN(n498) );
  XOR2_X1 U560 ( .A(KEYINPUT102), .B(KEYINPUT6), .Z(n459) );
  XNOR2_X1 U561 ( .A(n694), .B(n459), .ZN(n542) );
  XNOR2_X1 U562 ( .A(G110), .B(G107), .ZN(n461) );
  INV_X1 U563 ( .A(G104), .ZN(n460) );
  XNOR2_X1 U564 ( .A(n461), .B(n460), .ZN(n746) );
  INV_X1 U565 ( .A(n476), .ZN(n463) );
  XOR2_X1 U566 ( .A(n464), .B(n463), .Z(n753) );
  XOR2_X1 U567 ( .A(G146), .B(G140), .Z(n466) );
  NAND2_X1 U568 ( .A1(G227), .A2(n758), .ZN(n465) );
  XOR2_X1 U569 ( .A(n466), .B(n465), .Z(n467) );
  XNOR2_X1 U570 ( .A(n753), .B(n467), .ZN(n468) );
  XNOR2_X1 U571 ( .A(G128), .B(G119), .ZN(n471) );
  XNOR2_X1 U572 ( .A(n472), .B(n471), .ZN(n474) );
  XNOR2_X1 U573 ( .A(n475), .B(n754), .ZN(n479) );
  NAND2_X1 U574 ( .A1(G221), .A2(n527), .ZN(n477) );
  XOR2_X1 U575 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n481) );
  NAND2_X1 U576 ( .A1(G234), .A2(n496), .ZN(n480) );
  XNOR2_X1 U577 ( .A(n481), .B(n480), .ZN(n483) );
  NAND2_X1 U578 ( .A1(G217), .A2(n483), .ZN(n482) );
  NAND2_X1 U579 ( .A1(n483), .A2(G221), .ZN(n484) );
  XNOR2_X1 U580 ( .A(KEYINPUT21), .B(n484), .ZN(n691) );
  XNOR2_X1 U581 ( .A(KEYINPUT88), .B(KEYINPUT33), .ZN(n485) );
  XNOR2_X1 U582 ( .A(KEYINPUT16), .B(G122), .ZN(n487) );
  XOR2_X1 U583 ( .A(KEYINPUT91), .B(KEYINPUT89), .Z(n490) );
  XNOR2_X1 U584 ( .A(n490), .B(n489), .ZN(n492) );
  NAND2_X1 U585 ( .A1(n758), .A2(G224), .ZN(n491) );
  XNOR2_X1 U586 ( .A(n492), .B(n491), .ZN(n494) );
  XNOR2_X1 U587 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U588 ( .A1(n498), .A2(n497), .ZN(n500) );
  AND2_X1 U589 ( .A1(n500), .A2(G210), .ZN(n499) );
  NAND2_X1 U590 ( .A1(n500), .A2(G214), .ZN(n675) );
  XNOR2_X1 U591 ( .A(n501), .B(KEYINPUT92), .ZN(n502) );
  XNOR2_X1 U592 ( .A(KEYINPUT14), .B(n502), .ZN(n505) );
  NAND2_X1 U593 ( .A1(G902), .A2(n505), .ZN(n577) );
  NOR2_X1 U594 ( .A1(G898), .A2(n758), .ZN(n503) );
  XNOR2_X1 U595 ( .A(KEYINPUT93), .B(n503), .ZN(n747) );
  NOR2_X1 U596 ( .A1(n577), .A2(n747), .ZN(n504) );
  XNOR2_X1 U597 ( .A(n504), .B(KEYINPUT94), .ZN(n506) );
  NAND2_X1 U598 ( .A1(G952), .A2(n505), .ZN(n706) );
  NOR2_X1 U599 ( .A1(n706), .A2(G953), .ZN(n581) );
  XNOR2_X1 U600 ( .A(KEYINPUT13), .B(G475), .ZN(n520) );
  XOR2_X1 U601 ( .A(KEYINPUT98), .B(G122), .Z(n510) );
  XNOR2_X1 U602 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U603 ( .A(n754), .B(n511), .ZN(n518) );
  XOR2_X1 U604 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n513) );
  XNOR2_X1 U605 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U606 ( .A(n514), .B(KEYINPUT11), .Z(n516) );
  XNOR2_X1 U607 ( .A(G143), .B(G104), .ZN(n515) );
  XNOR2_X1 U608 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U609 ( .A(n518), .B(n517), .ZN(n638) );
  NOR2_X1 U610 ( .A1(G902), .A2(n638), .ZN(n519) );
  XOR2_X1 U611 ( .A(n520), .B(n519), .Z(n566) );
  INV_X1 U612 ( .A(n566), .ZN(n567) );
  XOR2_X1 U613 ( .A(G107), .B(G122), .Z(n522) );
  XNOR2_X1 U614 ( .A(n522), .B(n521), .ZN(n526) );
  XOR2_X1 U615 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n524) );
  XNOR2_X1 U616 ( .A(KEYINPUT7), .B(KEYINPUT100), .ZN(n523) );
  XNOR2_X1 U617 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U618 ( .A(n526), .B(n525), .Z(n529) );
  NAND2_X1 U619 ( .A1(G217), .A2(n527), .ZN(n528) );
  XNOR2_X1 U620 ( .A(n529), .B(n528), .ZN(n531) );
  XNOR2_X1 U621 ( .A(n530), .B(n531), .ZN(n728) );
  NOR2_X1 U622 ( .A1(G902), .A2(n728), .ZN(n532) );
  XNOR2_X1 U623 ( .A(G478), .B(n532), .ZN(n568) );
  INV_X1 U624 ( .A(n568), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n567), .A2(n565), .ZN(n600) );
  INV_X1 U626 ( .A(n600), .ZN(n533) );
  NAND2_X1 U627 ( .A1(n534), .A2(n533), .ZN(n536) );
  INV_X1 U628 ( .A(KEYINPUT35), .ZN(n535) );
  XNOR2_X2 U629 ( .A(n536), .B(n535), .ZN(n573) );
  INV_X1 U630 ( .A(KEYINPUT86), .ZN(n537) );
  NAND2_X1 U631 ( .A1(n573), .A2(n537), .ZN(n538) );
  NAND2_X1 U632 ( .A1(n566), .A2(n568), .ZN(n679) );
  NOR2_X1 U633 ( .A1(n679), .A2(n691), .ZN(n539) );
  XNOR2_X1 U634 ( .A(n539), .B(KEYINPUT103), .ZN(n540) );
  NOR2_X2 U635 ( .A1(n561), .A2(n540), .ZN(n541) );
  XNOR2_X1 U636 ( .A(KEYINPUT80), .B(n542), .ZN(n545) );
  INV_X1 U637 ( .A(KEYINPUT104), .ZN(n543) );
  XNOR2_X1 U638 ( .A(n389), .B(n543), .ZN(n690) );
  INV_X1 U639 ( .A(n690), .ZN(n556) );
  NOR2_X1 U640 ( .A1(n545), .A2(n556), .ZN(n546) );
  AND2_X1 U641 ( .A1(n688), .A2(n546), .ZN(n547) );
  NAND2_X1 U642 ( .A1(n554), .A2(n547), .ZN(n548) );
  AND2_X1 U643 ( .A1(n549), .A2(n621), .ZN(n550) );
  NAND2_X1 U644 ( .A1(n358), .A2(n550), .ZN(n645) );
  INV_X1 U645 ( .A(KEYINPUT44), .ZN(n572) );
  AND2_X1 U646 ( .A1(n572), .A2(KEYINPUT86), .ZN(n551) );
  AND2_X1 U647 ( .A1(n607), .A2(n621), .ZN(n553) );
  NAND2_X1 U648 ( .A1(n358), .A2(n553), .ZN(n555) );
  XNOR2_X1 U649 ( .A(n555), .B(KEYINPUT85), .ZN(n557) );
  INV_X1 U650 ( .A(n558), .ZN(n559) );
  NAND2_X1 U651 ( .A1(n384), .A2(n559), .ZN(n697) );
  NOR2_X1 U652 ( .A1(n372), .A2(n697), .ZN(n560) );
  XNOR2_X1 U653 ( .A(n560), .B(KEYINPUT31), .ZN(n669) );
  INV_X1 U654 ( .A(n372), .ZN(n564) );
  NOR2_X1 U655 ( .A1(n582), .A2(n384), .ZN(n563) );
  NAND2_X1 U656 ( .A1(n564), .A2(n563), .ZN(n656) );
  NAND2_X1 U657 ( .A1(n669), .A2(n656), .ZN(n569) );
  NOR2_X1 U658 ( .A1(n566), .A2(n565), .ZN(n664) );
  NOR2_X1 U659 ( .A1(n568), .A2(n567), .ZN(n660) );
  NOR2_X1 U660 ( .A1(n664), .A2(n660), .ZN(n682) );
  INV_X1 U661 ( .A(n682), .ZN(n604) );
  NAND2_X1 U662 ( .A1(n569), .A2(n604), .ZN(n570) );
  XNOR2_X1 U663 ( .A(n570), .B(KEYINPUT101), .ZN(n571) );
  NOR2_X1 U664 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U665 ( .A1(n630), .A2(n628), .ZN(n576) );
  NOR2_X1 U666 ( .A1(G900), .A2(n577), .ZN(n578) );
  NAND2_X1 U667 ( .A1(G953), .A2(n578), .ZN(n579) );
  XOR2_X1 U668 ( .A(KEYINPUT106), .B(n579), .Z(n580) );
  NOR2_X1 U669 ( .A1(n581), .A2(n580), .ZN(n589) );
  XNOR2_X1 U670 ( .A(n583), .B(KEYINPUT78), .ZN(n585) );
  AND2_X2 U671 ( .A1(n585), .A2(n584), .ZN(n599) );
  XOR2_X1 U672 ( .A(KEYINPUT76), .B(KEYINPUT38), .Z(n587) );
  INV_X1 U673 ( .A(n664), .ZN(n667) );
  XNOR2_X1 U674 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n588) );
  NOR2_X1 U675 ( .A1(n691), .A2(n589), .ZN(n590) );
  XNOR2_X1 U676 ( .A(KEYINPUT70), .B(n590), .ZN(n592) );
  XNOR2_X1 U677 ( .A(KEYINPUT28), .B(n593), .ZN(n595) );
  NAND2_X1 U678 ( .A1(n595), .A2(n594), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n676), .A2(n675), .ZN(n681) );
  XNOR2_X1 U680 ( .A(n596), .B(KEYINPUT41), .ZN(n707) );
  NOR2_X1 U681 ( .A1(n603), .A2(n707), .ZN(n597) );
  XNOR2_X1 U682 ( .A(n597), .B(KEYINPUT42), .ZN(n767) );
  XNOR2_X1 U683 ( .A(n598), .B(KEYINPUT46), .ZN(n617) );
  INV_X1 U684 ( .A(n599), .ZN(n601) );
  NOR2_X1 U685 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U686 ( .A1(n602), .A2(n586), .ZN(n647) );
  NAND2_X1 U687 ( .A1(n362), .A2(n604), .ZN(n613) );
  NAND2_X1 U688 ( .A1(n613), .A2(KEYINPUT47), .ZN(n605) );
  NAND2_X1 U689 ( .A1(n647), .A2(n605), .ZN(n606) );
  XNOR2_X1 U690 ( .A(n606), .B(KEYINPUT81), .ZN(n612) );
  NAND2_X1 U691 ( .A1(n619), .A2(n373), .ZN(n610) );
  XNOR2_X1 U692 ( .A(KEYINPUT36), .B(KEYINPUT111), .ZN(n609) );
  XNOR2_X1 U693 ( .A(n610), .B(n609), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n611), .A2(n688), .ZN(n673) );
  NAND2_X1 U695 ( .A1(n612), .A2(n673), .ZN(n615) );
  NOR2_X1 U696 ( .A1(KEYINPUT47), .A2(n613), .ZN(n614) );
  NOR2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n616) );
  INV_X1 U698 ( .A(n660), .ZN(n670) );
  XOR2_X1 U699 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n624) );
  NAND2_X1 U700 ( .A1(n619), .A2(n675), .ZN(n620) );
  XOR2_X1 U701 ( .A(KEYINPUT108), .B(n620), .Z(n622) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n624), .B(n623), .ZN(n626) );
  INV_X1 U704 ( .A(n586), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n644) );
  NAND2_X1 U706 ( .A1(n628), .A2(KEYINPUT2), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n721), .A2(G210), .ZN(n634) );
  XOR2_X1 U708 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n631) );
  XNOR2_X1 U709 ( .A(n359), .B(n631), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n634), .B(n633), .ZN(n636) );
  INV_X1 U711 ( .A(G952), .ZN(n635) );
  AND2_X1 U712 ( .A1(n635), .A2(G953), .ZN(n736) );
  NOR2_X2 U713 ( .A1(n636), .A2(n736), .ZN(n637) );
  XNOR2_X1 U714 ( .A(n637), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U715 ( .A1(n721), .A2(G475), .ZN(n640) );
  XNOR2_X1 U716 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U717 ( .A(n643), .B(n642), .ZN(G60) );
  XNOR2_X1 U718 ( .A(n644), .B(G140), .ZN(G42) );
  XNOR2_X1 U719 ( .A(n645), .B(G110), .ZN(G12) );
  XOR2_X1 U720 ( .A(G143), .B(KEYINPUT113), .Z(n646) );
  XNOR2_X1 U721 ( .A(n647), .B(n646), .ZN(G45) );
  NAND2_X1 U722 ( .A1(n721), .A2(G472), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n650), .B(n649), .ZN(n651) );
  NOR2_X2 U724 ( .A1(n651), .A2(n736), .ZN(n653) );
  XOR2_X1 U725 ( .A(KEYINPUT90), .B(KEYINPUT63), .Z(n652) );
  XNOR2_X1 U726 ( .A(n653), .B(n652), .ZN(G57) );
  XOR2_X1 U727 ( .A(G101), .B(n654), .Z(G3) );
  NOR2_X1 U728 ( .A1(n667), .A2(n656), .ZN(n655) );
  XOR2_X1 U729 ( .A(G104), .B(n655), .Z(G6) );
  NOR2_X1 U730 ( .A1(n670), .A2(n656), .ZN(n658) );
  XNOR2_X1 U731 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U733 ( .A(G107), .B(n659), .ZN(G9) );
  XOR2_X1 U734 ( .A(KEYINPUT29), .B(KEYINPUT112), .Z(n662) );
  NAND2_X1 U735 ( .A1(n362), .A2(n660), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U737 ( .A(G128), .B(n663), .ZN(G30) );
  NAND2_X1 U738 ( .A1(n362), .A2(n664), .ZN(n665) );
  XNOR2_X1 U739 ( .A(n665), .B(KEYINPUT114), .ZN(n666) );
  XNOR2_X1 U740 ( .A(G146), .B(n666), .ZN(G48) );
  NOR2_X1 U741 ( .A1(n667), .A2(n669), .ZN(n668) );
  XOR2_X1 U742 ( .A(G113), .B(n668), .Z(G15) );
  NOR2_X1 U743 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U744 ( .A(G116), .B(n671), .Z(G18) );
  XOR2_X1 U745 ( .A(G125), .B(KEYINPUT37), .Z(n672) );
  XNOR2_X1 U746 ( .A(n673), .B(n672), .ZN(G27) );
  XNOR2_X1 U747 ( .A(G134), .B(n674), .ZN(G36) );
  NOR2_X1 U748 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n677), .B(KEYINPUT116), .ZN(n678) );
  NOR2_X1 U750 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U751 ( .A(KEYINPUT117), .B(n680), .Z(n685) );
  NOR2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U753 ( .A(KEYINPUT118), .B(n683), .ZN(n684) );
  NOR2_X1 U754 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U755 ( .A1(n708), .A2(n686), .ZN(n703) );
  OR2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U757 ( .A(n689), .B(KEYINPUT50), .ZN(n696) );
  AND2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U759 ( .A(KEYINPUT49), .B(n692), .Z(n693) );
  NOR2_X1 U760 ( .A1(n384), .A2(n693), .ZN(n695) );
  NAND2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n698) );
  NAND2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n700) );
  XOR2_X1 U763 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n699) );
  XNOR2_X1 U764 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U765 ( .A1(n701), .A2(n707), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U767 ( .A(n704), .B(KEYINPUT52), .ZN(n705) );
  NOR2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n710) );
  NOR2_X1 U769 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U770 ( .A1(n710), .A2(n709), .ZN(n718) );
  NOR2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U772 ( .A1(n713), .A2(KEYINPUT2), .ZN(n715) );
  NOR2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U774 ( .A1(G953), .A2(n716), .ZN(n717) );
  NAND2_X1 U775 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U776 ( .A(KEYINPUT119), .B(n719), .ZN(n720) );
  XNOR2_X1 U777 ( .A(KEYINPUT53), .B(n720), .ZN(G75) );
  NAND2_X1 U778 ( .A1(n732), .A2(G469), .ZN(n726) );
  XOR2_X1 U779 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n724) );
  XNOR2_X1 U780 ( .A(n722), .B(KEYINPUT120), .ZN(n723) );
  XNOR2_X1 U781 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U782 ( .A(n726), .B(n725), .ZN(n727) );
  NOR2_X1 U783 ( .A1(n736), .A2(n727), .ZN(G54) );
  NAND2_X1 U784 ( .A1(n732), .A2(G478), .ZN(n730) );
  XOR2_X1 U785 ( .A(KEYINPUT121), .B(n728), .Z(n729) );
  XNOR2_X1 U786 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U787 ( .A1(n736), .A2(n731), .ZN(G63) );
  NAND2_X1 U788 ( .A1(n732), .A2(G217), .ZN(n733) );
  XNOR2_X1 U789 ( .A(n733), .B(n734), .ZN(n735) );
  NOR2_X1 U790 ( .A1(n736), .A2(n735), .ZN(G66) );
  NAND2_X1 U791 ( .A1(n737), .A2(n758), .ZN(n742) );
  NAND2_X1 U792 ( .A1(G224), .A2(G953), .ZN(n738) );
  XNOR2_X1 U793 ( .A(n738), .B(KEYINPUT122), .ZN(n739) );
  XNOR2_X1 U794 ( .A(KEYINPUT61), .B(n739), .ZN(n740) );
  NAND2_X1 U795 ( .A1(n740), .A2(G898), .ZN(n741) );
  NAND2_X1 U796 ( .A1(n742), .A2(n741), .ZN(n751) );
  XOR2_X1 U797 ( .A(G101), .B(KEYINPUT124), .Z(n743) );
  XNOR2_X1 U798 ( .A(n744), .B(n743), .ZN(n745) );
  XNOR2_X1 U799 ( .A(n746), .B(n745), .ZN(n748) );
  NAND2_X1 U800 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U801 ( .A(n749), .B(KEYINPUT125), .ZN(n750) );
  XNOR2_X1 U802 ( .A(n751), .B(n750), .ZN(n752) );
  XOR2_X1 U803 ( .A(KEYINPUT123), .B(n752), .Z(G69) );
  XOR2_X1 U804 ( .A(n754), .B(n753), .Z(n755) );
  XNOR2_X1 U805 ( .A(KEYINPUT126), .B(n755), .ZN(n756) );
  XNOR2_X1 U806 ( .A(n757), .B(n756), .ZN(n760) );
  NAND2_X1 U807 ( .A1(n759), .A2(n758), .ZN(n764) );
  XOR2_X1 U808 ( .A(G227), .B(n760), .Z(n761) );
  NAND2_X1 U809 ( .A1(n761), .A2(G900), .ZN(n762) );
  NAND2_X1 U810 ( .A1(n762), .A2(G953), .ZN(n763) );
  NAND2_X1 U811 ( .A1(n764), .A2(n763), .ZN(G72) );
  XOR2_X1 U812 ( .A(n765), .B(G131), .Z(G33) );
  XOR2_X1 U813 ( .A(n573), .B(G122), .Z(n766) );
  XNOR2_X1 U814 ( .A(n766), .B(KEYINPUT127), .ZN(G24) );
  XOR2_X1 U815 ( .A(n767), .B(G137), .Z(G39) );
  XNOR2_X1 U816 ( .A(n351), .B(G119), .ZN(G21) );
endmodule

