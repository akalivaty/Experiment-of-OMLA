

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U323 ( .A(n325), .B(n324), .ZN(n327) );
  XNOR2_X1 U324 ( .A(n410), .B(n323), .ZN(n324) );
  XNOR2_X1 U325 ( .A(n395), .B(n292), .ZN(n544) );
  XOR2_X1 U326 ( .A(n411), .B(n410), .Z(n517) );
  AND2_X1 U327 ( .A1(G232GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U328 ( .A(KEYINPUT111), .B(KEYINPUT48), .Z(n292) );
  XNOR2_X1 U329 ( .A(n334), .B(n291), .ZN(n335) );
  XOR2_X1 U330 ( .A(G43GAT), .B(G134GAT), .Z(n442) );
  INV_X1 U331 ( .A(KEYINPUT54), .ZN(n413) );
  XNOR2_X1 U332 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U333 ( .A(n342), .B(n371), .ZN(n343) );
  NOR2_X1 U334 ( .A1(n515), .A2(n415), .ZN(n567) );
  XNOR2_X1 U335 ( .A(n344), .B(n343), .ZN(n388) );
  XOR2_X1 U336 ( .A(n329), .B(n328), .Z(n574) );
  NOR2_X1 U337 ( .A1(n504), .A2(n513), .ZN(n510) );
  XNOR2_X1 U338 ( .A(KEYINPUT95), .B(n473), .ZN(n515) );
  XNOR2_X1 U339 ( .A(n453), .B(G190GAT), .ZN(n454) );
  XNOR2_X1 U340 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT1), .B(KEYINPUT93), .Z(n294) );
  XNOR2_X1 U342 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n293) );
  XNOR2_X1 U343 ( .A(n294), .B(n293), .ZN(n296) );
  XOR2_X1 U344 ( .A(G134GAT), .B(G148GAT), .Z(n295) );
  XNOR2_X1 U345 ( .A(n296), .B(n295), .ZN(n308) );
  XOR2_X1 U346 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n298) );
  XNOR2_X1 U347 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n300) );
  XNOR2_X1 U349 ( .A(G1GAT), .B(G127GAT), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n299), .B(G155GAT), .ZN(n321) );
  XOR2_X1 U351 ( .A(n300), .B(n321), .Z(n306) );
  XNOR2_X1 U352 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n301), .B(G120GAT), .ZN(n446) );
  XOR2_X1 U354 ( .A(KEYINPUT87), .B(G162GAT), .Z(n303) );
  XNOR2_X1 U355 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U357 ( .A(G141GAT), .B(n304), .Z(n430) );
  XNOR2_X1 U358 ( .A(n446), .B(n430), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n310) );
  NAND2_X1 U361 ( .A1(G225GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U363 ( .A(n311), .B(KEYINPUT94), .Z(n314) );
  XNOR2_X1 U364 ( .A(G29GAT), .B(KEYINPUT77), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n312), .B(G85GAT), .ZN(n338) );
  XNOR2_X1 U366 ( .A(n338), .B(KEYINPUT5), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n473) );
  XOR2_X1 U368 ( .A(KEYINPUT73), .B(KEYINPUT13), .Z(n316) );
  XNOR2_X1 U369 ( .A(G71GAT), .B(G78GAT), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U371 ( .A(G57GAT), .B(n317), .Z(n359) );
  XOR2_X1 U372 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n319) );
  XNOR2_X1 U373 ( .A(G64GAT), .B(KEYINPUT79), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n359), .B(n320), .ZN(n329) );
  XOR2_X1 U376 ( .A(G22GAT), .B(G15GAT), .Z(n367) );
  XOR2_X1 U377 ( .A(n321), .B(n367), .Z(n325) );
  XNOR2_X1 U378 ( .A(G8GAT), .B(G183GAT), .ZN(n322) );
  XOR2_X1 U379 ( .A(n322), .B(G211GAT), .Z(n410) );
  NAND2_X1 U380 ( .A1(G231GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U381 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n328) );
  INV_X1 U383 ( .A(n574), .ZN(n489) );
  XOR2_X1 U384 ( .A(G99GAT), .B(G106GAT), .Z(n352) );
  XOR2_X1 U385 ( .A(n352), .B(G218GAT), .Z(n331) );
  XNOR2_X1 U386 ( .A(G190GAT), .B(n442), .ZN(n330) );
  XNOR2_X1 U387 ( .A(n331), .B(n330), .ZN(n336) );
  XOR2_X1 U388 ( .A(KEYINPUT64), .B(KEYINPUT9), .Z(n333) );
  XNOR2_X1 U389 ( .A(G162GAT), .B(G92GAT), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U391 ( .A(n337), .B(KEYINPUT11), .ZN(n344) );
  XOR2_X1 U392 ( .A(n338), .B(KEYINPUT10), .Z(n342) );
  XOR2_X1 U393 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n340) );
  XNOR2_X1 U394 ( .A(G50GAT), .B(G36GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U396 ( .A(KEYINPUT7), .B(n341), .ZN(n371) );
  XNOR2_X1 U397 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n388), .B(n345), .ZN(n579) );
  NOR2_X1 U399 ( .A1(n489), .A2(n579), .ZN(n347) );
  INV_X1 U400 ( .A(KEYINPUT45), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n347), .B(n346), .ZN(n362) );
  XOR2_X1 U402 ( .A(G92GAT), .B(G64GAT), .Z(n405) );
  XOR2_X1 U403 ( .A(KEYINPUT74), .B(G85GAT), .Z(n349) );
  XNOR2_X1 U404 ( .A(G176GAT), .B(G120GAT), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U406 ( .A(n405), .B(n350), .Z(n354) );
  XNOR2_X1 U407 ( .A(G148GAT), .B(KEYINPUT75), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n351), .B(G204GAT), .ZN(n419) );
  XNOR2_X1 U409 ( .A(n419), .B(n352), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U411 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n356) );
  NAND2_X1 U412 ( .A1(G230GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U414 ( .A(n358), .B(n357), .Z(n361) );
  XNOR2_X1 U415 ( .A(n359), .B(KEYINPUT33), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n571) );
  NOR2_X1 U417 ( .A1(n362), .A2(n571), .ZN(n363) );
  XNOR2_X1 U418 ( .A(n363), .B(KEYINPUT109), .ZN(n385) );
  XOR2_X1 U419 ( .A(G141GAT), .B(G197GAT), .Z(n365) );
  XNOR2_X1 U420 ( .A(G29GAT), .B(G43GAT), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U422 ( .A(n366), .B(G113GAT), .Z(n369) );
  XNOR2_X1 U423 ( .A(G169GAT), .B(n367), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U425 ( .A(n371), .B(n370), .Z(n384) );
  XOR2_X1 U426 ( .A(KEYINPUT67), .B(G1GAT), .Z(n373) );
  XNOR2_X1 U427 ( .A(G8GAT), .B(KEYINPUT66), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U429 ( .A(KEYINPUT71), .B(KEYINPUT29), .Z(n375) );
  XNOR2_X1 U430 ( .A(KEYINPUT30), .B(KEYINPUT65), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U432 ( .A(n377), .B(n376), .Z(n382) );
  XOR2_X1 U433 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n379) );
  NAND2_X1 U434 ( .A1(G229GAT), .A2(G233GAT), .ZN(n378) );
  XNOR2_X1 U435 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U436 ( .A(KEYINPUT72), .B(n380), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U438 ( .A(n384), .B(n383), .Z(n503) );
  INV_X1 U439 ( .A(n503), .ZN(n568) );
  NOR2_X1 U440 ( .A1(n385), .A2(n568), .ZN(n387) );
  INV_X1 U441 ( .A(KEYINPUT110), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n394) );
  XOR2_X1 U443 ( .A(KEYINPUT41), .B(n571), .Z(n548) );
  NAND2_X1 U444 ( .A1(n568), .A2(n548), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n389), .B(KEYINPUT46), .ZN(n390) );
  XOR2_X1 U446 ( .A(KEYINPUT108), .B(n574), .Z(n558) );
  NAND2_X1 U447 ( .A1(n390), .A2(n558), .ZN(n391) );
  NOR2_X1 U448 ( .A1(n388), .A2(n391), .ZN(n392) );
  XNOR2_X1 U449 ( .A(KEYINPUT47), .B(n392), .ZN(n393) );
  NAND2_X1 U450 ( .A1(n394), .A2(n393), .ZN(n395) );
  INV_X1 U451 ( .A(n544), .ZN(n527) );
  XOR2_X1 U452 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n397) );
  XNOR2_X1 U453 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U455 ( .A(n398), .B(KEYINPUT82), .Z(n400) );
  XNOR2_X1 U456 ( .A(G169GAT), .B(G176GAT), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n438) );
  XOR2_X1 U458 ( .A(KEYINPUT21), .B(KEYINPUT86), .Z(n402) );
  XNOR2_X1 U459 ( .A(G197GAT), .B(G218GAT), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n420) );
  XOR2_X1 U461 ( .A(n420), .B(KEYINPUT96), .Z(n404) );
  NAND2_X1 U462 ( .A1(G226GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n406) );
  XOR2_X1 U464 ( .A(n406), .B(n405), .Z(n408) );
  XNOR2_X1 U465 ( .A(G36GAT), .B(G204GAT), .ZN(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n438), .B(n409), .ZN(n411) );
  INV_X1 U468 ( .A(n517), .ZN(n412) );
  NOR2_X1 U469 ( .A1(n527), .A2(n412), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U471 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n417) );
  NAND2_X1 U472 ( .A1(G228GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U474 ( .A(n418), .B(G211GAT), .Z(n422) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U477 ( .A(G155GAT), .B(G78GAT), .Z(n424) );
  XNOR2_X1 U478 ( .A(G50GAT), .B(G106GAT), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U480 ( .A(n426), .B(n425), .Z(n432) );
  XOR2_X1 U481 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n428) );
  XNOR2_X1 U482 ( .A(G22GAT), .B(KEYINPUT89), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n466) );
  NAND2_X1 U486 ( .A1(n567), .A2(n466), .ZN(n434) );
  XOR2_X1 U487 ( .A(KEYINPUT55), .B(KEYINPUT119), .Z(n433) );
  XNOR2_X1 U488 ( .A(n434), .B(n433), .ZN(n451) );
  XOR2_X1 U489 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n436) );
  XNOR2_X1 U490 ( .A(G71GAT), .B(G183GAT), .ZN(n435) );
  XNOR2_X1 U491 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n450) );
  XOR2_X1 U493 ( .A(G127GAT), .B(KEYINPUT20), .Z(n440) );
  XNOR2_X1 U494 ( .A(G15GAT), .B(G99GAT), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n442), .B(n441), .Z(n444) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U499 ( .A(n445), .B(KEYINPUT83), .Z(n448) );
  XNOR2_X1 U500 ( .A(n446), .B(KEYINPUT84), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n526) );
  NAND2_X1 U503 ( .A1(n451), .A2(n526), .ZN(n452) );
  XNOR2_X1 U504 ( .A(n452), .B(KEYINPUT120), .ZN(n559) );
  INV_X1 U505 ( .A(n559), .ZN(n556) );
  NAND2_X1 U506 ( .A1(n556), .A2(n388), .ZN(n455) );
  XOR2_X1 U507 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n453) );
  NAND2_X1 U508 ( .A1(n548), .A2(n556), .ZN(n459) );
  XOR2_X1 U509 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n457) );
  XOR2_X1 U510 ( .A(G176GAT), .B(KEYINPUT121), .Z(n456) );
  XNOR2_X1 U511 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U512 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  XOR2_X1 U513 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n479) );
  NOR2_X1 U514 ( .A1(n571), .A2(n503), .ZN(n460) );
  XOR2_X1 U515 ( .A(KEYINPUT76), .B(n460), .Z(n492) );
  NOR2_X1 U516 ( .A1(n388), .A2(n489), .ZN(n461) );
  XNOR2_X1 U517 ( .A(n461), .B(KEYINPUT16), .ZN(n476) );
  XNOR2_X1 U518 ( .A(KEYINPUT85), .B(n526), .ZN(n462) );
  XOR2_X1 U519 ( .A(n466), .B(KEYINPUT28), .Z(n521) );
  XNOR2_X1 U520 ( .A(KEYINPUT27), .B(n517), .ZN(n468) );
  NAND2_X1 U521 ( .A1(n515), .A2(n468), .ZN(n546) );
  NOR2_X1 U522 ( .A1(n521), .A2(n546), .ZN(n525) );
  NAND2_X1 U523 ( .A1(n462), .A2(n525), .ZN(n475) );
  NAND2_X1 U524 ( .A1(n517), .A2(n526), .ZN(n463) );
  NAND2_X1 U525 ( .A1(n463), .A2(n466), .ZN(n464) );
  XNOR2_X1 U526 ( .A(n464), .B(KEYINPUT25), .ZN(n465) );
  XOR2_X1 U527 ( .A(KEYINPUT98), .B(n465), .Z(n471) );
  NOR2_X1 U528 ( .A1(n466), .A2(n526), .ZN(n467) );
  XNOR2_X1 U529 ( .A(n467), .B(KEYINPUT26), .ZN(n566) );
  NAND2_X1 U530 ( .A1(n566), .A2(n468), .ZN(n469) );
  XOR2_X1 U531 ( .A(KEYINPUT97), .B(n469), .Z(n470) );
  NAND2_X1 U532 ( .A1(n471), .A2(n470), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n473), .A2(n472), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n488) );
  NAND2_X1 U535 ( .A1(n476), .A2(n488), .ZN(n504) );
  NOR2_X1 U536 ( .A1(n492), .A2(n504), .ZN(n477) );
  XOR2_X1 U537 ( .A(KEYINPUT99), .B(n477), .Z(n485) );
  NAND2_X1 U538 ( .A1(n485), .A2(n515), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U540 ( .A(G1GAT), .B(n480), .Z(G1324GAT) );
  NAND2_X1 U541 ( .A1(n485), .A2(n517), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n483) );
  NAND2_X1 U544 ( .A1(n485), .A2(n526), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U546 ( .A(G15GAT), .B(n484), .Z(G1326GAT) );
  NAND2_X1 U547 ( .A1(n485), .A2(n521), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n486), .B(KEYINPUT102), .ZN(n487) );
  XNOR2_X1 U549 ( .A(G22GAT), .B(n487), .ZN(G1327GAT) );
  XOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .Z(n495) );
  NAND2_X1 U551 ( .A1(n489), .A2(n488), .ZN(n490) );
  NOR2_X1 U552 ( .A1(n490), .A2(n579), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(KEYINPUT37), .ZN(n514) );
  NOR2_X1 U554 ( .A1(n492), .A2(n514), .ZN(n493) );
  XNOR2_X1 U555 ( .A(KEYINPUT38), .B(n493), .ZN(n501) );
  NAND2_X1 U556 ( .A1(n501), .A2(n515), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n501), .A2(n517), .ZN(n496) );
  XNOR2_X1 U559 ( .A(n496), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U560 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n500) );
  XOR2_X1 U561 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n498) );
  NAND2_X1 U562 ( .A1(n526), .A2(n501), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(G1330GAT) );
  NAND2_X1 U565 ( .A1(n501), .A2(n521), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n502), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n506) );
  NAND2_X1 U568 ( .A1(n548), .A2(n503), .ZN(n513) );
  NAND2_X1 U569 ( .A1(n510), .A2(n515), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n510), .A2(n517), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n510), .A2(n526), .ZN(n508) );
  XNOR2_X1 U574 ( .A(n508), .B(KEYINPUT106), .ZN(n509) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(n509), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U577 ( .A1(n510), .A2(n521), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  NOR2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n522) );
  NAND2_X1 U580 ( .A1(n522), .A2(n515), .ZN(n516) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  XOR2_X1 U582 ( .A(G92GAT), .B(KEYINPUT107), .Z(n519) );
  NAND2_X1 U583 ( .A1(n522), .A2(n517), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n519), .B(n518), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n522), .A2(n526), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  XOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT113), .Z(n531) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n528) );
  NOR2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U593 ( .A(n529), .B(KEYINPUT112), .Z(n535) );
  INV_X1 U594 ( .A(n535), .ZN(n539) );
  NAND2_X1 U595 ( .A1(n568), .A2(n539), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n533) );
  NAND2_X1 U598 ( .A1(n548), .A2(n539), .ZN(n532) );
  XNOR2_X1 U599 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U600 ( .A(G120GAT), .B(n534), .ZN(G1341GAT) );
  NOR2_X1 U601 ( .A1(n535), .A2(n558), .ZN(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U606 ( .A1(n388), .A2(n539), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n543) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT117), .Z(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n544), .A2(n566), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n568), .A2(n554), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n552) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U616 ( .A1(n554), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n574), .A2(n554), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U621 ( .A1(n554), .A2(n388), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n555), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U623 ( .A1(n568), .A2(n556), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(n557), .ZN(G1348GAT) );
  INV_X1 U625 ( .A(KEYINPUT122), .ZN(n561) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G183GAT), .B(n562), .ZN(G1350GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n564) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT124), .B(n565), .Z(n570) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n578) );
  INV_X1 U634 ( .A(n578), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n575), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U638 ( .A1(n575), .A2(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  XNOR2_X1 U640 ( .A(G211GAT), .B(KEYINPUT126), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

