//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(new_n208), .A2(new_n209), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  INV_X1    g0019(.A(G97), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n216), .B1(new_n209), .B2(new_n208), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT64), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n235), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G20), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G77), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n252), .B1(new_n214), .B2(G68), .C1(new_n254), .C2(new_n202), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n213), .B1(new_n206), .B2(new_n250), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT11), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT68), .A2(G1), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT68), .A2(G1), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G68), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT12), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n256), .B1(new_n261), .B2(G20), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G68), .ZN(new_n268));
  XOR2_X1   g0068(.A(new_n268), .B(KEYINPUT71), .Z(new_n269));
  NAND3_X1  g0069(.A1(new_n258), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G226), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G97), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G41), .A2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(G274), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n280), .B1(new_n283), .B2(new_n261), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(new_n287), .B2(G238), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT13), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT13), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n281), .A2(new_n291), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G200), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n290), .A2(new_n296), .A3(new_n292), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n270), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n267), .A2(G77), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(G77), .B2(new_n262), .ZN(new_n300));
  INV_X1    g0100(.A(new_n256), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT15), .B(G87), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  AOI22_X1  g0103(.A1(new_n303), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n304));
  XNOR2_X1  g0104(.A(KEYINPUT8), .B(G58), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n254), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n301), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n300), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n274), .A2(G232), .A3(new_n275), .ZN(new_n310));
  INV_X1    g0110(.A(G107), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n274), .A2(G1698), .ZN(new_n312));
  INV_X1    g0112(.A(G238), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n310), .B1(new_n311), .B2(new_n274), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n280), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n286), .B1(new_n287), .B2(G244), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n317), .A2(G190), .ZN(new_n318));
  AOI21_X1  g0118(.A(G200), .B1(new_n315), .B2(new_n316), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n309), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n309), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n315), .A2(G179), .A3(new_n316), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n315), .B2(new_n316), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n321), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n324), .B1(new_n290), .B2(new_n292), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n329), .A2(KEYINPUT72), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n328), .A2(new_n331), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n290), .A2(G179), .A3(new_n292), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI211_X1 g0135(.A(new_n298), .B(new_n327), .C1(new_n335), .C2(new_n270), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n287), .A2(G226), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n285), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n274), .A2(G222), .A3(new_n275), .ZN(new_n339));
  INV_X1    g0139(.A(G223), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n339), .B1(new_n225), .B2(new_n274), .C1(new_n312), .C2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n338), .B1(new_n341), .B2(new_n280), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(new_n294), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT70), .B1(new_n342), .B2(G190), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n342), .A2(KEYINPUT70), .A3(G190), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n267), .A2(G50), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(G50), .B2(new_n262), .ZN(new_n349));
  INV_X1    g0149(.A(new_n305), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n251), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n253), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n301), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT9), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT69), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n347), .B(new_n356), .C1(new_n357), .C2(KEYINPUT10), .ZN(new_n358));
  INV_X1    g0158(.A(new_n343), .ZN(new_n359));
  INV_X1    g0159(.A(new_n346), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n356), .B(new_n359), .C1(new_n360), .C2(new_n344), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n357), .B(new_n359), .C1(new_n360), .C2(new_n344), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT10), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n342), .A2(G179), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n324), .B2(new_n342), .ZN(new_n366));
  INV_X1    g0166(.A(new_n354), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n358), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n336), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n262), .A2(new_n305), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n267), .B2(new_n305), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(G58), .A2(G68), .ZN(new_n374));
  OAI21_X1  g0174(.A(G20), .B1(new_n374), .B2(new_n201), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g0177(.A(KEYINPUT75), .B(G20), .C1(new_n374), .C2(new_n201), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n253), .A2(G159), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT73), .B1(new_n250), .B2(KEYINPUT3), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(new_n271), .A3(G33), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n383), .A3(new_n273), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n214), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n264), .B1(new_n385), .B2(KEYINPUT7), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(KEYINPUT74), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT74), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n381), .A2(new_n383), .A3(new_n388), .A4(new_n273), .ZN(new_n389));
  NOR2_X1   g0189(.A1(KEYINPUT7), .A2(G20), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n380), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n301), .B1(new_n392), .B2(KEYINPUT16), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n274), .B2(G20), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n272), .A2(new_n273), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n264), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n394), .B1(new_n399), .B2(new_n380), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n373), .B1(new_n393), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G41), .ZN(new_n402));
  OAI211_X1 g0202(.A(G1), .B(G13), .C1(new_n250), .C2(new_n402), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT68), .B(G1), .ZN(new_n404));
  OAI211_X1 g0204(.A(G232), .B(new_n403), .C1(new_n404), .C2(new_n282), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n405), .A2(KEYINPUT77), .A3(new_n285), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT77), .B1(new_n405), .B2(new_n285), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT78), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n405), .A2(new_n285), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT77), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n405), .A2(KEYINPUT77), .A3(new_n285), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  MUX2_X1   g0214(.A(new_n340), .B(new_n224), .S(G1698), .Z(new_n415));
  OAI22_X1  g0215(.A1(new_n384), .A2(new_n415), .B1(new_n250), .B2(new_n218), .ZN(new_n416));
  AOI21_X1  g0216(.A(G190), .B1(new_n416), .B2(new_n280), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n408), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n280), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n411), .A2(new_n413), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n294), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n401), .A2(KEYINPUT17), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT17), .B1(new_n401), .B2(new_n422), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(G179), .B1(new_n416), .B2(new_n280), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n408), .A2(new_n414), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n420), .A2(new_n324), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n386), .A2(new_n391), .ZN(new_n430));
  INV_X1    g0230(.A(new_n380), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(KEYINPUT16), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(new_n400), .A3(new_n256), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n372), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(new_n434), .A3(KEYINPUT18), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n427), .A2(new_n428), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n436), .B1(new_n401), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n425), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(KEYINPUT79), .B1(new_n370), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT79), .ZN(new_n442));
  INV_X1    g0242(.A(new_n440), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n336), .A2(new_n369), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n441), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n261), .A2(G33), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n262), .A2(new_n447), .A3(G116), .A4(new_n301), .ZN(new_n448));
  INV_X1    g0248(.A(G116), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n261), .A2(G13), .A3(G20), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(G20), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n256), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT86), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT86), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n256), .A2(new_n456), .A3(new_n453), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(G20), .B1(G33), .B2(G283), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(G33), .B2(new_n220), .ZN(new_n460));
  AOI21_X1  g0260(.A(KEYINPUT20), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n256), .A2(new_n456), .A3(new_n453), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n456), .B1(new_n256), .B2(new_n453), .ZN(new_n463));
  OAI211_X1 g0263(.A(KEYINPUT20), .B(new_n460), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n452), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  OR2_X1    g0266(.A1(KEYINPUT68), .A2(G1), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G41), .ZN(new_n469));
  NAND2_X1  g0269(.A1(KEYINPUT68), .A2(G1), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n467), .A2(new_n469), .A3(G45), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT84), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT84), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n261), .A2(new_n473), .A3(G45), .A4(new_n469), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n402), .A2(KEYINPUT5), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(G270), .A3(new_n403), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n403), .A2(G274), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n474), .A2(new_n472), .A3(new_n478), .A4(new_n475), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n221), .A2(G1698), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(G264), .B2(G1698), .ZN(new_n481));
  XOR2_X1   g0281(.A(KEYINPUT85), .B(G303), .Z(new_n482));
  OAI22_X1  g0282(.A1(new_n481), .A2(new_n384), .B1(new_n274), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n280), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n477), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n466), .A2(new_n485), .A3(G169), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT21), .ZN(new_n487));
  AND3_X1   g0287(.A1(new_n486), .A2(KEYINPUT87), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n487), .B1(new_n486), .B2(KEYINPUT87), .ZN(new_n489));
  INV_X1    g0289(.A(G179), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n491), .A2(new_n466), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n488), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n485), .A2(G190), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n294), .B2(new_n485), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n495), .A2(new_n466), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT19), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n214), .B1(new_n278), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G87), .A2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n311), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n214), .A2(G33), .A3(G97), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n499), .A2(new_n501), .B1(new_n498), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n381), .A2(new_n383), .A3(new_n214), .A4(new_n273), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n264), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n256), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n262), .A2(new_n447), .A3(new_n301), .A4(new_n303), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n262), .A2(new_n303), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G244), .A2(G1698), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n313), .B2(G1698), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n512), .A2(new_n381), .A3(new_n383), .A4(new_n273), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n403), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n219), .B1(new_n261), .B2(G45), .ZN(new_n517));
  AND4_X1   g0317(.A1(G45), .A2(new_n467), .A3(G274), .A4(new_n470), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n403), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(new_n519), .A3(new_n490), .ZN(new_n520));
  INV_X1    g0320(.A(G45), .ZN(new_n521));
  OAI21_X1  g0321(.A(G250), .B1(new_n404), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n261), .A2(G45), .A3(G274), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n280), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n324), .B1(new_n524), .B2(new_n515), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n510), .A2(new_n520), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n516), .A2(new_n519), .A3(G190), .ZN(new_n527));
  OAI21_X1  g0327(.A(G200), .B1(new_n524), .B2(new_n515), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n262), .A2(new_n301), .A3(new_n447), .ZN(new_n529));
  OR2_X1    g0329(.A1(new_n529), .A2(new_n218), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n508), .B1(new_n505), .B2(new_n256), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n527), .A2(new_n528), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n476), .A2(G257), .A3(new_n403), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n226), .A2(G1698), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n381), .A2(new_n383), .A3(new_n273), .A4(new_n535), .ZN(new_n536));
  XNOR2_X1  g0336(.A(KEYINPUT83), .B(KEYINPUT4), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n272), .A2(new_n273), .A3(G250), .A4(G1698), .ZN(new_n539));
  AND2_X1   g0339(.A1(KEYINPUT4), .A2(G244), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n272), .A2(new_n273), .A3(new_n540), .A4(new_n275), .ZN(new_n541));
  INV_X1    g0341(.A(G283), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n539), .B(new_n541), .C1(new_n250), .C2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n280), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n534), .A2(new_n544), .A3(new_n479), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n294), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n534), .A2(new_n544), .A3(new_n296), .A4(new_n479), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n396), .A2(new_n398), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G107), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n253), .A2(G77), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT6), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n220), .A2(new_n311), .ZN(new_n553));
  NOR2_X1   g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT80), .ZN(new_n556));
  NAND2_X1  g0356(.A1(KEYINPUT6), .A2(G97), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n556), .B1(new_n557), .B2(G107), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n311), .A2(KEYINPUT80), .A3(KEYINPUT6), .A4(G97), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT81), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT81), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n555), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n550), .B(new_n551), .C1(new_n565), .C2(new_n214), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n262), .A2(new_n447), .A3(G97), .A4(new_n301), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(G97), .B2(new_n262), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT82), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT82), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n567), .B(new_n570), .C1(G97), .C2(new_n262), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n566), .A2(new_n256), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n533), .B1(new_n548), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n545), .A2(G169), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n490), .B2(new_n545), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n566), .A2(new_n256), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n569), .A2(new_n571), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n476), .A2(G264), .A3(new_n403), .ZN(new_n581));
  MUX2_X1   g0381(.A(new_n219), .B(new_n221), .S(G1698), .Z(new_n582));
  INV_X1    g0382(.A(G294), .ZN(new_n583));
  OAI22_X1  g0383(.A1(new_n384), .A2(new_n582), .B1(new_n250), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n280), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n581), .A2(new_n479), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(new_n490), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT90), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT90), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n586), .B2(G169), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n588), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n529), .A2(new_n311), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT25), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n263), .B2(new_n311), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n262), .A2(KEYINPUT25), .A3(G107), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT23), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n214), .B2(G107), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n311), .A2(KEYINPUT23), .A3(G20), .ZN(new_n599));
  INV_X1    g0399(.A(new_n514), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n598), .A2(new_n599), .B1(new_n600), .B2(new_n214), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT22), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(new_n214), .A3(G87), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT88), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n604), .A2(new_n605), .A3(new_n272), .A4(new_n273), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT88), .B1(new_n397), .B2(new_n603), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT22), .B1(new_n504), .B2(new_n218), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT89), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n610), .B1(new_n608), .B2(new_n609), .ZN(new_n613));
  OAI211_X1 g0413(.A(KEYINPUT24), .B(new_n601), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n256), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n608), .A2(new_n609), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT89), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n611), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT24), .B1(new_n618), .B2(new_n601), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n596), .B1(new_n615), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n591), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n586), .A2(new_n294), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n581), .A2(new_n296), .A3(new_n479), .A4(new_n585), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n624), .B(new_n596), .C1(new_n615), .C2(new_n619), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n580), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n446), .A2(new_n497), .A3(new_n626), .ZN(G372));
  INV_X1    g0427(.A(KEYINPUT91), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT18), .B1(new_n429), .B2(new_n434), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n401), .A2(new_n437), .A3(new_n436), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n435), .A2(new_n438), .A3(KEYINPUT91), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n298), .ZN(new_n634));
  INV_X1    g0434(.A(new_n325), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n309), .B1(new_n635), .B2(new_n322), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n335), .A2(new_n270), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n425), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n358), .A2(new_n364), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n639), .A2(new_n640), .B1(new_n367), .B2(new_n366), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n489), .A2(new_n492), .ZN(new_n642));
  INV_X1    g0442(.A(new_n488), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n621), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n625), .A2(new_n573), .A3(new_n579), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT26), .B1(new_n579), .B2(new_n533), .ZN(new_n648));
  INV_X1    g0448(.A(new_n533), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n649), .A2(new_n575), .A3(new_n578), .A4(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n648), .A2(new_n526), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n641), .B1(new_n446), .B2(new_n654), .ZN(G369));
  NAND2_X1  g0455(.A1(new_n642), .A2(new_n643), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n214), .A2(G13), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n261), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G343), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n466), .ZN(new_n665));
  XOR2_X1   g0465(.A(new_n665), .B(KEYINPUT92), .Z(new_n666));
  NOR2_X1   g0466(.A1(new_n656), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n497), .B2(new_n666), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(G330), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n621), .A2(new_n663), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n621), .A2(new_n625), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n620), .A2(new_n664), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n656), .A2(new_n663), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(new_n671), .A3(new_n672), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n621), .B2(new_n664), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n674), .A2(new_n678), .ZN(G399));
  NAND3_X1  g0479(.A1(new_n500), .A2(new_n311), .A3(new_n449), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n207), .A2(new_n402), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n682), .A3(G1), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n211), .B2(new_n682), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT93), .Z(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n664), .B1(new_n647), .B2(new_n652), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n688), .A2(KEYINPUT29), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n688), .A2(KEYINPUT29), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n524), .A2(new_n515), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G179), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n485), .A2(new_n545), .A3(new_n586), .A4(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n581), .A2(new_n692), .A3(new_n585), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n696), .A2(new_n545), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n697), .A2(new_n491), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(KEYINPUT94), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT30), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n698), .B2(KEYINPUT94), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n695), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT31), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n700), .A2(new_n702), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n694), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n705), .B1(new_n707), .B2(new_n664), .ZN(new_n708));
  INV_X1    g0508(.A(new_n497), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n671), .A3(new_n580), .A4(new_n663), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n704), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G330), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n691), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n686), .B1(new_n713), .B2(new_n284), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT95), .Z(G364));
  NAND2_X1  g0515(.A1(new_n657), .A2(G45), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n682), .A2(new_n716), .A3(G1), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n669), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n668), .A2(G330), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G13), .A2(G33), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n668), .A2(G20), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n213), .B1(G20), .B2(new_n324), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n214), .A2(new_n296), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(G179), .A3(new_n294), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G322), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n214), .A2(G190), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n729), .A2(new_n490), .A3(G200), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(G311), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n727), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n490), .A2(new_n294), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n728), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT33), .B(G317), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n274), .B(new_n733), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n294), .A2(G179), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n728), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n728), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI22_X1  g0544(.A1(G283), .A2(new_n741), .B1(new_n744), .B2(G329), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n734), .A2(new_n724), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n724), .A2(new_n739), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(G326), .A2(new_n747), .B1(new_n749), .B2(G303), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n742), .A2(G190), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G294), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n738), .A2(new_n745), .A3(new_n750), .A4(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT97), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n274), .B1(new_n731), .B2(new_n225), .ZN(new_n756));
  INV_X1    g0556(.A(new_n752), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n220), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n746), .A2(new_n202), .B1(new_n735), .B2(new_n264), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G159), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n743), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT32), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n740), .A2(new_n311), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n748), .A2(new_n218), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n764), .B(new_n765), .C1(G58), .C2(new_n726), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n760), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n754), .B1(new_n755), .B2(new_n767), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n767), .A2(new_n755), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n723), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n721), .A2(G20), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n723), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n387), .A2(new_n389), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n207), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n244), .A2(G45), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n211), .A2(new_n521), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n274), .A2(new_n207), .ZN(new_n779));
  INV_X1    g0579(.A(G355), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n779), .A2(new_n780), .B1(G116), .B2(new_n207), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT96), .Z(new_n782));
  OAI21_X1  g0582(.A(new_n772), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n717), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n770), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n718), .A2(new_n719), .B1(new_n722), .B2(new_n785), .ZN(G396));
  NAND2_X1  g0586(.A1(new_n664), .A2(new_n321), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n636), .B1(new_n320), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n326), .A2(new_n664), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OR3_X1    g0590(.A1(new_n687), .A2(KEYINPUT98), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n645), .B1(new_n493), .B2(new_n621), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n648), .A2(new_n526), .A3(new_n651), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n663), .B(new_n790), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(KEYINPUT98), .B1(new_n687), .B2(new_n790), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n707), .A2(new_n705), .A3(new_n664), .ZN(new_n798));
  OAI21_X1  g0598(.A(KEYINPUT31), .B1(new_n703), .B2(new_n663), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n626), .A2(new_n497), .A3(new_n664), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G330), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n784), .B1(new_n797), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n803), .B2(new_n797), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n723), .A2(new_n720), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n717), .B1(new_n225), .B2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n723), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G107), .A2(new_n749), .B1(new_n744), .B2(G311), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n809), .B(new_n397), .C1(new_n218), .C2(new_n740), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n731), .A2(new_n449), .B1(new_n583), .B2(new_n725), .ZN(new_n811));
  INV_X1    g0611(.A(G303), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n746), .A2(new_n812), .B1(new_n735), .B2(new_n542), .ZN(new_n813));
  NOR4_X1   g0613(.A1(new_n810), .A2(new_n811), .A3(new_n758), .A4(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n726), .A2(G143), .B1(new_n736), .B2(G150), .ZN(new_n815));
  INV_X1    g0615(.A(G137), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n815), .B1(new_n816), .B2(new_n746), .C1(new_n761), .C2(new_n731), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT34), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G50), .A2(new_n749), .B1(new_n741), .B2(G68), .ZN(new_n819));
  INV_X1    g0619(.A(G132), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n820), .B2(new_n743), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n774), .B(new_n821), .C1(G58), .C2(new_n752), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n814), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n807), .B1(new_n808), .B2(new_n823), .C1(new_n790), .C2(new_n721), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n805), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(G384));
  INV_X1    g0626(.A(KEYINPUT35), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n565), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n562), .A2(KEYINPUT35), .A3(new_n564), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n828), .A2(G116), .A3(new_n215), .A4(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT36), .Z(new_n831));
  OR3_X1    g0631(.A1(new_n211), .A2(new_n225), .A3(new_n374), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n202), .A2(G68), .ZN(new_n833));
  AOI211_X1 g0633(.A(G13), .B(new_n261), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n788), .A2(new_n789), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n270), .B(new_n664), .C1(new_n335), .C2(new_n298), .ZN(new_n837));
  INV_X1    g0637(.A(new_n333), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n334), .B1(new_n328), .B2(new_n331), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n270), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n270), .A2(new_n664), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n840), .A2(new_n634), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n836), .B1(new_n837), .B2(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n394), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n392), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n373), .B1(new_n847), .B2(new_n393), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(new_n661), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n440), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n432), .A2(new_n256), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n392), .A2(new_n846), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n372), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI22_X1  g0654(.A1(new_n854), .A2(new_n429), .B1(new_n401), .B2(new_n422), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n849), .B1(new_n855), .B2(KEYINPUT100), .ZN(new_n856));
  INV_X1    g0656(.A(new_n422), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n857), .A2(new_n434), .B1(new_n848), .B2(new_n437), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT100), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n851), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT37), .B1(new_n429), .B2(new_n434), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n401), .A2(new_n422), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT101), .B1(new_n434), .B2(new_n662), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT101), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n865), .B(new_n661), .C1(new_n433), .C2(new_n372), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n862), .B(new_n863), .C1(new_n864), .C2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT38), .B(new_n850), .C1(new_n861), .C2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n864), .A2(new_n866), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n631), .A2(new_n425), .A3(new_n632), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n429), .A2(new_n434), .A3(KEYINPUT91), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n628), .B1(new_n401), .B2(new_n437), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n870), .A2(new_n871), .B1(new_n876), .B2(new_n867), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n869), .B1(new_n877), .B2(KEYINPUT38), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n845), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n856), .A2(new_n860), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n868), .B1(new_n881), .B2(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(new_n849), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n425), .B2(new_n439), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n880), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT40), .B1(new_n885), .B2(new_n869), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n879), .A2(KEYINPUT40), .B1(new_n845), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n445), .A2(new_n711), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n889), .A2(new_n802), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n885), .A2(new_n869), .ZN(new_n891));
  INV_X1    g0691(.A(new_n789), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n794), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n837), .A2(new_n842), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(KEYINPUT99), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT99), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n893), .B2(new_n894), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n891), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n840), .A2(new_n664), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT39), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n869), .B(new_n901), .C1(new_n877), .C2(KEYINPUT38), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n901), .B1(new_n885), .B2(new_n869), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n633), .A2(new_n662), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n899), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n445), .B1(new_n689), .B2(new_n690), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n908), .A2(new_n641), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n907), .B(new_n909), .ZN(new_n910));
  OAI22_X1  g0710(.A1(new_n890), .A2(new_n910), .B1(new_n261), .B2(new_n657), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n890), .A2(new_n910), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n835), .B1(new_n911), .B2(new_n912), .ZN(G367));
  NOR2_X1   g0713(.A1(new_n572), .A2(new_n663), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n572), .B2(new_n548), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n579), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n677), .A2(new_n916), .ZN(new_n917));
  OR3_X1    g0717(.A1(new_n917), .A2(KEYINPUT103), .A3(KEYINPUT42), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT103), .B1(new_n917), .B2(KEYINPUT42), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n579), .B1(new_n916), .B2(new_n621), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n917), .A2(KEYINPUT42), .B1(new_n920), .B2(new_n663), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT43), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n530), .A2(new_n531), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n664), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n649), .A2(KEYINPUT102), .A3(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n526), .B2(new_n925), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT102), .B1(new_n649), .B2(new_n925), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n922), .B1(new_n923), .B2(new_n929), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n927), .A2(KEYINPUT43), .A3(new_n928), .ZN(new_n931));
  OR2_X1    g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  INV_X1    g0733(.A(new_n674), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n579), .A2(new_n663), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n915), .B2(new_n579), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g0737(.A1(new_n932), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n937), .B1(new_n932), .B2(new_n933), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n682), .B(KEYINPUT41), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n678), .A2(new_n936), .ZN(new_n942));
  NOR2_X1   g0742(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  AND2_X1   g0744(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n678), .A2(new_n936), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT45), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n674), .A2(KEYINPUT105), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n947), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  OAI211_X1 g0752(.A(KEYINPUT105), .B(new_n674), .C1(new_n946), .C2(new_n949), .ZN(new_n953));
  INV_X1    g0753(.A(new_n713), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n669), .A2(new_n673), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n934), .A2(new_n676), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n676), .B1(new_n934), .B2(new_n955), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n952), .A2(new_n953), .A3(new_n954), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n941), .B1(new_n959), .B2(new_n954), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n716), .A2(G1), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n940), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n929), .A2(new_n771), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n740), .A2(new_n225), .B1(new_n743), .B2(new_n816), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n397), .B(new_n964), .C1(G58), .C2(new_n749), .ZN(new_n965));
  AOI22_X1  g0765(.A1(new_n730), .A2(G50), .B1(new_n736), .B2(G159), .ZN(new_n966));
  AOI22_X1  g0766(.A1(new_n726), .A2(G150), .B1(new_n747), .B2(G143), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n752), .A2(G68), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n749), .A2(G116), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT46), .ZN(new_n971));
  INV_X1    g0771(.A(G317), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n743), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n740), .A2(new_n220), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(G107), .C2(new_n752), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n730), .A2(G283), .B1(new_n736), .B2(G294), .ZN(new_n976));
  INV_X1    g0776(.A(new_n482), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n977), .A2(new_n726), .B1(new_n747), .B2(G311), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n971), .A2(new_n975), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n969), .B1(new_n979), .B2(new_n773), .ZN(new_n980));
  XNOR2_X1  g0780(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n808), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n980), .B2(new_n981), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n772), .B1(new_n207), .B2(new_n302), .C1(new_n239), .C2(new_n775), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n963), .A2(new_n784), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n962), .A2(new_n985), .ZN(G387));
  OAI22_X1  g0786(.A1(new_n725), .A2(new_n972), .B1(new_n735), .B2(new_n732), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n731), .A2(new_n482), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(G322), .C2(new_n747), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n989), .A2(KEYINPUT48), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(KEYINPUT48), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n749), .A2(G294), .B1(new_n752), .B2(G283), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(KEYINPUT107), .B(KEYINPUT49), .Z(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n744), .A2(G326), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n741), .A2(G116), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n995), .A2(new_n774), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n731), .A2(new_n264), .B1(new_n202), .B2(new_n725), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n974), .B(new_n999), .C1(new_n350), .C2(new_n736), .ZN(new_n1000));
  INV_X1    g0800(.A(G150), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n748), .A2(new_n225), .B1(new_n743), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G159), .B2(new_n747), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n303), .A2(new_n752), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1000), .A2(new_n773), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n808), .B1(new_n998), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n305), .A2(G50), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT50), .ZN(new_n1008));
  AOI211_X1 g0808(.A(G45), .B(new_n680), .C1(G68), .C2(G77), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n775), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n235), .B2(new_n521), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(G107), .B2(new_n207), .C1(new_n681), .C2(new_n779), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n717), .B(new_n1006), .C1(new_n772), .C2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT108), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n673), .A2(new_n771), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1014), .A2(new_n1015), .B1(new_n958), .B2(new_n961), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n958), .A2(new_n954), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n713), .B1(new_n956), .B2(new_n957), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n682), .B(KEYINPUT109), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1016), .A2(new_n1020), .ZN(G393));
  NAND3_X1  g0821(.A1(new_n947), .A2(new_n674), .A3(new_n950), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n934), .B1(new_n946), .B2(new_n949), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1022), .A2(new_n1017), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n959), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n752), .A2(G77), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n202), .B2(new_n735), .C1(new_n218), .C2(new_n740), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n731), .A2(new_n305), .B1(new_n264), .B2(new_n748), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(G143), .C2(new_n744), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n725), .A2(new_n761), .B1(new_n746), .B2(new_n1001), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1029), .A2(new_n773), .A3(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n725), .A2(new_n732), .B1(new_n746), .B2(new_n972), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT52), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n977), .A2(new_n736), .B1(new_n744), .B2(G322), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n730), .A2(G294), .B1(new_n749), .B2(G283), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n274), .B(new_n764), .C1(G116), .C2(new_n752), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n808), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n772), .B1(new_n220), .B2(new_n207), .C1(new_n248), .C2(new_n775), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n784), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1040), .B(new_n1042), .C1(new_n936), .C2(new_n771), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n961), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1025), .A2(new_n1045), .ZN(G390));
  INV_X1    g0846(.A(new_n894), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n712), .B2(new_n836), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n711), .A2(G330), .A3(new_n843), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT112), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1048), .B(new_n1049), .C1(new_n1050), .C2(new_n893), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n893), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n894), .B1(new_n803), .B2(new_n790), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1049), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n445), .A2(G330), .A3(new_n711), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n908), .A2(new_n1056), .A3(new_n641), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n1051), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n883), .B1(new_n858), .B2(new_n859), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n855), .A2(KEYINPUT100), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT37), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n867), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT38), .B1(new_n1062), .B2(new_n850), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n869), .ZN(new_n1064));
  OAI21_X1  g0864(.A(KEYINPUT39), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n900), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n789), .B1(new_n687), .B2(new_n790), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1066), .B1(new_n1067), .B2(new_n1047), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1065), .A2(new_n1068), .A3(new_n902), .ZN(new_n1069));
  AND4_X1   g0869(.A1(KEYINPUT111), .A2(new_n895), .A3(new_n878), .A4(new_n1066), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n900), .B1(new_n893), .B2(new_n894), .ZN(new_n1071));
  AOI21_X1  g0871(.A(KEYINPUT111), .B1(new_n1071), .B2(new_n878), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1069), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n1054), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1069), .B(new_n1049), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1058), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n1019), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1051), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT113), .ZN(new_n1079));
  AND3_X1   g0879(.A1(new_n1074), .A2(new_n1079), .A3(new_n1075), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1079), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT114), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1071), .A2(new_n878), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT111), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1071), .A2(KEYINPUT111), .A3(new_n878), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1049), .B1(new_n1089), .B2(new_n1069), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1075), .ZN(new_n1091));
  OAI21_X1  g0891(.A(KEYINPUT113), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1074), .A2(new_n1079), .A3(new_n1075), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(KEYINPUT114), .A3(new_n1078), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1077), .B1(new_n1084), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1074), .A2(new_n961), .A3(new_n1075), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1065), .A2(new_n720), .A3(new_n902), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n806), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n784), .B1(new_n350), .B2(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n731), .A2(new_n220), .B1(new_n740), .B2(new_n264), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n1101), .A2(new_n274), .A3(new_n765), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G283), .A2(new_n747), .B1(new_n736), .B2(G107), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n726), .A2(G116), .B1(new_n744), .B2(G294), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1102), .A2(new_n1026), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT54), .B(G143), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n731), .A2(new_n1106), .B1(new_n816), .B2(new_n735), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G159), .B2(new_n752), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT115), .ZN(new_n1109));
  INV_X1    g0909(.A(G128), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n725), .A2(new_n820), .B1(new_n746), .B2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT117), .Z(new_n1112));
  NAND3_X1  g0912(.A1(new_n749), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT53), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n748), .B2(new_n1001), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1113), .A2(new_n1115), .B1(G125), .B2(new_n744), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n274), .B1(new_n740), .B2(new_n202), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT116), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1112), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1105), .B1(new_n1109), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1100), .B1(new_n1120), .B2(new_n723), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1098), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1097), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1096), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(G378));
  NAND2_X1  g0925(.A1(new_n1076), .A2(new_n1057), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n367), .A2(new_n662), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n369), .B(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1128), .B(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT120), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n907), .A2(new_n1133), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1132), .A2(new_n899), .A3(new_n905), .A4(new_n906), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n887), .A2(new_n802), .B1(new_n1131), .B2(new_n1130), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT57), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1126), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1126), .B2(new_n1141), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1019), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1137), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n961), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1130), .A2(new_n720), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n730), .A2(G137), .B1(new_n736), .B2(G132), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT119), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n748), .A2(new_n1106), .ZN(new_n1152));
  INV_X1    g0952(.A(G125), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n725), .A2(new_n1110), .B1(new_n746), .B2(new_n1153), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(G150), .C2(new_n752), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1151), .A2(new_n1155), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n744), .A2(G124), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G33), .B(G41), .C1(new_n741), .C2(G159), .ZN(new_n1160));
  AND4_X1   g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n730), .A2(new_n303), .B1(new_n749), .B2(G77), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G116), .A2(new_n747), .B1(new_n736), .B2(G97), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n726), .A2(G107), .B1(new_n744), .B2(G283), .ZN(new_n1164));
  AND4_X1   g0964(.A1(new_n968), .A2(new_n1162), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n773), .A2(G41), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n741), .A2(G58), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT118), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT58), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1166), .ZN(new_n1171));
  AOI21_X1  g0971(.A(G50), .B1(new_n250), .B2(new_n402), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1169), .A2(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n1170), .B2(new_n1169), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n723), .B1(new_n1161), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n717), .B1(new_n202), .B2(new_n806), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1149), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1148), .A2(KEYINPUT121), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT121), .B1(new_n1148), .B2(new_n1177), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1145), .A2(new_n1180), .ZN(G375));
  NAND2_X1  g0981(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(G1), .B2(new_n716), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1047), .A2(new_n720), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n784), .B1(G68), .B2(new_n1099), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n725), .A2(new_n542), .B1(new_n748), .B2(new_n220), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n274), .B(new_n1186), .C1(G77), .C2(new_n741), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G116), .A2(new_n736), .B1(new_n744), .B2(G303), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n730), .A2(G107), .B1(new_n747), .B2(G294), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1187), .A2(new_n1004), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n735), .A2(new_n1106), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G132), .B2(new_n747), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n730), .A2(G150), .B1(new_n749), .B2(G159), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n725), .A2(new_n816), .B1(new_n743), .B2(new_n1110), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G50), .B2(new_n752), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1168), .A2(new_n1192), .A3(new_n1193), .A4(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1190), .B1(new_n1196), .B2(new_n774), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1185), .B1(new_n1197), .B2(new_n723), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1183), .B1(new_n1184), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1057), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n941), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n1202), .A3(new_n1078), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1199), .A2(new_n1203), .ZN(G381));
  OAI21_X1  g1004(.A(KEYINPUT122), .B1(new_n1096), .B2(new_n1123), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1077), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT114), .B1(new_n1094), .B2(new_n1078), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1083), .B(new_n1058), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT122), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1123), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1205), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(G375), .ZN(new_n1214));
  INV_X1    g1014(.A(G390), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n962), .A2(new_n1215), .A3(new_n985), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(G393), .A2(G396), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(G381), .A2(new_n1218), .A3(G384), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1213), .A2(new_n1214), .A3(new_n1217), .A4(new_n1219), .ZN(G407));
  INV_X1    g1020(.A(G213), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(G343), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1213), .A2(new_n1214), .A3(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(G407), .A2(new_n1223), .A3(G213), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT123), .ZN(G409));
  NAND2_X1  g1025(.A1(G393), .A2(G396), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1218), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1215), .B1(new_n962), .B2(new_n985), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1228), .B1(new_n1217), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G387), .A2(G390), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(new_n1216), .A3(new_n1227), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1126), .A2(new_n1141), .A3(new_n1202), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1234), .A2(new_n1148), .A3(new_n1177), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1205), .A2(new_n1212), .A3(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1145), .B(new_n1180), .C1(new_n1096), .C2(new_n1123), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT62), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1222), .ZN(new_n1240));
  OAI211_X1 g1040(.A(KEYINPUT124), .B(new_n1078), .C1(new_n1200), .C2(KEYINPUT60), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1019), .C1(new_n1242), .C2(new_n1201), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1201), .A2(new_n1242), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT124), .B1(new_n1244), .B2(new_n1078), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1199), .B1(new_n1243), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n825), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G384), .B(new_n1199), .C1(new_n1243), .C2(new_n1245), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .A4(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1222), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1222), .A2(G2897), .ZN(new_n1254));
  AND3_X1   g1054(.A1(new_n1247), .A2(new_n1248), .A3(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1254), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1251), .B(new_n1252), .C1(new_n1253), .C2(new_n1257), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1222), .B(new_n1249), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1259), .A2(new_n1239), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1233), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1253), .A2(KEYINPUT125), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1257), .B1(new_n1253), .B2(KEYINPUT125), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1230), .A2(new_n1252), .A3(new_n1232), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1259), .B2(KEYINPUT63), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1253), .A2(new_n1250), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT63), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1264), .A2(new_n1266), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1261), .A2(new_n1270), .ZN(G405));
  NAND3_X1  g1071(.A1(G375), .A2(new_n1205), .A3(new_n1212), .ZN(new_n1272));
  OR2_X1    g1072(.A1(new_n1272), .A2(KEYINPUT126), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1237), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1272), .B1(new_n1274), .B2(KEYINPUT126), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1273), .A2(new_n1275), .A3(new_n1233), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1233), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n1276), .A2(new_n1277), .B1(KEYINPUT127), .B2(new_n1249), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1233), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1249), .A2(KEYINPUT127), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1273), .A2(new_n1275), .A3(new_n1233), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1278), .A2(new_n1284), .ZN(G402));
endmodule


