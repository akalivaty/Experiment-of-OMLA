//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1155;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT67), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G235), .A3(G237), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT69), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n460), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n465), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT3), .B(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(new_n460), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n472), .A2(new_n478), .ZN(G160));
  NOR2_X1   g054(.A1(new_n461), .A2(new_n462), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n460), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  INV_X1    g059(.A(G100), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n485), .A2(new_n460), .A3(KEYINPUT70), .ZN(new_n486));
  AOI21_X1  g061(.A(KEYINPUT70), .B1(new_n485), .B2(new_n460), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G112), .B2(new_n460), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n482), .A2(new_n484), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(KEYINPUT4), .B(G138), .C1(new_n461), .C2(new_n462), .ZN(new_n491));
  NAND2_X1  g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(G114), .A2(G2104), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n475), .B2(G126), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n496), .B2(new_n460), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n463), .A2(new_n469), .A3(G138), .A4(new_n460), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(G164));
  AND2_X1   g074(.A1(KEYINPUT72), .A2(KEYINPUT6), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT72), .A2(KEYINPUT6), .ZN(new_n501));
  OAI21_X1  g076(.A(G651), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n502), .B(KEYINPUT73), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT6), .ZN(new_n505));
  XNOR2_X1  g080(.A(new_n505), .B(KEYINPUT71), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G88), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n503), .A2(G543), .A3(new_n506), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G50), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n517), .A2(new_n504), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n513), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n513), .A2(new_n516), .A3(new_n521), .A4(new_n518), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(G166));
  NAND2_X1  g098(.A1(new_n512), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT77), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT75), .B(G51), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n503), .A2(G543), .A3(new_n506), .A4(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT76), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n530), .A2(KEYINPUT76), .A3(new_n531), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n528), .A2(KEYINPUT78), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT78), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n524), .A2(new_n534), .A3(new_n527), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n537), .B2(new_n532), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n535), .A2(new_n538), .ZN(G168));
  NAND2_X1  g114(.A1(new_n512), .A2(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n515), .A2(G52), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n504), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(new_n512), .A2(G81), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n515), .A2(G43), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n504), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT79), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n553), .A2(new_n557), .ZN(G188));
  NAND4_X1  g133(.A1(new_n503), .A2(G91), .A3(new_n506), .A4(new_n510), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(new_n504), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n503), .A2(G53), .A3(G543), .A4(new_n506), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n562), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  AND2_X1   g142(.A1(new_n535), .A2(new_n538), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  OR2_X1    g144(.A1(new_n510), .A2(G74), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n515), .A2(G49), .B1(G651), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n512), .A2(G87), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G288));
  INV_X1    g148(.A(G48), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n514), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT80), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n511), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n512), .A2(G86), .B1(G651), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n576), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n581), .B1(new_n576), .B2(new_n580), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n512), .A2(G85), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n515), .A2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OR2_X1    g163(.A1(new_n588), .A2(new_n504), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(G290));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  NOR2_X1   g166(.A1(G301), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n512), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n512), .A2(KEYINPUT10), .A3(G92), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n504), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n515), .B2(G54), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n592), .B1(new_n602), .B2(new_n591), .ZN(G284));
  AOI21_X1  g178(.A(new_n592), .B1(new_n602), .B2(new_n591), .ZN(G321));
  NAND2_X1  g179(.A1(G299), .A2(new_n591), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G168), .B2(new_n591), .ZN(G280));
  XNOR2_X1  g181(.A(G280), .B(KEYINPUT82), .ZN(G297));
  INV_X1    g182(.A(G860), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n601), .B1(G559), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT83), .ZN(G148));
  NOR2_X1   g185(.A1(new_n550), .A2(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n601), .A2(G559), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n463), .A2(new_n469), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n473), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT12), .Z(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT13), .Z(new_n619));
  INV_X1    g194(.A(G2100), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  MUX2_X1   g197(.A(G99), .B(G111), .S(G2105), .Z(new_n623));
  AOI22_X1  g198(.A1(new_n483), .A2(G123), .B1(G2104), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G135), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n476), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT84), .B(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n621), .A2(new_n622), .A3(new_n628), .ZN(G156));
  INV_X1    g204(.A(G14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2451), .B(G2454), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT85), .B(KEYINPUT16), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT15), .B(G2435), .Z(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT86), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2430), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n630), .B1(new_n637), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n637), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT87), .ZN(G401));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT89), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT88), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2084), .B(G2090), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n650), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  INV_X1    g230(.A(new_n653), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n650), .B2(new_n652), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT90), .B(KEYINPUT17), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n650), .B(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n657), .B1(new_n659), .B2(new_n652), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n652), .A3(new_n656), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n655), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2096), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n620), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n666), .A2(new_n669), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT20), .Z(new_n673));
  AOI211_X1 g248(.A(new_n671), .B(new_n673), .C1(new_n666), .C2(new_n670), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT91), .ZN(new_n678));
  XOR2_X1   g253(.A(G1991), .B(G1996), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n676), .B(new_n680), .ZN(G229));
  OR2_X1    g256(.A1(G6), .A2(G16), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(G305), .B2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT32), .B(G1981), .Z(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(G22), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G166), .B2(new_n683), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1971), .ZN(new_n691));
  MUX2_X1   g266(.A(G23), .B(G288), .S(G16), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT33), .B(G1976), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n687), .A2(new_n688), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(G25), .A2(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n483), .A2(G119), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT92), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G95), .B(G107), .S(G2105), .Z(new_n701));
  AOI22_X1  g276(.A1(new_n481), .A2(G131), .B1(G2104), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT93), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n697), .B1(new_n705), .B2(G29), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n683), .A2(G24), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT94), .Z(new_n710));
  INV_X1    g285(.A(G290), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n683), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n708), .B1(G1986), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G1986), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n696), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n688), .B1(new_n687), .B2(new_n695), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT36), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n481), .A2(G139), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n473), .A2(G103), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(KEYINPUT25), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(KEYINPUT25), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n719), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT95), .ZN(new_n724));
  NAND2_X1  g299(.A1(G115), .A2(G2104), .ZN(new_n725));
  INV_X1    g300(.A(G127), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n615), .B2(new_n726), .ZN(new_n727));
  AND3_X1   g302(.A1(new_n727), .A2(KEYINPUT96), .A3(G2105), .ZN(new_n728));
  AOI21_X1  g303(.A(KEYINPUT96), .B1(new_n727), .B2(G2105), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n724), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  MUX2_X1   g305(.A(G33), .B(new_n730), .S(G29), .Z(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(G2072), .Z(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G26), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT28), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n481), .A2(G140), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n483), .A2(G128), .ZN(new_n737));
  MUX2_X1   g312(.A(G104), .B(G116), .S(G2105), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G2104), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n735), .B1(new_n741), .B2(new_n733), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2067), .ZN(new_n743));
  NOR2_X1   g318(.A1(G29), .A2(G35), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G162), .B2(G29), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT29), .Z(new_n746));
  INV_X1    g321(.A(G2090), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n481), .A2(G141), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT97), .Z(new_n750));
  AND2_X1   g325(.A1(new_n473), .A2(G105), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT26), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n751), .B(new_n753), .C1(G129), .C2(new_n483), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(new_n733), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n733), .B2(G32), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n743), .B(new_n748), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G27), .A2(G29), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G164), .B2(G29), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n746), .A2(new_n747), .B1(G2078), .B2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(new_n762), .ZN(new_n764));
  INV_X1    g339(.A(G2078), .ZN(new_n765));
  OR2_X1    g340(.A1(KEYINPUT24), .A2(G34), .ZN(new_n766));
  NAND2_X1  g341(.A1(KEYINPUT24), .A2(G34), .ZN(new_n767));
  AOI21_X1  g342(.A(G29), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G160), .B2(G29), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n764), .A2(new_n765), .B1(G2084), .B2(new_n769), .ZN(new_n770));
  AND4_X1   g345(.A1(new_n732), .A2(new_n760), .A3(new_n763), .A4(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G4), .A2(G16), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n602), .B2(G16), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1348), .ZN(new_n774));
  NOR2_X1   g349(.A1(G16), .A2(G19), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n551), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1341), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  OAI22_X1  g353(.A1(new_n758), .A2(new_n759), .B1(G2084), .B2(new_n769), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n683), .A2(G5), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G171), .B2(new_n683), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G1961), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(KEYINPUT100), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n683), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT23), .Z(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G299), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G1956), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n783), .B2(KEYINPUT100), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n771), .A2(new_n778), .A3(new_n784), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G286), .A2(new_n683), .ZN(new_n792));
  OR2_X1    g367(.A1(G16), .A2(G21), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n792), .B1(KEYINPUT98), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(KEYINPUT98), .B2(new_n792), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(G1966), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(G1966), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT31), .B(G11), .Z(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT30), .B(G28), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n798), .B1(new_n733), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n626), .B2(new_n733), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n781), .B2(G1961), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n796), .A2(new_n797), .A3(new_n802), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(KEYINPUT99), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(KEYINPUT99), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n791), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n718), .A2(new_n806), .ZN(G311));
  NAND2_X1  g382(.A1(new_n718), .A2(new_n806), .ZN(G150));
  NAND2_X1  g383(.A1(new_n602), .A2(G559), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT38), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n515), .A2(G55), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n512), .A2(G93), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n811), .B(new_n812), .C1(new_n504), .C2(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(KEYINPUT101), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(KEYINPUT101), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n815), .A2(new_n550), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n551), .A2(new_n814), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n810), .B(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n822), .A2(new_n608), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n815), .A2(new_n816), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(G145));
  XNOR2_X1  g403(.A(new_n730), .B(new_n756), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n703), .B(KEYINPUT93), .ZN(new_n830));
  INV_X1    g405(.A(new_n618), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n705), .A2(new_n618), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n481), .A2(G142), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n483), .A2(G130), .ZN(new_n835));
  MUX2_X1   g410(.A(G106), .B(G118), .S(G2105), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G2104), .ZN(new_n837));
  AND3_X1   g412(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n832), .A2(new_n833), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n839), .B1(new_n832), .B2(new_n833), .ZN(new_n842));
  XNOR2_X1  g417(.A(G164), .B(new_n740), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n841), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n832), .A2(new_n833), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n838), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n843), .B1(new_n847), .B2(new_n840), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n829), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(G160), .B(new_n489), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n626), .Z(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n844), .B1(new_n841), .B2(new_n842), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n847), .A2(new_n840), .A3(new_n843), .ZN(new_n854));
  INV_X1    g429(.A(new_n829), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n849), .A2(new_n852), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT102), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n849), .A2(new_n859), .A3(new_n852), .A4(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n849), .A2(new_n856), .ZN(new_n862));
  AOI21_X1  g437(.A(G37), .B1(new_n862), .B2(new_n851), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g440(.A(new_n584), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(G303), .A3(new_n582), .ZN(new_n867));
  OAI21_X1  g442(.A(G166), .B1(new_n583), .B2(new_n584), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(G288), .B(G290), .Z(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(KEYINPUT103), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(new_n874), .A3(new_n871), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(new_n869), .B2(new_n871), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n867), .A2(new_n868), .A3(KEYINPUT104), .A4(new_n870), .ZN(new_n878));
  AOI22_X1  g453(.A1(new_n873), .A2(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n879), .A2(KEYINPUT42), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n819), .B(new_n612), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n602), .A2(new_n566), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n601), .A2(G299), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(KEYINPUT41), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(new_n887), .A3(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n885), .B1(new_n881), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n879), .A2(KEYINPUT42), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n880), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n890), .B1(new_n880), .B2(new_n891), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI211_X1 g470(.A(KEYINPUT105), .B(new_n890), .C1(new_n880), .C2(new_n891), .ZN(new_n896));
  OAI21_X1  g471(.A(G868), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n825), .A2(new_n591), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(G295));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n898), .ZN(G331));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n877), .A2(new_n878), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n874), .B1(new_n869), .B2(new_n871), .ZN(new_n903));
  INV_X1    g478(.A(new_n875), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n884), .A2(KEYINPUT106), .A3(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(G286), .A2(G301), .ZN(new_n907));
  NAND2_X1  g482(.A1(G168), .A2(G171), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n819), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n819), .B1(new_n907), .B2(new_n908), .ZN(new_n911));
  OAI221_X1 g486(.A(new_n906), .B1(new_n889), .B2(KEYINPUT106), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n908), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n820), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n914), .A2(new_n883), .A3(new_n882), .A4(new_n909), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n905), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n889), .B1(new_n910), .B2(new_n911), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n915), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n917), .B1(new_n919), .B2(new_n879), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n901), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n905), .A2(new_n915), .A3(new_n918), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n879), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT43), .A4(new_n917), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT44), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT43), .B1(new_n916), .B2(new_n920), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n922), .A2(new_n923), .A3(new_n917), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n926), .B1(KEYINPUT43), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n925), .B1(KEYINPUT44), .B2(new_n928), .ZN(G397));
  NOR2_X1   g504(.A1(G290), .A2(G1986), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(G164), .B2(G1384), .ZN(new_n932));
  INV_X1    g507(.A(new_n478), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n470), .A2(new_n471), .ZN(new_n934));
  OAI211_X1 g509(.A(G40), .B(new_n933), .C1(new_n934), .C2(new_n460), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n930), .A2(KEYINPUT48), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT48), .ZN(new_n938));
  INV_X1    g513(.A(new_n930), .ZN(new_n939));
  INV_X1    g514(.A(new_n936), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AND2_X1   g516(.A1(new_n755), .A2(G1996), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n755), .A2(G1996), .ZN(new_n943));
  INV_X1    g518(.A(G2067), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n740), .B(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n942), .A2(new_n943), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n705), .A2(new_n707), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n705), .A2(new_n707), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n937), .B(new_n941), .C1(new_n951), .C2(new_n940), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n949), .B1(new_n947), .B2(new_n940), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(G2067), .B2(new_n740), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n954), .A2(KEYINPUT126), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n936), .B1(new_n954), .B2(KEYINPUT126), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n940), .B1(new_n756), .B2(new_n945), .ZN(new_n958));
  OR3_X1    g533(.A1(new_n940), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT46), .B1(new_n940), .B2(G1996), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT47), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n957), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G40), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n472), .A2(new_n964), .A3(new_n478), .ZN(new_n965));
  OAI21_X1  g540(.A(G126), .B1(new_n461), .B2(new_n462), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n460), .B1(new_n966), .B2(new_n494), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT4), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n498), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n493), .ZN(new_n970));
  AOI21_X1  g545(.A(G1384), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n965), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(G8), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT109), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1976), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n571), .A2(new_n976), .A3(new_n572), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT49), .ZN(new_n978));
  INV_X1    g553(.A(G1981), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n576), .A2(new_n580), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n979), .B1(new_n576), .B2(new_n580), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n982), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n984), .A2(KEYINPUT49), .A3(new_n980), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n983), .A2(new_n985), .A3(new_n975), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n983), .A2(new_n985), .A3(KEYINPUT113), .A4(new_n975), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n977), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n980), .B(KEYINPUT114), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n975), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n989), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n571), .A2(G1976), .A3(new_n572), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n995), .A2(KEYINPUT110), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n995), .A2(KEYINPUT110), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n974), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n994), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n996), .A2(new_n997), .ZN(new_n1001));
  OAI211_X1 g576(.A(KEYINPUT111), .B(KEYINPUT52), .C1(new_n1001), .C2(new_n974), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT52), .B1(G288), .B2(new_n976), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n1003), .B(KEYINPUT112), .Z(new_n1004));
  AOI22_X1  g579(.A1(new_n1000), .A2(new_n1002), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G303), .A2(G8), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n971), .A2(KEYINPUT45), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n932), .A2(new_n1009), .A3(new_n965), .ZN(new_n1010));
  INV_X1    g585(.A(G1971), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1010), .A2(KEYINPUT107), .A3(new_n1011), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n969), .A2(new_n970), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n965), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n971), .A2(KEYINPUT108), .A3(new_n1017), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT108), .B1(new_n971), .B2(new_n1017), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1014), .B(new_n1015), .C1(new_n1024), .C2(G2090), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1025), .A2(G8), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n993), .A2(new_n1005), .A3(new_n1008), .A4(new_n1026), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n992), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1006), .B(KEYINPUT55), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n935), .B1(new_n1017), .B2(new_n971), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(new_n1017), .B2(new_n971), .ZN(new_n1031));
  XNOR2_X1  g606(.A(new_n1031), .B(KEYINPUT115), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1012), .B1(new_n1032), .B2(G2090), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(G8), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1029), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1008), .A2(G8), .A3(new_n1025), .ZN(new_n1036));
  AND4_X1   g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n993), .A4(new_n1005), .ZN(new_n1037));
  INV_X1    g612(.A(G1966), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n965), .B(KEYINPUT116), .C1(new_n971), .C2(KEYINPUT45), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n1009), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT116), .B1(new_n932), .B2(new_n965), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1038), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT117), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1044), .B(new_n1038), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G2084), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT108), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n1048), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1030), .A2(new_n1047), .A3(new_n1023), .A4(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1050), .B(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1046), .A2(G168), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(G8), .A3(G168), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT63), .B1(new_n1037), .B2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1036), .A2(new_n993), .A3(KEYINPUT63), .A4(new_n1005), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1026), .A2(KEYINPUT119), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1026), .A2(KEYINPUT119), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1008), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1057), .A2(new_n1054), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1028), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1010), .B2(G2078), .ZN(new_n1064));
  XOR2_X1   g639(.A(new_n1064), .B(KEYINPUT125), .Z(new_n1065));
  INV_X1    g640(.A(G1961), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1024), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n965), .B1(new_n971), .B2(KEYINPUT45), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(new_n1009), .A3(new_n1039), .ZN(new_n1071));
  OR3_X1    g646(.A1(new_n1071), .A2(new_n1063), .A3(G2078), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1065), .A2(new_n1067), .A3(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1073), .A2(G301), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1045), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1044), .B1(new_n1071), .B2(new_n1038), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1022), .A2(new_n1051), .A3(new_n1047), .A4(new_n1023), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1050), .A2(KEYINPUT118), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(G286), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(KEYINPUT51), .A3(G8), .A4(new_n1053), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1053), .A2(G8), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT51), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1082), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1087), .A2(new_n1088), .A3(KEYINPUT62), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT62), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1080), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT51), .B1(new_n1091), .B2(G168), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(new_n1083), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT51), .B1(new_n1053), .B2(G8), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT124), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1082), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1090), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1074), .B1(new_n1089), .B2(new_n1097), .ZN(new_n1098));
  XOR2_X1   g673(.A(G301), .B(KEYINPUT54), .Z(new_n1099));
  INV_X1    g674(.A(new_n1010), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(KEYINPUT53), .A3(new_n765), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1065), .A2(new_n1067), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1073), .B2(new_n1099), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n1104));
  NAND3_X1  g679(.A1(G299), .A2(new_n1104), .A3(KEYINPUT57), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n566), .B2(KEYINPUT120), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1031), .A2(new_n788), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT56), .B(G2072), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1100), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n972), .A2(G2067), .ZN(new_n1114));
  INV_X1    g689(.A(G1348), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1114), .B1(new_n1024), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1113), .B1(new_n601), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1105), .A2(new_n1107), .A3(new_n1109), .A4(new_n1111), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1119), .B(new_n1120), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1113), .A2(KEYINPUT61), .A3(new_n1118), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1116), .A2(new_n1123), .A3(new_n602), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT58), .B(G1341), .Z(new_n1125));
  NAND2_X1  g700(.A1(new_n972), .A2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1010), .B2(G1996), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1127), .A2(new_n551), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT59), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1124), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1122), .A2(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1116), .A2(new_n601), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1116), .A2(new_n601), .ZN(new_n1136));
  OAI21_X1  g711(.A(KEYINPUT60), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT61), .B1(new_n1113), .B2(new_n1118), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g715(.A(KEYINPUT123), .B(KEYINPUT61), .C1(new_n1113), .C2(new_n1118), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1134), .B(new_n1137), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1103), .B1(new_n1121), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1098), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1062), .B1(new_n1145), .B2(new_n1037), .ZN(new_n1146));
  XOR2_X1   g721(.A(G290), .B(G1986), .Z(new_n1147));
  AOI21_X1  g722(.A(new_n940), .B1(new_n951), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n963), .B1(new_n1146), .B2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g724(.A1(new_n647), .A2(G319), .ZN(new_n1151));
  OR3_X1    g725(.A1(G229), .A2(G227), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g726(.A(new_n1152), .B1(new_n861), .B2(new_n863), .ZN(new_n1153));
  NAND3_X1  g727(.A1(new_n921), .A2(new_n1153), .A3(new_n924), .ZN(G225));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n1155));
  XNOR2_X1  g729(.A(G225), .B(new_n1155), .ZN(G308));
endmodule


