//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071;
  XNOR2_X1  g000(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT69), .A2(G237), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT69), .A2(G237), .ZN(new_n189));
  AOI21_X1  g003(.A(G953), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  AOI21_X1  g006(.A(G143), .B1(new_n190), .B2(G214), .ZN(new_n193));
  OAI21_X1  g007(.A(G131), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT17), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n188), .A2(new_n189), .ZN(new_n196));
  INV_X1    g010(.A(G953), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(G214), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G143), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(new_n191), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n194), .A2(new_n195), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(G140), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G125), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G125), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G140), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n206), .B1(new_n210), .B2(new_n204), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g027(.A(G146), .B(new_n206), .C1(new_n210), .C2(new_n204), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n201), .B1(new_n200), .B2(new_n191), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(KEYINPUT17), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n203), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT18), .A2(G131), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n219), .B1(new_n200), .B2(new_n191), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n210), .A2(G146), .ZN(new_n222));
  XNOR2_X1  g036(.A(G125), .B(G140), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(new_n212), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n200), .A2(new_n191), .A3(new_n219), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n221), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(KEYINPUT84), .B(G104), .Z(new_n228));
  XNOR2_X1  g042(.A(G113), .B(G122), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n218), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(new_n225), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(new_n220), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT19), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n223), .B(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n214), .B1(new_n236), .B2(G146), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(new_n194), .B2(new_n202), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n230), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n232), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(G475), .A2(G902), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n187), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n241), .ZN(new_n243));
  AOI211_X1 g057(.A(KEYINPUT20), .B(new_n243), .C1(new_n232), .C2(new_n239), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n218), .A2(new_n227), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n230), .ZN(new_n246));
  AOI21_X1  g060(.A(G902), .B1(new_n246), .B2(new_n232), .ZN(new_n247));
  INV_X1    g061(.A(G475), .ZN(new_n248));
  OAI22_X1  g062(.A1(new_n242), .A2(new_n244), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(G143), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n199), .A2(G128), .ZN(new_n252));
  OR3_X1    g066(.A1(new_n251), .A2(new_n252), .A3(G134), .ZN(new_n253));
  OAI21_X1  g067(.A(G134), .B1(new_n251), .B2(new_n252), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT85), .ZN(new_n256));
  INV_X1    g070(.A(G116), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(G122), .ZN(new_n258));
  INV_X1    g072(.A(G122), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT85), .A3(G116), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n257), .A2(G122), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT14), .ZN(new_n263));
  OR3_X1    g077(.A1(new_n259), .A2(KEYINPUT14), .A3(G116), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G107), .ZN(new_n266));
  INV_X1    g080(.A(G107), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n261), .A2(new_n267), .A3(new_n262), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n255), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n199), .A2(G128), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT13), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n252), .B2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n273), .A2(KEYINPUT86), .B1(KEYINPUT13), .B2(new_n251), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT86), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n275), .B(new_n271), .C1(new_n252), .C2(new_n272), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n270), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n261), .A2(new_n267), .A3(new_n262), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n267), .B1(new_n261), .B2(new_n262), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n253), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n269), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT88), .ZN(new_n282));
  INV_X1    g096(.A(G234), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT9), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT9), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G234), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT78), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n287), .B1(new_n284), .B2(new_n286), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT87), .ZN(new_n291));
  INV_X1    g105(.A(G217), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(G953), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n291), .B1(new_n290), .B2(new_n293), .ZN(new_n295));
  OR2_X1    g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT88), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n269), .B(new_n297), .C1(new_n277), .C2(new_n280), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n282), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G902), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n273), .A2(KEYINPUT86), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n251), .A2(KEYINPUT13), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n276), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G134), .ZN(new_n304));
  INV_X1    g118(.A(new_n279), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n268), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n306), .A3(new_n253), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n294), .A2(new_n295), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n307), .A2(new_n308), .A3(new_n297), .A4(new_n269), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n299), .A2(new_n300), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G478), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(KEYINPUT15), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n310), .B(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n197), .A2(G952), .ZN(new_n314));
  NAND2_X1  g128(.A1(G234), .A2(G237), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(G902), .A3(G953), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT21), .B(G898), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n317), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n249), .A2(new_n313), .A3(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(KEYINPUT67), .B(G119), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(G128), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n250), .A2(G119), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n323), .A2(G128), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT76), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n323), .A2(G128), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n327), .A2(new_n324), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT76), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(new_n325), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT24), .B(G110), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n250), .A2(KEYINPUT23), .A3(G119), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n323), .A2(G128), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n330), .B(new_n339), .C1(new_n340), .C2(KEYINPUT23), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G110), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n338), .A2(new_n215), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT22), .B(G137), .ZN(new_n344));
  INV_X1    g158(.A(G221), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n345), .A2(new_n283), .A3(G953), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n344), .B(new_n346), .Z(new_n347));
  NAND3_X1  g161(.A1(new_n329), .A2(new_n334), .A3(new_n336), .ZN(new_n348));
  OR2_X1    g162(.A1(new_n341), .A2(G110), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT77), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT77), .B1(new_n348), .B2(new_n349), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n214), .A2(new_n224), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n343), .B(new_n347), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n347), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n348), .A2(new_n349), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n354), .B1(new_n360), .B2(new_n350), .ZN(new_n361));
  INV_X1    g175(.A(new_n343), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n356), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n292), .B1(G234), .B2(new_n300), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(G902), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n366), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n355), .A2(new_n363), .A3(new_n300), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT25), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n355), .A2(new_n363), .A3(KEYINPUT25), .A4(new_n300), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n370), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n369), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G214), .B1(G237), .B2(G902), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G104), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT3), .B1(new_n380), .B2(G107), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n267), .A3(G104), .ZN(new_n383));
  INV_X1    g197(.A(G101), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n380), .A2(G107), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n381), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n380), .A2(G107), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n267), .A2(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n323), .A2(G116), .ZN(new_n391));
  INV_X1    g205(.A(G119), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(G116), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  XOR2_X1   g208(.A(KEYINPUT2), .B(G113), .Z(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT68), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n393), .B1(new_n323), .B2(G116), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT68), .A3(new_n395), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n390), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(KEYINPUT5), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n402), .B(G113), .C1(KEYINPUT5), .C2(new_n391), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G101), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT4), .A3(new_n386), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n408), .A3(G101), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n399), .A2(new_n395), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n398), .B2(new_n400), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n404), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G122), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n404), .B(new_n414), .C1(new_n412), .C2(new_n410), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(KEYINPUT6), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n412), .ZN(new_n419));
  INV_X1    g233(.A(new_n410), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n419), .A2(new_n420), .B1(new_n403), .B2(new_n401), .ZN(new_n421));
  OR3_X1    g235(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n414), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n212), .A2(G143), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n199), .A2(G146), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT1), .B1(new_n199), .B2(G146), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(G128), .A3(new_n426), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n423), .B(new_n424), .C1(KEYINPUT1), .C2(new_n250), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n208), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n423), .A2(new_n424), .A3(KEYINPUT0), .A4(G128), .ZN(new_n430));
  XNOR2_X1  g244(.A(G143), .B(G146), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT0), .B(G128), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n429), .B1(new_n433), .B2(new_n208), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n197), .A2(G224), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n434), .B(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n418), .A2(new_n422), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(KEYINPUT7), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT82), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n434), .A2(new_n439), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n438), .A2(KEYINPUT82), .ZN(new_n441));
  MUX2_X1   g255(.A(new_n434), .B(new_n440), .S(new_n441), .Z(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(new_n421), .B2(new_n414), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n414), .B(KEYINPUT8), .ZN(new_n444));
  OAI21_X1  g258(.A(G113), .B1(new_n391), .B2(KEYINPUT5), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n445), .B1(new_n402), .B2(KEYINPUT81), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(KEYINPUT81), .B2(new_n402), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n447), .A2(new_n401), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n386), .A2(new_n389), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n398), .A2(new_n400), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n449), .B1(new_n450), .B2(new_n403), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n444), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(G902), .B1(new_n443), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n437), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G210), .B1(G237), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n437), .A2(new_n453), .A3(new_n455), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n379), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n345), .B1(new_n290), .B2(new_n300), .ZN(new_n460));
  XOR2_X1   g274(.A(G110), .B(G140), .Z(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT79), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n197), .A2(G227), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n427), .A2(new_n428), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n390), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n427), .A2(new_n386), .A3(new_n389), .A4(new_n428), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G137), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(KEYINPUT11), .A3(G134), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n270), .A2(G137), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT11), .ZN(new_n473));
  OAI211_X1 g287(.A(KEYINPUT64), .B(new_n473), .C1(new_n270), .C2(G137), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n469), .A2(G134), .ZN(new_n476));
  AOI21_X1  g290(.A(KEYINPUT64), .B1(new_n476), .B2(new_n473), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n472), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G131), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n472), .B(new_n201), .C1(new_n475), .C2(new_n477), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n468), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT12), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n468), .A2(new_n481), .A3(KEYINPUT12), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n467), .B(KEYINPUT10), .ZN(new_n487));
  INV_X1    g301(.A(new_n433), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n407), .A2(new_n488), .A3(new_n409), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n470), .A2(new_n471), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n473), .B1(new_n270), .B2(G137), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT64), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI211_X1 g307(.A(G131), .B(new_n490), .C1(new_n493), .C2(new_n474), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n474), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n201), .B1(new_n495), .B2(new_n472), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT80), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT80), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n479), .A2(new_n498), .A3(new_n480), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n487), .A2(new_n489), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n464), .B1(new_n486), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n427), .A2(new_n428), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(KEYINPUT10), .A3(new_n449), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT10), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n467), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n489), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n481), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n500), .A2(new_n507), .A3(new_n464), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(G469), .B1(new_n509), .B2(G902), .ZN(new_n510));
  INV_X1    g324(.A(new_n464), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n506), .A2(new_n481), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n497), .A2(new_n499), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(new_n506), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n511), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n486), .A2(new_n500), .A3(new_n464), .ZN(new_n516));
  AOI21_X1  g330(.A(G902), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(G469), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n460), .B1(new_n510), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n459), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n377), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT74), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n476), .A2(new_n471), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G131), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n480), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT66), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT66), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n480), .A2(new_n528), .A3(new_n525), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n502), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n488), .B1(new_n494), .B2(new_n496), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT65), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n481), .A2(KEYINPUT65), .A3(new_n488), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n502), .A2(new_n480), .A3(new_n525), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n531), .A2(KEYINPUT30), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n419), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n190), .A2(G210), .ZN(new_n541));
  XOR2_X1   g355(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT26), .B(G101), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n412), .A2(new_n531), .A3(new_n538), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n540), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT31), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n539), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n535), .B2(new_n536), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n547), .B1(new_n553), .B2(new_n419), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(KEYINPUT31), .A3(new_n546), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT72), .ZN(new_n556));
  XOR2_X1   g370(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT65), .B1(new_n481), .B2(new_n488), .ZN(new_n559));
  AOI211_X1 g373(.A(new_n532), .B(new_n433), .C1(new_n479), .C2(new_n480), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n412), .B1(new_n561), .B2(new_n530), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n556), .B(new_n558), .C1(new_n562), .C2(new_n547), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n547), .B1(new_n535), .B2(new_n419), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT72), .B1(new_n564), .B2(new_n557), .ZN(new_n565));
  OR2_X1    g379(.A1(new_n547), .A2(KEYINPUT28), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI22_X1  g381(.A1(new_n551), .A2(new_n555), .B1(new_n567), .B2(new_n545), .ZN(new_n568));
  NOR2_X1   g382(.A1(G472), .A2(G902), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT32), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT32), .ZN(new_n572));
  AND4_X1   g386(.A1(KEYINPUT31), .A2(new_n540), .A3(new_n546), .A4(new_n548), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT31), .B1(new_n554), .B2(new_n546), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n566), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n564), .A2(new_n557), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(new_n556), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n546), .B1(new_n578), .B2(new_n565), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n572), .B(new_n569), .C1(new_n575), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n571), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G472), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n540), .A2(new_n548), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT29), .B1(new_n583), .B2(new_n545), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n563), .A2(new_n565), .A3(new_n546), .A4(new_n566), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n412), .B1(new_n538), .B2(new_n531), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT28), .B1(new_n547), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT29), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n545), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n566), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n591), .A2(KEYINPUT73), .A3(new_n300), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT73), .B1(new_n591), .B2(new_n300), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n582), .B1(new_n586), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n523), .B1(new_n581), .B2(new_n596), .ZN(new_n597));
  AOI211_X1 g411(.A(KEYINPUT74), .B(new_n595), .C1(new_n571), .C2(new_n580), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n322), .B(new_n522), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  NAND2_X1  g414(.A1(new_n551), .A2(new_n555), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n567), .A2(new_n545), .ZN(new_n602));
  AOI21_X1  g416(.A(G902), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI22_X1  g417(.A1(new_n603), .A2(new_n582), .B1(new_n568), .B2(new_n570), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT92), .ZN(new_n606));
  INV_X1    g420(.A(new_n321), .ZN(new_n607));
  INV_X1    g421(.A(new_n458), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n455), .B1(new_n437), .B2(new_n453), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n607), .B(new_n378), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n299), .A2(new_n611), .A3(new_n309), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n269), .B(KEYINPUT89), .C1(new_n277), .C2(new_n280), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT90), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n296), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n614), .B1(new_n294), .B2(new_n295), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n616), .A2(KEYINPUT89), .B1(new_n307), .B2(new_n269), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT33), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n311), .A2(G902), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n612), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT91), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n310), .A2(new_n311), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n612), .A2(new_n618), .A3(KEYINPUT91), .A4(new_n619), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n249), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n606), .B1(new_n610), .B2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n610), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT92), .ZN(new_n629));
  INV_X1    g443(.A(new_n520), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n369), .A2(new_n630), .A3(new_n375), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n605), .A2(new_n627), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  INV_X1    g448(.A(new_n610), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n605), .A2(new_n635), .A3(new_n631), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n232), .A2(new_n239), .ZN(new_n637));
  INV_X1    g451(.A(new_n187), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n637), .A2(new_n638), .A3(new_n243), .ZN(new_n639));
  OAI22_X1  g453(.A1(new_n639), .A2(new_n242), .B1(new_n248), .B2(new_n247), .ZN(new_n640));
  INV_X1    g454(.A(new_n313), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT35), .B(G107), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NOR2_X1   g459(.A1(new_n361), .A2(new_n362), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n357), .A2(KEYINPUT36), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n648), .A2(new_n367), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n375), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n521), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n605), .A2(new_n652), .A3(new_n322), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT93), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT37), .B(G110), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  OR2_X1    g470(.A1(new_n318), .A2(G900), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n316), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n640), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n313), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n652), .B(new_n662), .C1(new_n597), .C2(new_n598), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  NOR2_X1   g478(.A1(new_n608), .A2(new_n609), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n665), .B(KEYINPUT38), .Z(new_n666));
  NOR2_X1   g480(.A1(new_n554), .A2(new_n545), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n547), .A2(new_n587), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n300), .B1(new_n668), .B2(new_n546), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT94), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n581), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n375), .A2(new_n650), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n249), .A2(new_n313), .A3(new_n378), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n666), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT95), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n666), .A2(new_n672), .A3(KEYINPUT95), .A4(new_n675), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n658), .B(KEYINPUT39), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n520), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n681), .B(KEYINPUT40), .Z(new_n682));
  AND3_X1   g496(.A1(new_n678), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n199), .ZN(G45));
  AND2_X1   g498(.A1(new_n620), .A2(new_n621), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n624), .A2(new_n623), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n249), .B(new_n658), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT96), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n625), .A2(KEYINPUT96), .A3(new_n249), .A4(new_n658), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n652), .B(new_n692), .C1(new_n597), .C2(new_n598), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G146), .ZN(G48));
  NAND2_X1  g508(.A1(new_n601), .A2(new_n602), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n572), .B1(new_n695), .B2(new_n569), .ZN(new_n696));
  AOI211_X1 g510(.A(KEYINPUT32), .B(new_n570), .C1(new_n601), .C2(new_n602), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n596), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT74), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n581), .A2(new_n523), .A3(new_n596), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n377), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(G469), .B1(new_n517), .B2(KEYINPUT97), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT97), .ZN(new_n703));
  AOI211_X1 g517(.A(new_n703), .B(G902), .C1(new_n515), .C2(new_n516), .ZN(new_n704));
  OAI211_X1 g518(.A(KEYINPUT98), .B(new_n519), .C1(new_n702), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n515), .A2(new_n516), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n300), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n703), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT98), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n517), .A2(KEYINPUT97), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n708), .A2(new_n709), .A3(G469), .A4(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n460), .B1(new_n705), .B2(new_n711), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n629), .A2(new_n627), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n701), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND2_X1  g530(.A1(new_n705), .A2(new_n711), .ZN(new_n717));
  INV_X1    g531(.A(new_n460), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n459), .A3(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n719), .A2(new_n321), .A3(new_n642), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n720), .B(new_n376), .C1(new_n597), .C2(new_n598), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT99), .B(G116), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G18));
  NOR2_X1   g537(.A1(new_n719), .A2(new_n651), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n322), .B(new_n724), .C1(new_n597), .C2(new_n598), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  AND4_X1   g540(.A1(new_n607), .A2(new_n717), .A3(new_n459), .A4(new_n718), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n638), .B1(new_n637), .B2(new_n243), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT20), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n240), .A2(new_n729), .A3(new_n241), .ZN(new_n730));
  INV_X1    g544(.A(new_n232), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n231), .B1(new_n218), .B2(new_n227), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n300), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n728), .A2(new_n730), .B1(G475), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n641), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n695), .A2(new_n300), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT100), .B(G472), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n566), .A2(new_n588), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n601), .B1(new_n546), .B2(new_n738), .ZN(new_n739));
  AOI22_X1  g553(.A1(new_n736), .A2(new_n737), .B1(new_n569), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n727), .A2(new_n376), .A3(new_n735), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  AND3_X1   g556(.A1(new_n689), .A2(KEYINPUT101), .A3(new_n690), .ZN(new_n743));
  AOI21_X1  g557(.A(KEYINPUT101), .B1(new_n689), .B2(new_n690), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n745), .A2(new_n724), .A3(new_n740), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G125), .ZN(G27));
  NOR3_X1   g561(.A1(new_n608), .A2(new_n609), .A3(new_n379), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(KEYINPUT42), .A3(new_n520), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n743), .A2(new_n744), .A3(new_n749), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT102), .B1(new_n696), .B2(new_n697), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT102), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n571), .A2(new_n752), .A3(new_n580), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n751), .A2(new_n596), .A3(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n750), .A2(new_n754), .A3(new_n376), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n699), .A2(new_n700), .ZN(new_n756));
  INV_X1    g570(.A(new_n748), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n757), .A2(new_n630), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n756), .A2(new_n376), .A3(new_n745), .A4(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT42), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n755), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n201), .ZN(G33));
  NAND3_X1  g576(.A1(new_n701), .A2(new_n662), .A3(new_n758), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  INV_X1    g578(.A(KEYINPUT43), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n625), .A2(new_n765), .A3(new_n734), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n765), .B1(new_n625), .B2(new_n734), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n604), .A2(new_n768), .A3(KEYINPUT44), .A4(new_n673), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT103), .ZN(new_n770));
  OAI21_X1  g584(.A(G472), .B1(new_n568), .B2(G902), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n695), .A2(new_n569), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n651), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT103), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n774), .A3(KEYINPUT44), .A4(new_n768), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n770), .A2(new_n775), .A3(new_n748), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT104), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT104), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n770), .A2(new_n775), .A3(new_n778), .A4(new_n748), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n604), .A2(new_n768), .A3(new_n673), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT105), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n780), .A2(KEYINPUT105), .A3(new_n781), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n777), .A2(KEYINPUT106), .A3(new_n779), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n788), .B1(new_n501), .B2(new_n508), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n500), .A2(new_n507), .A3(new_n464), .ZN(new_n790));
  INV_X1    g604(.A(new_n506), .ZN(new_n791));
  INV_X1    g605(.A(new_n513), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n791), .A2(new_n792), .B1(new_n484), .B2(new_n485), .ZN(new_n793));
  OAI211_X1 g607(.A(KEYINPUT45), .B(new_n790), .C1(new_n793), .C2(new_n464), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n794), .A3(G469), .ZN(new_n795));
  NAND2_X1  g609(.A1(G469), .A2(G902), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT46), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n796), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n519), .A3(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(new_n718), .A3(new_n680), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n787), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n776), .A2(KEYINPUT104), .B1(new_n784), .B2(new_n785), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT106), .B1(new_n803), .B2(new_n779), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n469), .ZN(G39));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  INV_X1    g621(.A(new_n799), .ZN(new_n808));
  INV_X1    g622(.A(new_n519), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n808), .A2(new_n797), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n807), .B1(new_n810), .B2(new_n460), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n800), .A2(KEYINPUT47), .A3(new_n718), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n691), .A2(new_n376), .A3(new_n757), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n699), .A3(new_n700), .A4(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(KEYINPUT107), .B(G140), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n815), .B(new_n816), .ZN(G42));
  NAND3_X1  g631(.A1(new_n376), .A2(new_n378), .A3(new_n718), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n665), .B(KEYINPUT38), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n734), .A3(new_n625), .ZN(new_n820));
  INV_X1    g634(.A(new_n717), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n818), .B(new_n820), .C1(KEYINPUT49), .C2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n672), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n821), .A2(KEYINPUT49), .ZN(new_n824));
  XOR2_X1   g638(.A(new_n824), .B(KEYINPUT108), .Z(new_n825));
  NAND3_X1  g639(.A1(new_n822), .A2(new_n823), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n641), .A2(new_n249), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n605), .A2(new_n635), .A3(new_n631), .A4(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n741), .A2(new_n828), .A3(new_n653), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n829), .B1(new_n701), .B2(new_n713), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n721), .A2(new_n725), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n605), .A2(new_n628), .A3(new_n631), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n599), .A2(KEYINPUT109), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(KEYINPUT109), .B1(new_n599), .B2(new_n832), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n830), .B(new_n831), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n665), .A2(new_n674), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n630), .A2(new_n659), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT110), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n837), .A2(new_n651), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n838), .B1(new_n837), .B2(new_n651), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n672), .B(new_n836), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n663), .A2(new_n693), .A3(new_n746), .A4(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n835), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n640), .A2(new_n313), .A3(new_n659), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n756), .A2(new_n846), .B1(new_n740), .B2(new_n745), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n758), .A2(new_n673), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n763), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n845), .A2(new_n849), .A3(new_n761), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT101), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n691), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n689), .A2(KEYINPUT101), .A3(new_n690), .ZN(new_n854));
  AND4_X1   g668(.A1(new_n724), .A2(new_n740), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n652), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n699), .B2(new_n700), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n855), .B1(new_n857), .B2(new_n662), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n851), .B1(new_n859), .B2(KEYINPUT52), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n844), .A2(new_n850), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n599), .A2(new_n832), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT109), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n599), .A2(KEYINPUT109), .A3(new_n832), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n741), .A2(new_n828), .A3(new_n653), .ZN(new_n867));
  AND4_X1   g681(.A1(new_n714), .A2(new_n867), .A3(new_n721), .A4(new_n725), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT52), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n858), .A2(new_n871), .A3(new_n693), .A4(new_n841), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n376), .B(new_n758), .C1(new_n597), .C2(new_n598), .ZN(new_n873));
  INV_X1    g687(.A(new_n745), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n760), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n755), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n873), .A2(new_n661), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n846), .B1(new_n597), .B2(new_n598), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n745), .A2(new_n740), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n848), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n872), .A2(new_n877), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n851), .B1(new_n870), .B2(new_n883), .ZN(new_n884));
  XOR2_X1   g698(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n885));
  NAND3_X1  g699(.A1(new_n861), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n851), .B1(new_n858), .B2(new_n871), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n844), .A2(new_n850), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n888), .B1(new_n890), .B2(new_n884), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT51), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n813), .B1(new_n460), .B2(new_n717), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n766), .A2(new_n767), .A3(new_n316), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n740), .A2(new_n895), .A3(new_n376), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n894), .A2(new_n757), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n712), .ZN(new_n898));
  NOR4_X1   g712(.A1(new_n898), .A2(new_n377), .A3(new_n316), .A4(new_n757), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n625), .A2(new_n249), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n823), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n898), .A2(new_n757), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n895), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n740), .A2(new_n673), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n897), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT112), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n898), .B2(new_n378), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n712), .A2(KEYINPUT112), .A3(new_n379), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n819), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT113), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n896), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n910), .A2(new_n911), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT114), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT50), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT50), .B1(new_n915), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n906), .B1(new_n919), .B2(KEYINPUT115), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT115), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n917), .A2(new_n918), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n893), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n595), .B1(new_n581), .B2(KEYINPUT102), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n377), .B1(new_n924), .B2(new_n753), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n895), .A3(new_n902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT48), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n899), .A2(new_n249), .A3(new_n625), .A4(new_n823), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n896), .A2(new_n719), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n927), .A2(new_n314), .A3(new_n928), .A4(new_n929), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n897), .A2(new_n905), .A3(new_n893), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n919), .B2(new_n931), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n892), .A2(new_n923), .A3(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(G952), .A2(G953), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT116), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n826), .B1(new_n933), .B2(new_n935), .ZN(G75));
  NOR2_X1   g750(.A1(new_n197), .A2(G952), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n300), .B1(new_n861), .B2(new_n884), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT56), .B1(new_n939), .B2(G210), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n418), .A2(new_n422), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(new_n436), .Z(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT55), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n938), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(G210), .ZN(new_n946));
  AOI211_X1 g760(.A(new_n946), .B(new_n300), .C1(new_n861), .C2(new_n884), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n947), .A2(KEYINPUT56), .A3(new_n943), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT117), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n940), .A2(new_n944), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n943), .B1(new_n947), .B2(KEYINPUT56), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT117), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n950), .A2(new_n951), .A3(new_n952), .A4(new_n938), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n949), .A2(new_n953), .ZN(G51));
  XOR2_X1   g768(.A(new_n796), .B(KEYINPUT57), .Z(new_n955));
  AOI21_X1  g769(.A(new_n885), .B1(new_n861), .B2(new_n884), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n887), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n706), .ZN(new_n958));
  INV_X1    g772(.A(new_n795), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n939), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n937), .B1(new_n958), .B2(new_n960), .ZN(G54));
  AND2_X1   g775(.A1(KEYINPUT58), .A2(G475), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n939), .A2(new_n240), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n240), .B1(new_n939), .B2(new_n962), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n963), .A2(new_n964), .A3(new_n937), .ZN(G60));
  INV_X1    g779(.A(KEYINPUT118), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n612), .A2(new_n618), .ZN(new_n967));
  NAND2_X1  g781(.A1(G478), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT59), .Z(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n861), .A2(new_n884), .ZN(new_n972));
  INV_X1    g786(.A(new_n885), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n971), .B1(new_n974), .B2(new_n886), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n966), .B1(new_n975), .B2(new_n937), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n970), .B1(new_n887), .B2(new_n956), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n977), .A2(KEYINPUT118), .A3(new_n938), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n967), .B1(new_n892), .B2(new_n969), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(G63));
  XNOR2_X1  g794(.A(KEYINPUT119), .B(KEYINPUT60), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n292), .A2(new_n300), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n984), .B1(new_n861), .B2(new_n884), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n938), .B1(new_n985), .B2(new_n365), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n648), .A2(new_n649), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n985), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n987), .A2(KEYINPUT120), .A3(new_n988), .A4(new_n990), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n988), .A2(KEYINPUT120), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n988), .A2(KEYINPUT120), .ZN(new_n993));
  INV_X1    g807(.A(new_n990), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n992), .B(new_n993), .C1(new_n994), .C2(new_n986), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n991), .A2(new_n995), .ZN(G66));
  INV_X1    g810(.A(G224), .ZN(new_n997));
  OAI21_X1  g811(.A(G953), .B1(new_n320), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n835), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n998), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n941), .B1(G898), .B2(new_n197), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(G69));
  INV_X1    g816(.A(KEYINPUT125), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n553), .B(new_n236), .Z(new_n1004));
  NOR2_X1   g818(.A1(new_n197), .A2(G900), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT122), .ZN(new_n1006));
  AND4_X1   g820(.A1(new_n718), .A2(new_n836), .A3(new_n800), .A4(new_n680), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1006), .B1(new_n925), .B2(new_n1007), .ZN(new_n1008));
  AND4_X1   g822(.A1(new_n1006), .A2(new_n754), .A3(new_n376), .A4(new_n1007), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n763), .B(new_n815), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1010), .A2(new_n761), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n663), .A2(new_n693), .A3(new_n746), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(KEYINPUT121), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT121), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n663), .A2(new_n693), .A3(new_n1014), .A4(new_n746), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1011), .B(new_n1016), .C1(new_n804), .C2(new_n802), .ZN(new_n1017));
  AOI211_X1 g831(.A(KEYINPUT123), .B(new_n1005), .C1(new_n1017), .C2(new_n197), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT123), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n815), .B1(new_n873), .B2(new_n661), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n925), .A2(new_n1007), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(KEYINPUT122), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n925), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1016), .A2(new_n1024), .A3(new_n877), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n197), .B1(new_n805), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1005), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1019), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n1003), .B(new_n1004), .C1(new_n1018), .C2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n197), .B1(G227), .B2(G900), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1004), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(KEYINPUT123), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1026), .A2(new_n1019), .A3(new_n1027), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1031), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(new_n827), .ZN(new_n1036));
  AOI211_X1 g850(.A(new_n681), .B(new_n757), .C1(new_n626), .C2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n701), .A2(new_n1037), .ZN(new_n1038));
  AND2_X1   g852(.A1(new_n1038), .A2(new_n815), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n683), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT62), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI211_X1 g856(.A(KEYINPUT62), .B(new_n683), .C1(new_n1013), .C2(new_n1015), .ZN(new_n1043));
  NOR3_X1   g857(.A1(new_n1042), .A2(new_n805), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1031), .B1(new_n1044), .B2(G953), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1045), .A2(KEYINPUT125), .ZN(new_n1046));
  OAI211_X1 g860(.A(new_n1029), .B(new_n1030), .C1(new_n1035), .C2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1004), .B1(new_n1018), .B2(new_n1028), .ZN(new_n1048));
  AND2_X1   g862(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1049));
  OAI21_X1  g863(.A(KEYINPUT62), .B1(new_n1049), .B2(new_n683), .ZN(new_n1050));
  INV_X1    g864(.A(new_n804), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1051), .A2(new_n801), .A3(new_n787), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1053));
  NAND4_X1  g867(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .A4(new_n1039), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1054), .A2(new_n197), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n1030), .B1(new_n1055), .B2(new_n1031), .ZN(new_n1056));
  AND3_X1   g870(.A1(new_n1048), .A2(new_n1056), .A3(KEYINPUT124), .ZN(new_n1057));
  AOI21_X1  g871(.A(KEYINPUT124), .B1(new_n1048), .B2(new_n1056), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1047), .B1(new_n1057), .B2(new_n1058), .ZN(G72));
  NOR2_X1   g873(.A1(new_n1017), .A2(new_n835), .ZN(new_n1060));
  XOR2_X1   g874(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1061));
  NOR2_X1   g875(.A1(new_n582), .A2(new_n300), .ZN(new_n1062));
  XNOR2_X1  g876(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  OAI211_X1 g877(.A(new_n545), .B(new_n554), .C1(new_n1060), .C2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n890), .A2(new_n884), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n583), .A2(new_n545), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n1063), .B1(new_n1066), .B2(new_n549), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n937), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1064), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g883(.A(new_n1063), .ZN(new_n1070));
  OAI21_X1  g884(.A(new_n1070), .B1(new_n1054), .B2(new_n835), .ZN(new_n1071));
  AOI21_X1  g885(.A(new_n1069), .B1(new_n667), .B2(new_n1071), .ZN(G57));
endmodule


