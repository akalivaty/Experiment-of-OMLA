//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT65), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n208), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n211), .B1(new_n214), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0024(.A(G238), .B(G244), .Z(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G226), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G250), .B(G257), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G87), .B(G97), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G107), .B(G116), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT67), .Z(new_n237));
  INV_X1    g0037(.A(G50), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G68), .ZN(new_n239));
  INV_X1    g0039(.A(G68), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n237), .B(new_n244), .ZN(G351));
  NAND2_X1  g0045(.A1(G33), .A2(G41), .ZN(new_n246));
  NAND3_X1  g0046(.A1(new_n246), .A2(G1), .A3(G13), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G232), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G1698), .ZN(new_n250));
  OAI211_X1 g0050(.A(new_n248), .B(new_n250), .C1(G226), .C2(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G97), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n247), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  OAI21_X1  g0057(.A(G274), .B1(new_n257), .B2(new_n212), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT68), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  AND2_X1   g0061(.A1(G1), .A2(G13), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(new_n246), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT68), .ZN(new_n264));
  INV_X1    g0064(.A(G41), .ZN(new_n265));
  INV_X1    g0065(.A(G45), .ZN(new_n266));
  AOI21_X1  g0066(.A(G1), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n263), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n247), .A2(new_n259), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G238), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT72), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n269), .A2(KEYINPUT72), .A3(new_n272), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n256), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI211_X1 g0079(.A(KEYINPUT13), .B(new_n256), .C1(new_n275), .C2(new_n276), .ZN(new_n280));
  OAI21_X1  g0080(.A(G169), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT14), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT73), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(new_n277), .B2(new_n278), .ZN(new_n284));
  INV_X1    g0084(.A(new_n256), .ZN(new_n285));
  INV_X1    g0085(.A(new_n276), .ZN(new_n286));
  AOI21_X1  g0086(.A(KEYINPUT72), .B1(new_n269), .B2(new_n272), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n288), .A2(KEYINPUT73), .A3(KEYINPUT13), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n277), .A2(new_n278), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n284), .A2(new_n289), .A3(G179), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(KEYINPUT13), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n290), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT14), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(new_n294), .A3(G169), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n282), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G20), .A2(G33), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n297), .A2(G50), .B1(G20), .B2(new_n240), .ZN(new_n298));
  INV_X1    g0098(.A(G77), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n206), .A2(G33), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n212), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n304), .A2(KEYINPUT11), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n302), .A2(new_n212), .ZN(new_n306));
  INV_X1    g0106(.A(G13), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(G1), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G20), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT70), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n306), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NOR3_X1   g0111(.A1(new_n307), .A2(new_n206), .A3(G1), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT70), .B1(new_n312), .B2(new_n303), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n205), .A2(G20), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(G68), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n312), .A2(new_n240), .ZN(new_n317));
  XNOR2_X1  g0117(.A(new_n317), .B(KEYINPUT12), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n304), .A2(KEYINPUT11), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n305), .A2(new_n316), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n296), .A2(new_n320), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n258), .A2(KEYINPUT68), .A3(new_n259), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n264), .B1(new_n263), .B2(new_n267), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(G226), .B2(new_n271), .ZN(new_n325));
  INV_X1    g0125(.A(G1698), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n248), .A2(G222), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n248), .A2(G223), .A3(G1698), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n327), .B(new_n328), .C1(new_n299), .C2(new_n248), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n257), .A2(new_n212), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n333), .A2(G169), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n202), .A2(G20), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT8), .B(G58), .ZN(new_n336));
  INV_X1    g0136(.A(G150), .ZN(new_n337));
  INV_X1    g0137(.A(new_n297), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n336), .A2(new_n300), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n306), .B1(new_n335), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n312), .A2(new_n303), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n238), .B1(new_n205), .B2(G20), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n342), .A2(new_n343), .B1(new_n238), .B2(new_n312), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n332), .A2(G179), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n334), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n248), .A2(G232), .A3(new_n326), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n248), .A2(G238), .A3(G1698), .ZN(new_n350));
  AND2_X1   g0150(.A1(KEYINPUT3), .A2(G33), .ZN(new_n351));
  NOR2_X1   g0151(.A1(KEYINPUT3), .A2(G33), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G107), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n349), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT69), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n247), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n356), .B2(new_n355), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n324), .B1(G244), .B2(new_n271), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G200), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n314), .A2(G77), .A3(new_n315), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n336), .A2(new_n338), .B1(new_n206), .B2(new_n299), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n300), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n303), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n312), .A2(new_n299), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n362), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G190), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n361), .B(new_n369), .C1(new_n370), .C2(new_n360), .ZN(new_n371));
  INV_X1    g0171(.A(G169), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n360), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G179), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n358), .A2(new_n359), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n368), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n371), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n325), .B2(new_n331), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n333), .B2(G190), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n335), .A2(new_n340), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n303), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT71), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n383), .A3(new_n344), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT9), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT71), .B1(new_n341), .B2(new_n345), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n385), .B1(new_n384), .B2(new_n386), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n380), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT10), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT10), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n380), .B(new_n391), .C1(new_n387), .C2(new_n388), .ZN(new_n392));
  AOI211_X1 g0192(.A(new_n348), .B(new_n377), .C1(new_n390), .C2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT7), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n248), .B2(G20), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n353), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n240), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G58), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n399), .A2(new_n240), .ZN(new_n400));
  NOR2_X1   g0200(.A1(G58), .A2(G68), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n297), .A2(G159), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n394), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT7), .B1(new_n353), .B2(new_n206), .ZN(new_n406));
  NOR4_X1   g0206(.A1(new_n351), .A2(new_n352), .A3(new_n395), .A4(G20), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n404), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(KEYINPUT16), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n410), .A3(new_n303), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n336), .B1(new_n205), .B2(G20), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n412), .A2(new_n342), .B1(new_n312), .B2(new_n336), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT74), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n411), .A2(KEYINPUT74), .A3(new_n413), .ZN(new_n416));
  NOR2_X1   g0216(.A1(G223), .A2(G1698), .ZN(new_n417));
  INV_X1    g0217(.A(G226), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(new_n418), .B2(G1698), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n248), .B1(G33), .B2(G87), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT75), .B1(new_n420), .B2(new_n247), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(G1698), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(G223), .B2(G1698), .ZN(new_n423));
  INV_X1    g0223(.A(G87), .ZN(new_n424));
  OAI22_X1  g0224(.A1(new_n423), .A2(new_n353), .B1(new_n252), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT75), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(new_n426), .A3(new_n330), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n421), .A2(new_n427), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n322), .A2(new_n323), .B1(new_n249), .B2(new_n270), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(G179), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n260), .A2(new_n268), .B1(new_n271), .B2(G232), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n425), .A2(new_n330), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n428), .A2(new_n430), .B1(new_n372), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n415), .A2(new_n416), .A3(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n435), .A2(KEYINPUT18), .ZN(new_n436));
  INV_X1    g0236(.A(new_n413), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n408), .A2(new_n409), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n306), .B1(new_n438), .B2(new_n394), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n437), .B1(new_n439), .B2(new_n410), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n420), .A2(new_n247), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n378), .B1(new_n429), .B2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n421), .A2(new_n431), .A3(new_n370), .A4(new_n427), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT17), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n440), .A2(new_n444), .B1(KEYINPUT76), .B2(new_n445), .ZN(new_n446));
  XOR2_X1   g0246(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n447));
  AND4_X1   g0247(.A1(new_n411), .A2(new_n444), .A3(new_n413), .A4(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n435), .A2(KEYINPUT18), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n436), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n293), .A2(G200), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n284), .A2(new_n289), .A3(G190), .A4(new_n290), .ZN(new_n455));
  INV_X1    g0255(.A(new_n320), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AND4_X1   g0257(.A1(new_n321), .A2(new_n393), .A3(new_n453), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT78), .ZN(new_n460));
  XNOR2_X1  g0260(.A(G97), .B(G107), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT6), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n462), .A2(new_n253), .A3(G107), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n466), .A2(G20), .B1(G77), .B2(new_n297), .ZN(new_n467));
  OAI21_X1  g0267(.A(G107), .B1(new_n406), .B2(new_n407), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n306), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n309), .A2(G97), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n205), .A2(G33), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT77), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n342), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n471), .B1(new_n475), .B2(new_n253), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n460), .B1(new_n469), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n464), .B1(new_n462), .B2(new_n461), .ZN(new_n478));
  OAI22_X1  g0278(.A1(new_n478), .A2(new_n206), .B1(new_n299), .B2(new_n338), .ZN(new_n479));
  INV_X1    g0279(.A(G107), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n480), .B1(new_n396), .B2(new_n397), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n303), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n476), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT78), .ZN(new_n484));
  XNOR2_X1  g0284(.A(KEYINPUT5), .B(G41), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n266), .A2(G1), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(new_n258), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n487), .A2(G257), .A3(new_n247), .ZN(new_n489));
  OAI211_X1 g0289(.A(G244), .B(new_n326), .C1(new_n351), .C2(new_n352), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n248), .A2(KEYINPUT4), .A3(G244), .A4(new_n326), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n248), .A2(G250), .A3(G1698), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n492), .A2(new_n493), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  AOI211_X1 g0296(.A(new_n488), .B(new_n489), .C1(new_n496), .C2(new_n330), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(G200), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n489), .B1(new_n496), .B2(new_n330), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n485), .A2(new_n486), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n263), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n499), .A2(new_n370), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n477), .B(new_n484), .C1(new_n498), .C2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n499), .A2(G179), .A3(new_n501), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n497), .B2(new_n372), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n482), .A2(new_n483), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n248), .A2(new_n206), .A3(G68), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT19), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(new_n300), .B2(new_n253), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n424), .A2(new_n253), .A3(new_n480), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT79), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT79), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n514), .A2(new_n424), .A3(new_n253), .A4(new_n480), .ZN(new_n515));
  NAND3_X1  g0315(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n513), .A2(new_n515), .B1(new_n206), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n303), .B1(new_n511), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n364), .A2(new_n312), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n474), .A2(G87), .A3(new_n342), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n247), .A2(G274), .A3(new_n486), .ZN(new_n522));
  OAI21_X1  g0322(.A(G250), .B1(new_n266), .B2(G1), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(new_n330), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n248), .A2(G238), .A3(new_n326), .ZN(new_n525));
  OAI211_X1 g0325(.A(G244), .B(G1698), .C1(new_n351), .C2(new_n352), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G116), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n524), .B1(new_n528), .B2(new_n330), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n521), .B1(G190), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g0330(.A1(new_n529), .A2(new_n378), .ZN(new_n531));
  AOI211_X1 g0331(.A(G179), .B(new_n524), .C1(new_n330), .C2(new_n528), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n528), .A2(new_n330), .ZN(new_n533));
  INV_X1    g0333(.A(new_n524), .ZN(new_n534));
  AOI21_X1  g0334(.A(G169), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n518), .B(new_n519), .C1(new_n475), .C2(new_n364), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n530), .A2(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n503), .A2(new_n507), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n309), .A2(G107), .ZN(new_n540));
  XNOR2_X1  g0340(.A(new_n540), .B(KEYINPUT25), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n474), .A2(G107), .A3(new_n342), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n206), .B(G87), .C1(new_n351), .C2(new_n352), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT22), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT22), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n248), .A2(new_n546), .A3(new_n206), .A4(G87), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT83), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n527), .B2(G20), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT23), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n206), .B2(G107), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n480), .A2(KEYINPUT23), .A3(G20), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n206), .A2(KEYINPUT83), .A3(G33), .A4(G116), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n548), .A2(new_n550), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT84), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n554), .A2(new_n550), .A3(new_n555), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n558), .B1(new_n545), .B2(new_n547), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT84), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n557), .A2(KEYINPUT24), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n559), .A2(new_n560), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n306), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n543), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n330), .B1(new_n486), .B2(new_n485), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n488), .B1(G264), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n248), .A2(G257), .A3(G1698), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n248), .A2(G250), .A3(new_n326), .ZN(new_n570));
  INV_X1    g0370(.A(G294), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n570), .C1(new_n252), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n330), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n372), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(G179), .B2(new_n574), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n566), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n556), .A2(KEYINPUT84), .A3(new_n564), .ZN(new_n578));
  INV_X1    g0378(.A(new_n561), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT24), .B1(new_n559), .B2(new_n560), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n578), .B(new_n303), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n543), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n568), .A2(new_n573), .A3(new_n370), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n487), .A2(G264), .A3(new_n247), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n501), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n585), .B1(new_n330), .B2(new_n572), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n583), .B1(new_n586), .B2(G200), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n581), .A2(new_n582), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(KEYINPUT85), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT85), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n566), .A2(new_n590), .A3(new_n587), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n577), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AND4_X1   g0392(.A1(G116), .A2(new_n311), .A3(new_n474), .A4(new_n313), .ZN(new_n593));
  INV_X1    g0393(.A(G116), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n308), .A2(G20), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n302), .A2(new_n212), .B1(G20), .B2(new_n594), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n494), .B(new_n206), .C1(G33), .C2(new_n253), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n596), .A2(KEYINPUT20), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT20), .B1(new_n596), .B2(new_n597), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n593), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n567), .A2(G270), .B1(new_n500), .B2(new_n263), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n248), .A2(G264), .A3(G1698), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n353), .A2(G303), .ZN(new_n604));
  OAI211_X1 g0404(.A(G257), .B(new_n326), .C1(new_n351), .C2(new_n352), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n330), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n601), .A2(new_n608), .A3(new_n374), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n372), .B1(new_n602), .B2(new_n607), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n311), .A2(new_n474), .A3(new_n313), .A4(G116), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(new_n595), .C1(new_n599), .C2(new_n598), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT80), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n609), .B1(new_n614), .B2(KEYINPUT21), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT81), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n602), .A2(new_n607), .A3(G190), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n601), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n378), .B1(new_n602), .B2(new_n607), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n619), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n621), .A2(KEYINPUT81), .A3(new_n601), .A4(new_n617), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT80), .ZN(new_n624));
  AOI211_X1 g0424(.A(new_n624), .B(KEYINPUT21), .C1(new_n610), .C2(new_n612), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n615), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(KEYINPUT82), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT82), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n612), .A2(G179), .A3(new_n607), .A4(new_n602), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n624), .B1(new_n610), .B2(new_n612), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT21), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n633), .A2(new_n625), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n629), .B1(new_n634), .B2(new_n623), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n539), .B(new_n592), .C1(new_n628), .C2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n459), .A2(new_n636), .ZN(G372));
  OAI211_X1 g0437(.A(new_n615), .B(new_n626), .C1(new_n566), .C2(new_n576), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n589), .A2(new_n591), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n539), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n521), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n529), .A2(G190), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n531), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n529), .A2(new_n374), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n537), .B(new_n644), .C1(G169), .C2(new_n529), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n505), .A2(new_n643), .A3(new_n645), .A4(new_n506), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  OAI21_X1  g0447(.A(KEYINPUT86), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n477), .A2(new_n484), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n505), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n643), .A2(new_n645), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n499), .A2(new_n501), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G169), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(new_n504), .B1(new_n482), .B2(new_n483), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT86), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n538), .A2(new_n655), .A3(new_n656), .A4(KEYINPUT26), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n648), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n640), .A2(new_n658), .A3(new_n645), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n458), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n433), .A2(new_n372), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n421), .A2(new_n431), .A3(new_n374), .A4(new_n427), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT18), .B1(new_n440), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n411), .A2(new_n413), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT18), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n434), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n376), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n296), .A2(new_n320), .B1(new_n457), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n664), .B(new_n667), .C1(new_n669), .C2(new_n449), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n390), .A2(new_n392), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n348), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n660), .A2(new_n672), .ZN(G369));
  NAND2_X1  g0473(.A1(new_n308), .A2(new_n206), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  XOR2_X1   g0475(.A(new_n675), .B(KEYINPUT87), .Z(new_n676));
  OAI21_X1  g0476(.A(G213), .B1(new_n674), .B2(KEYINPUT27), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n601), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n628), .B2(new_n635), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n634), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n592), .B1(new_n566), .B2(new_n682), .ZN(new_n689));
  INV_X1    g0489(.A(new_n577), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n682), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n634), .A2(new_n681), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n592), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n577), .A2(new_n682), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(KEYINPUT88), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT88), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n694), .A2(new_n698), .A3(new_n695), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n692), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n209), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n513), .A2(new_n594), .A3(new_n515), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n704), .A2(G1), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n215), .B2(new_n704), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n659), .A2(new_n682), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(KEYINPUT29), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT26), .B1(new_n650), .B2(new_n651), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n538), .A2(new_n655), .A3(new_n647), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n640), .A2(new_n645), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n712), .B1(new_n715), .B2(new_n682), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G330), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n681), .A2(KEYINPUT31), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n529), .A2(G179), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n653), .A2(new_n608), .A3(new_n574), .A4(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(KEYINPUT89), .B1(new_n608), .B2(new_n374), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n529), .A2(new_n568), .A3(new_n573), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT89), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n602), .A2(new_n607), .A3(new_n724), .A4(G179), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n722), .A2(new_n723), .A3(new_n499), .A4(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n721), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n726), .A2(new_n727), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n719), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT90), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n726), .A2(new_n732), .A3(new_n727), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(KEYINPUT90), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n729), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n681), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n731), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n627), .A2(KEYINPUT82), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n634), .A2(new_n629), .A3(new_n623), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n741), .A2(new_n539), .A3(new_n592), .A4(new_n682), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n718), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n717), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT91), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n717), .A2(KEYINPUT91), .A3(new_n744), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n709), .B1(new_n749), .B2(G1), .ZN(new_n750));
  XOR2_X1   g0550(.A(new_n750), .B(KEYINPUT92), .Z(G364));
  NOR2_X1   g0551(.A1(new_n307), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n205), .B1(new_n752), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n703), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n688), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(G330), .B2(new_n686), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n212), .B1(G20), .B2(new_n372), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G179), .A2(G200), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n206), .B1(new_n759), .B2(G190), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n571), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n206), .A2(new_n374), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(new_n370), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(KEYINPUT33), .A2(G317), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(KEYINPUT33), .A2(G317), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n763), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n761), .B(new_n767), .C1(G326), .C2(new_n769), .ZN(new_n770));
  OR3_X1    g0570(.A1(new_n206), .A2(KEYINPUT95), .A3(G190), .ZN(new_n771));
  OAI21_X1  g0571(.A(KEYINPUT95), .B1(new_n206), .B2(G190), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n771), .A2(new_n759), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G329), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n206), .A2(new_n370), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n374), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n353), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n378), .A2(G179), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n206), .A2(G190), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n777), .ZN(new_n785));
  INV_X1    g0585(.A(G311), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n782), .A2(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n771), .A2(new_n772), .A3(new_n781), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n780), .B(new_n787), .C1(G283), .C2(new_n789), .ZN(new_n790));
  AND3_X1   g0590(.A1(new_n770), .A2(new_n775), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(KEYINPUT97), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n248), .B1(new_n782), .B2(new_n424), .C1(new_n240), .C2(new_n763), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n760), .B(KEYINPUT96), .Z(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n253), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n794), .B(new_n797), .C1(G50), .C2(new_n769), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n778), .A2(new_n399), .B1(new_n785), .B2(new_n299), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT94), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n799), .A2(KEYINPUT94), .B1(new_n789), .B2(G107), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n798), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G159), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n773), .A2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT32), .Z(new_n805));
  OAI21_X1  g0605(.A(new_n793), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n792), .A2(KEYINPUT97), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n758), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n755), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n209), .A2(new_n248), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n810), .B1(KEYINPUT93), .B2(G355), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(KEYINPUT93), .B2(G355), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n244), .A2(new_n266), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n702), .A2(new_n248), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n814), .B1(G45), .B2(new_n215), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n812), .B1(G116), .B2(new_n209), .C1(new_n813), .C2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(G13), .A2(G33), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(G20), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n819), .A2(new_n758), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n809), .B1(new_n816), .B2(new_n820), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n819), .B(KEYINPUT98), .Z(new_n822));
  OAI211_X1 g0622(.A(new_n808), .B(new_n821), .C1(new_n686), .C2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n757), .A2(new_n823), .ZN(G396));
  NAND2_X1  g0624(.A1(new_n376), .A2(KEYINPUT100), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT100), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n373), .A2(new_n826), .A3(new_n368), .A4(new_n375), .ZN(new_n827));
  AND3_X1   g0627(.A1(new_n825), .A2(new_n827), .A3(new_n371), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n681), .A2(new_n368), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n828), .A2(new_n829), .B1(new_n668), .B2(new_n681), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n710), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n659), .A2(new_n682), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n755), .B1(new_n833), .B2(new_n744), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n744), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n758), .A2(new_n817), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT99), .Z(new_n837));
  OAI21_X1  g0637(.A(new_n755), .B1(new_n837), .B2(G77), .ZN(new_n838));
  INV_X1    g0638(.A(new_n778), .ZN(new_n839));
  INV_X1    g0639(.A(new_n785), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G143), .A2(new_n839), .B1(new_n840), .B2(G159), .ZN(new_n841));
  INV_X1    g0641(.A(G137), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n842), .B2(new_n768), .C1(new_n337), .C2(new_n763), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT34), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n789), .A2(G68), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n248), .B1(new_n760), .B2(new_n399), .C1(new_n238), .C2(new_n782), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(G132), .B2(new_n774), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n843), .A2(new_n844), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n788), .A2(new_n424), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(G311), .B2(new_n774), .ZN(new_n852));
  INV_X1    g0652(.A(new_n782), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n248), .B1(new_n853), .B2(G107), .ZN(new_n854));
  AOI22_X1  g0654(.A1(G294), .A2(new_n839), .B1(new_n840), .B2(G116), .ZN(new_n855));
  INV_X1    g0655(.A(new_n763), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G303), .A2(new_n769), .B1(new_n856), .B2(G283), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n852), .A2(new_n854), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  OAI22_X1  g0658(.A1(new_n849), .A2(new_n850), .B1(new_n797), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n838), .B1(new_n859), .B2(new_n758), .ZN(new_n860));
  INV_X1    g0660(.A(new_n830), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n860), .B1(new_n861), .B2(new_n818), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n835), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G384));
  AND2_X1   g0664(.A1(new_n466), .A2(KEYINPUT35), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n466), .A2(KEYINPUT35), .ZN(new_n866));
  NOR4_X1   g0666(.A1(new_n865), .A2(new_n866), .A3(new_n214), .A4(new_n594), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT36), .ZN(new_n868));
  OR3_X1    g0668(.A1(new_n400), .A2(new_n215), .A3(new_n299), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n205), .B(G13), .C1(new_n869), .C2(new_n239), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n681), .A2(new_n320), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n321), .A2(new_n457), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n457), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n320), .B(new_n681), .C1(new_n874), .C2(new_n296), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n830), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n733), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n732), .B1(new_n726), .B2(new_n727), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n877), .A2(new_n728), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n737), .B1(new_n879), .B2(new_n682), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n681), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n742), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n876), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT40), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT16), .B1(new_n408), .B2(new_n409), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT101), .B1(new_n885), .B2(new_n306), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT101), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n405), .A2(new_n887), .A3(new_n303), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n410), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n413), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT102), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT102), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n889), .A2(new_n892), .A3(new_n413), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n678), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n452), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n444), .A2(new_n411), .A3(new_n413), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n889), .A2(new_n892), .A3(new_n413), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n892), .B1(new_n889), .B2(new_n413), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n902), .B2(new_n434), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n897), .B1(new_n903), .B2(new_n894), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n415), .A2(new_n416), .A3(new_n678), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT37), .B1(new_n440), .B2(new_n444), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n435), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(KEYINPUT38), .B(new_n896), .C1(new_n904), .C2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT38), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n891), .A2(new_n434), .A3(new_n893), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n894), .A2(new_n911), .A3(new_n898), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n908), .B1(new_n912), .B2(KEYINPUT37), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n449), .B1(KEYINPUT18), .B2(new_n435), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n894), .B1(new_n914), .B2(new_n436), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n910), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n909), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n883), .A2(new_n884), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n912), .A2(KEYINPUT37), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n919), .A2(new_n907), .B1(new_n452), .B2(new_n895), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n411), .A2(KEYINPUT74), .A3(new_n413), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n921), .A2(new_n414), .A3(new_n679), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n898), .B1(new_n440), .B2(new_n663), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT37), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n907), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n664), .B(new_n667), .C1(new_n446), .C2(new_n448), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n922), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n928), .A2(KEYINPUT103), .A3(new_n910), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT103), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n924), .A2(new_n907), .B1(new_n926), .B2(new_n922), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n930), .B1(new_n931), .B2(KEYINPUT38), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n920), .A2(KEYINPUT38), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n876), .A2(new_n882), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT40), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n918), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n458), .A2(new_n882), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n718), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n937), .B2(new_n936), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n909), .A2(new_n916), .A3(KEYINPUT39), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n321), .A2(new_n681), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n940), .B(new_n941), .C1(new_n933), .C2(KEYINPUT39), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n678), .B1(new_n664), .B2(new_n667), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n681), .B1(new_n825), .B2(new_n827), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n832), .A2(new_n945), .B1(new_n873), .B2(new_n875), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n943), .B1(new_n917), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n458), .B1(new_n711), .B2(new_n716), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n672), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n948), .B(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n939), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n205), .B2(new_n752), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n939), .A2(new_n951), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n871), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT104), .Z(G367));
  OAI21_X1  g0756(.A(new_n820), .B1(new_n209), .B2(new_n364), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n814), .B2(new_n232), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n778), .A2(new_n337), .B1(new_n785), .B2(new_n238), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n353), .B(new_n959), .C1(G58), .C2(new_n853), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n795), .A2(G68), .ZN(new_n961));
  AOI22_X1  g0761(.A1(G143), .A2(new_n769), .B1(new_n856), .B2(G159), .ZN(new_n962));
  AOI22_X1  g0762(.A1(G77), .A2(new_n789), .B1(new_n774), .B2(G137), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n960), .A2(new_n961), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  AOI22_X1  g0764(.A1(G311), .A2(new_n769), .B1(new_n856), .B2(G294), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n782), .A2(new_n594), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n965), .B1(KEYINPUT46), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(KEYINPUT108), .B(G317), .ZN(new_n968));
  AOI22_X1  g0768(.A1(G97), .A2(new_n789), .B1(new_n774), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n353), .B1(new_n778), .B2(new_n783), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G283), .B2(new_n840), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n760), .A2(new_n480), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n966), .B2(KEYINPUT46), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n969), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n964), .B1(new_n967), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n809), .B(new_n958), .C1(new_n976), .C2(new_n758), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n538), .B1(new_n641), .B2(new_n682), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n681), .A2(new_n537), .A3(new_n536), .A4(new_n521), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(new_n822), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT107), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n649), .A2(new_n681), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n503), .A2(new_n984), .A3(new_n507), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n649), .A2(new_n681), .A3(new_n505), .ZN(new_n986));
  AND2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(new_n697), .B2(new_n699), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT45), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n697), .A2(new_n699), .A3(new_n987), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT44), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n692), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n694), .B1(new_n691), .B2(new_n693), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n687), .B(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n747), .B2(new_n748), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n989), .A2(new_n692), .A3(new_n992), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n994), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n999), .A2(new_n749), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n703), .B(KEYINPUT41), .Z(new_n1001));
  OAI21_X1  g0801(.A(new_n753), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(KEYINPUT106), .B1(new_n692), .B2(new_n987), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT106), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n987), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n688), .A2(new_n1004), .A3(new_n691), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  OR3_X1    g0810(.A1(new_n694), .A2(new_n987), .A3(KEYINPUT105), .ZN(new_n1011));
  OAI21_X1  g0811(.A(KEYINPUT105), .B1(new_n694), .B2(new_n987), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n507), .B1(new_n987), .B2(new_n690), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1013), .A2(KEYINPUT42), .B1(new_n682), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(KEYINPUT42), .B2(new_n1013), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n1017));
  AND2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1003), .A2(new_n1008), .A3(new_n1006), .ZN(new_n1019));
  AND3_X1   g0819(.A1(new_n1010), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1018), .B1(new_n1010), .B2(new_n1019), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n983), .B1(new_n1002), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1001), .B1(new_n999), .B2(new_n749), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1022), .B(new_n983), .C1(new_n754), .C2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n982), .B1(new_n1023), .B2(new_n1026), .ZN(G387));
  NOR2_X1   g0827(.A1(new_n997), .A2(new_n704), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n996), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n749), .B2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n229), .A2(G45), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n814), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1031), .A2(new_n1032), .B1(new_n706), .B2(new_n810), .ZN(new_n1033));
  OR3_X1    g0833(.A1(new_n336), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1034));
  OAI21_X1  g0834(.A(KEYINPUT50), .B1(new_n336), .B2(G50), .ZN(new_n1035));
  AOI21_X1  g0835(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n706), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1033), .A2(new_n1037), .B1(new_n480), .B2(new_n702), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n820), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n755), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(G283), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n782), .A2(new_n571), .B1(new_n760), .B2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n839), .A2(new_n968), .B1(new_n840), .B2(G303), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n786), .B2(new_n763), .C1(new_n779), .C2(new_n768), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n1045), .B2(new_n1044), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT49), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n788), .A2(new_n594), .ZN(new_n1051));
  AOI211_X1 g0851(.A(new_n248), .B(new_n1051), .C1(G326), .C2(new_n774), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1049), .A2(new_n1050), .A3(new_n1052), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n796), .A2(new_n364), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n782), .A2(new_n299), .B1(new_n785), .B2(new_n240), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n353), .B(new_n1055), .C1(G50), .C2(new_n839), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n336), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G159), .A2(new_n769), .B1(new_n856), .B2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G97), .A2(new_n789), .B1(new_n774), .B2(G150), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1054), .A2(new_n1056), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1040), .B1(new_n1061), .B2(new_n758), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n691), .B2(new_n822), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT109), .Z(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n1029), .B2(new_n754), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1030), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT110), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT110), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1030), .A2(new_n1068), .A3(new_n1065), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(G393));
  INV_X1    g0870(.A(new_n998), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1071), .A2(new_n993), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n754), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n795), .A2(G77), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1074), .B1(new_n238), .B2(new_n763), .C1(new_n336), .C2(new_n785), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT111), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n768), .A2(new_n337), .B1(new_n778), .B2(new_n803), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT51), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n774), .A2(G143), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n353), .B(new_n851), .C1(G68), .C2(new_n853), .ZN(new_n1080));
  AND4_X1   g0880(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n769), .A2(G317), .B1(new_n839), .B2(G311), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT52), .Z(new_n1083));
  NAND2_X1  g0883(.A1(new_n789), .A2(G107), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n353), .B1(new_n785), .B2(new_n571), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n763), .A2(new_n783), .B1(new_n760), .B2(new_n594), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(G283), .C2(new_n853), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n774), .A2(G322), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1083), .A2(new_n1084), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT112), .Z(new_n1090));
  OAI21_X1  g0890(.A(new_n758), .B1(new_n1081), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n987), .A2(new_n819), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n814), .A2(new_n236), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1039), .B1(G97), .B2(new_n702), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n809), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1091), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1073), .A2(new_n1096), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1072), .A2(new_n997), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n704), .B1(new_n1072), .B2(new_n997), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(G390));
  OAI21_X1  g0901(.A(new_n755), .B1(new_n837), .B2(new_n1057), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n846), .B1(new_n571), .B2(new_n773), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT115), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n248), .B1(new_n853), .B2(G87), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G116), .A2(new_n839), .B1(new_n840), .B2(G97), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G283), .A2(new_n769), .B1(new_n856), .B2(G107), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1074), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n782), .A2(new_n337), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT53), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n774), .A2(G125), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n238), .C2(new_n788), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n795), .A2(G159), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n839), .A2(G132), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(KEYINPUT54), .B(G143), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n353), .B1(new_n840), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(G128), .A2(new_n769), .B1(new_n856), .B2(G137), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1113), .A2(new_n1114), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1104), .A2(new_n1108), .B1(new_n1112), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1102), .B1(new_n1120), .B2(new_n758), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n909), .A2(new_n916), .A3(KEYINPUT39), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n929), .A2(new_n932), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT39), .B1(new_n1123), .B2(new_n909), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1121), .B1(new_n1125), .B2(new_n818), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT116), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n876), .A2(G330), .A3(new_n882), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n832), .A2(new_n945), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n873), .A2(new_n875), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n941), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT39), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT103), .B1(new_n928), .B2(new_n910), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n931), .A2(new_n930), .A3(KEYINPUT38), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n913), .A2(new_n915), .A3(new_n910), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1132), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1131), .B1(new_n1137), .B2(new_n940), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n715), .A2(new_n682), .A3(new_n828), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1139), .A2(new_n945), .B1(new_n873), .B2(new_n875), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n933), .A2(new_n1140), .A3(new_n941), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1128), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1123), .A2(new_n909), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n941), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1139), .A2(new_n945), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1130), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1143), .B(new_n1144), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n743), .A2(new_n861), .A3(new_n1130), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1147), .B(new_n1148), .C1(new_n1125), .C2(new_n1131), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1142), .A2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1127), .B1(new_n753), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT117), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1127), .B(KEYINPUT117), .C1(new_n753), .C2(new_n1150), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT114), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n458), .A2(G330), .A3(new_n882), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n949), .A2(new_n1157), .A3(new_n672), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1130), .B1(new_n743), .B2(new_n861), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1129), .B1(new_n1128), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n882), .A2(G330), .A3(new_n861), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1146), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1162), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1158), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n1142), .B2(new_n1149), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(KEYINPUT113), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1165), .A2(KEYINPUT113), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1142), .A2(new_n1149), .A3(new_n1164), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n703), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1156), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n1165), .A2(KEYINPUT113), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1171), .B1(new_n1173), .B2(new_n1166), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT114), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1155), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(G378));
  INV_X1    g0977(.A(KEYINPUT119), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n348), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n671), .A2(new_n1179), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n384), .A2(new_n386), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(new_n679), .ZN(new_n1182));
  OR2_X1    g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1183), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT118), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n942), .A2(new_n947), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1191), .B1(new_n942), .B2(new_n947), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n718), .B1(new_n918), .B2(new_n935), .ZN(new_n1194));
  NOR3_X1   g0994(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n884), .B1(new_n883), .B2(new_n1143), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n882), .A2(new_n1130), .A3(new_n884), .A4(new_n861), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n909), .B2(new_n916), .ZN(new_n1198));
  OAI21_X1  g0998(.A(G330), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1191), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n948), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n942), .A2(new_n947), .A3(new_n1191), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1199), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1178), .B1(new_n1195), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1194), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1201), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(new_n1206), .A3(KEYINPUT119), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1204), .A2(new_n754), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT120), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1188), .A2(new_n817), .A3(new_n1189), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n755), .B1(new_n837), .B2(G50), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G33), .A2(G41), .ZN(new_n1212));
  AOI211_X1 g1012(.A(G50), .B(new_n1212), .C1(new_n353), .C2(new_n265), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n763), .A2(new_n253), .B1(new_n768), .B2(new_n594), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n778), .A2(new_n480), .B1(new_n785), .B2(new_n364), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n265), .B(new_n353), .C1(new_n782), .C2(new_n299), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G58), .A2(new_n789), .B1(new_n774), .B2(G283), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n961), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT58), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1213), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(G128), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1222), .A2(new_n778), .B1(new_n782), .B2(new_n1115), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1223), .B1(G137), .B2(new_n840), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G125), .A2(new_n769), .B1(new_n856), .B2(G132), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n796), .C2(new_n337), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1212), .B1(new_n788), .B2(new_n803), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(G124), .B2(new_n774), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1226), .A2(KEYINPUT59), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1221), .B1(new_n1220), .B2(new_n1219), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1211), .B1(new_n1232), .B2(new_n758), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1210), .A2(new_n1233), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1208), .A2(new_n1209), .A3(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1209), .B1(new_n1208), .B2(new_n1234), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1205), .A2(new_n1206), .A3(KEYINPUT119), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT119), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1158), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1170), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT121), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1170), .A2(KEYINPUT121), .A3(new_n1240), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT57), .B1(new_n1239), .B2(new_n1245), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1205), .A2(new_n1206), .A3(KEYINPUT57), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1170), .A2(KEYINPUT121), .A3(new_n1240), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT121), .B1(new_n1170), .B2(new_n1240), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1247), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n703), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n1235), .A2(new_n1236), .B1(new_n1246), .B2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT122), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1252), .A2(KEYINPUT122), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(G375));
  NAND2_X1  g1056(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1257), .A2(new_n1240), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1258), .A2(new_n1001), .A3(new_n1164), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n753), .B(KEYINPUT123), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1257), .A2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n755), .B1(new_n837), .B2(G68), .ZN(new_n1262));
  XOR2_X1   g1062(.A(new_n1262), .B(KEYINPUT124), .Z(new_n1263));
  OAI22_X1  g1063(.A1(new_n778), .A2(new_n1041), .B1(new_n785), .B2(new_n480), .ZN(new_n1264));
  AOI211_X1 g1064(.A(new_n248), .B(new_n1264), .C1(G97), .C2(new_n853), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(G294), .A2(new_n769), .B1(new_n856), .B2(G116), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(G77), .A2(new_n789), .B1(new_n774), .B2(G303), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1054), .A2(new_n1265), .A3(new_n1266), .A4(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n796), .A2(new_n238), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n842), .A2(new_n778), .B1(new_n782), .B2(new_n803), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n353), .B(new_n1270), .C1(G150), .C2(new_n840), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G132), .A2(new_n769), .B1(new_n856), .B2(new_n1116), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(G58), .A2(new_n789), .B1(new_n774), .B2(G128), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1268), .B1(new_n1269), .B2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1263), .B1(new_n758), .B2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1130), .B2(new_n818), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1261), .A2(new_n1277), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1259), .A2(new_n1278), .ZN(G381));
  NAND4_X1  g1079(.A1(new_n1067), .A2(new_n757), .A3(new_n823), .A4(new_n1069), .ZN(new_n1280));
  NOR4_X1   g1080(.A1(new_n1280), .A2(G390), .A3(G384), .A4(G381), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1022), .B1(new_n1024), .B2(new_n754), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT107), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1025), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1155), .A2(new_n1174), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1281), .A2(new_n1284), .A3(new_n982), .A4(new_n1285), .ZN(new_n1286));
  OR2_X1    g1086(.A1(G375), .A2(new_n1286), .ZN(G407));
  NAND3_X1  g1087(.A1(new_n1285), .A2(G213), .A3(new_n680), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G407), .B(G213), .C1(G375), .C2(new_n1288), .ZN(G409));
  NOR2_X1   g1089(.A1(new_n1195), .A2(new_n1203), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1290), .A2(new_n1260), .B1(new_n1210), .B2(new_n1233), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1239), .A2(new_n1245), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1291), .B1(new_n1292), .B2(new_n1001), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1285), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1252), .B2(new_n1176), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT125), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n680), .A2(G213), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1294), .B(KEYINPUT125), .C1(new_n1252), .C2(new_n1176), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1164), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(new_n1258), .A3(KEYINPUT60), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n703), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1258), .B1(KEYINPUT60), .B2(new_n1301), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  OR3_X1    g1105(.A1(new_n1305), .A2(new_n863), .A3(new_n1278), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n863), .B1(new_n1305), .B2(new_n1278), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n680), .A2(G213), .A3(G2897), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1311), .A2(new_n1308), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1300), .B1(new_n1309), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G393), .A2(G396), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(new_n1280), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G390), .B1(new_n1284), .B2(new_n982), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n982), .ZN(new_n1317));
  AOI211_X1 g1117(.A(new_n1317), .B(new_n1100), .C1(new_n1283), .C2(new_n1025), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1315), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(G387), .A2(new_n1100), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1315), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1284), .A2(new_n982), .A3(G390), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT61), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1319), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  AND2_X1   g1125(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1310), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1325), .B1(new_n1326), .B2(new_n1328), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1297), .A2(new_n1298), .A3(new_n1311), .A4(new_n1299), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1327), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1313), .A2(new_n1329), .A3(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1312), .A2(new_n1309), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1324), .B1(new_n1326), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT62), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1330), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1326), .A2(KEYINPUT62), .A3(new_n1311), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1334), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1319), .A2(new_n1323), .ZN(new_n1339));
  XOR2_X1   g1139(.A(new_n1339), .B(KEYINPUT126), .Z(new_n1340));
  OAI21_X1  g1140(.A(new_n1332), .B1(new_n1338), .B2(new_n1340), .ZN(G405));
  AND3_X1   g1141(.A1(new_n1319), .A2(new_n1323), .A3(new_n1310), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1310), .B1(new_n1319), .B2(new_n1323), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1255), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1346), .A2(new_n1253), .A3(new_n1285), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT127), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(G375), .A2(KEYINPUT127), .A3(new_n1285), .ZN(new_n1350));
  OR2_X1    g1150(.A1(new_n1252), .A2(new_n1176), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1349), .A2(new_n1350), .A3(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1345), .A2(new_n1352), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1344), .A2(new_n1351), .A3(new_n1349), .A4(new_n1350), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1353), .A2(new_n1354), .ZN(G402));
endmodule


