//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n796, new_n797, new_n798, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT67), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT66), .B(G190gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G183gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT24), .ZN(new_n207));
  INV_X1    g006(.A(G183gat), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n209), .A2(KEYINPUT66), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(KEYINPUT66), .ZN(new_n211));
  OAI211_X1 g010(.A(KEYINPUT67), .B(new_n208), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n205), .A2(new_n207), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT68), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n205), .A2(new_n212), .A3(KEYINPUT68), .A4(new_n207), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(G169gat), .B2(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(new_n225), .B2(KEYINPUT23), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n217), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n207), .B1(G183gat), .B2(G190gat), .ZN(new_n231));
  XOR2_X1   g030(.A(KEYINPUT64), .B(G176gat), .Z(new_n232));
  INV_X1    g031(.A(G169gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(KEYINPUT23), .A3(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n223), .A2(new_n231), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n224), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n217), .A2(KEYINPUT69), .A3(new_n227), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n230), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n239));
  INV_X1    g038(.A(new_n204), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT27), .B(G183gat), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n242), .B(KEYINPUT28), .Z(new_n243));
  INV_X1    g042(.A(KEYINPUT26), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT71), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n246), .B(new_n221), .C1(new_n244), .C2(new_n225), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n247), .A3(new_n206), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n238), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(G127gat), .B(G134gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n250), .B1(KEYINPUT72), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n252), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n202), .B1(new_n249), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n249), .A2(new_n256), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n238), .A2(KEYINPUT73), .A3(new_n255), .A4(new_n248), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G227gat), .A2(G233gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT33), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G15gat), .B(G43gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT74), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n265), .B(G71gat), .ZN(new_n266));
  INV_X1    g065(.A(G99gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n257), .A2(new_n261), .A3(new_n258), .A4(new_n259), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT34), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n271), .A2(KEYINPUT34), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n262), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(KEYINPUT32), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n274), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n279), .B(new_n272), .C1(new_n263), .C2(new_n269), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n275), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n278), .B1(new_n275), .B2(new_n280), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT29), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n249), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G226gat), .A2(G233gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT76), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(KEYINPUT77), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT77), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT29), .B1(new_n238), .B2(new_n248), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n290), .B1(new_n291), .B2(new_n287), .ZN(new_n292));
  NAND2_X1  g091(.A1(G211gat), .A2(G218gat), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G197gat), .B(G204gat), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n295), .B2(KEYINPUT22), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(G211gat), .B2(G218gat), .ZN(new_n297));
  INV_X1    g096(.A(G211gat), .ZN(new_n298));
  INV_X1    g097(.A(G218gat), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT22), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n295), .B1(new_n300), .B2(new_n294), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n249), .A2(new_n287), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n289), .A2(new_n292), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT78), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n249), .ZN(new_n307));
  MUX2_X1   g106(.A(new_n291), .B(new_n307), .S(new_n287), .Z(new_n308));
  OR2_X1    g107(.A1(new_n308), .A2(new_n302), .ZN(new_n309));
  XNOR2_X1  g108(.A(G8gat), .B(G36gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(G64gat), .B(G92gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n306), .A2(KEYINPUT30), .A3(new_n309), .A4(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n289), .A2(new_n292), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n315), .A2(new_n305), .A3(new_n302), .A4(new_n303), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n304), .A2(KEYINPUT78), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n316), .A2(new_n309), .A3(new_n317), .A4(new_n313), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT30), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(new_n309), .A3(new_n317), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n312), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n314), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT6), .ZN(new_n324));
  INV_X1    g123(.A(G148gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G141gat), .ZN(new_n326));
  XOR2_X1   g125(.A(KEYINPUT82), .B(G141gat), .Z(new_n327));
  OAI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(new_n325), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT83), .ZN(new_n329));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330));
  INV_X1    g129(.A(G155gat), .ZN(new_n331));
  INV_X1    g130(.A(G162gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n330), .B1(new_n333), .B2(KEYINPUT2), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G141gat), .B(G148gat), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(KEYINPUT80), .ZN(new_n337));
  INV_X1    g136(.A(new_n330), .ZN(new_n338));
  XOR2_X1   g137(.A(KEYINPUT81), .B(KEYINPUT2), .Z(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n330), .B(KEYINPUT79), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n340), .A2(new_n333), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n335), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(KEYINPUT3), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n256), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT5), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n255), .A3(new_n342), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353));
  OR3_X1    g152(.A1(new_n352), .A2(KEYINPUT85), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n353), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n351), .A2(KEYINPUT4), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(KEYINPUT85), .A3(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n349), .A2(new_n350), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n355), .A2(KEYINPUT84), .A3(new_n356), .ZN(new_n359));
  OR3_X1    g158(.A1(new_n351), .A2(KEYINPUT84), .A3(KEYINPUT4), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n359), .A2(new_n347), .A3(new_n348), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n256), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n351), .ZN(new_n363));
  INV_X1    g162(.A(new_n348), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n350), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n358), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368));
  INV_X1    g167(.A(G85gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT0), .B(G57gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(new_n371), .Z(new_n372));
  OAI21_X1  g171(.A(new_n324), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n367), .A2(new_n372), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT86), .ZN(new_n377));
  XOR2_X1   g176(.A(KEYINPUT31), .B(G50gat), .Z(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G228gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n302), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n344), .B2(KEYINPUT29), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT29), .B1(new_n381), .B2(KEYINPUT87), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(KEYINPUT87), .B2(new_n297), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT3), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n385), .A2(new_n386), .B1(new_n335), .B2(new_n342), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n380), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n381), .A2(KEYINPUT29), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n389), .A2(KEYINPUT88), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n386), .B1(new_n389), .B2(KEYINPUT88), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n343), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n382), .A2(new_n392), .A3(G228gat), .A4(G233gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G22gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n394), .A2(G22gat), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n379), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n379), .A2(KEYINPUT89), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n395), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(KEYINPUT89), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n283), .A2(new_n323), .A3(new_n375), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT91), .ZN(new_n406));
  NOR3_X1   g205(.A1(new_n281), .A2(new_n282), .A3(new_n403), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT91), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n407), .A2(new_n408), .A3(new_n375), .A4(new_n323), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(KEYINPUT35), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n314), .A2(new_n320), .A3(new_n322), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n373), .B(new_n374), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n403), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n282), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT36), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n275), .A2(new_n280), .A3(new_n278), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n415), .A2(new_n416), .ZN(new_n419));
  NAND2_X1  g218(.A1(KEYINPUT75), .A2(KEYINPUT36), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n419), .B(new_n420), .C1(new_n281), .C2(new_n282), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n413), .A2(new_n418), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT90), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT39), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n363), .A2(new_n364), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n347), .A2(new_n357), .A3(new_n354), .ZN(new_n426));
  AOI211_X1 g225(.A(new_n424), .B(new_n425), .C1(new_n426), .C2(new_n364), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n424), .A3(new_n364), .ZN(new_n428));
  INV_X1    g227(.A(new_n372), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n423), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT40), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n411), .A2(new_n433), .A3(new_n374), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT37), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n316), .A2(new_n435), .A3(new_n309), .A4(new_n317), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n315), .A2(new_n381), .A3(new_n303), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n437), .B(KEYINPUT37), .C1(new_n381), .C2(new_n308), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT38), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n436), .A2(new_n438), .A3(new_n439), .A4(new_n312), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n412), .A2(new_n318), .A3(new_n440), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n436), .A2(new_n312), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n321), .A2(KEYINPUT37), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n439), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n434), .B(new_n404), .C1(new_n441), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n422), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT35), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n405), .A2(KEYINPUT91), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n410), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT17), .ZN(new_n450));
  OR3_X1    g249(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n451), .A2(new_n452), .B1(G29gat), .B2(G36gat), .ZN(new_n453));
  INV_X1    g252(.A(G50gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(G43gat), .ZN(new_n455));
  INV_X1    g254(.A(G43gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(G50gat), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT93), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n455), .B2(new_n457), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT15), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G43gat), .B(G50gat), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(KEYINPUT15), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n453), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n455), .A2(new_n457), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT93), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n463), .A2(new_n458), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT15), .ZN(new_n469));
  INV_X1    g268(.A(new_n453), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n450), .B1(new_n465), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n464), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n470), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n459), .A2(new_n460), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n453), .B1(new_n475), .B2(KEYINPUT15), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n474), .A2(new_n476), .A3(KEYINPUT94), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT94), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n465), .B2(new_n471), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n450), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT95), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT94), .B1(new_n474), .B2(new_n476), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n478), .A3(new_n471), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT95), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n450), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n472), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488));
  INV_X1    g287(.A(G92gat), .ZN(new_n489));
  AOI22_X1  g288(.A1(KEYINPUT8), .A2(new_n488), .B1(new_n369), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT7), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(new_n369), .B2(new_n489), .ZN(new_n492));
  NAND3_X1  g291(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  XOR2_X1   g293(.A(G99gat), .B(G106gat), .Z(new_n495));
  OR2_X1    g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT98), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n495), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT99), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n494), .A2(KEYINPUT98), .A3(new_n495), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n500), .B1(new_n499), .B2(new_n501), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n487), .A2(KEYINPUT100), .A3(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(G190gat), .B(G218gat), .Z(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT101), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT100), .B1(new_n502), .B2(new_n503), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n484), .B1(new_n487), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n505), .B(new_n509), .C1(new_n511), .C2(new_n504), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT41), .ZN(new_n513));
  NAND2_X1  g312(.A1(G232gat), .A2(G233gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n472), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n485), .B1(new_n484), .B2(new_n450), .ZN(new_n517));
  AOI211_X1 g316(.A(KEYINPUT95), .B(KEYINPUT17), .C1(new_n482), .C2(new_n483), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n510), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n484), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n504), .ZN(new_n522));
  AOI22_X1  g321(.A1(new_n521), .A2(new_n522), .B1(new_n508), .B2(new_n507), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n514), .A2(new_n513), .ZN(new_n524));
  NAND3_X1  g323(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .A4(new_n505), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n506), .A2(KEYINPUT101), .ZN(new_n527));
  XNOR2_X1  g326(.A(G134gat), .B(G162gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n515), .A2(new_n526), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n529), .B1(new_n515), .B2(new_n526), .ZN(new_n531));
  XNOR2_X1  g330(.A(G127gat), .B(G155gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(G231gat), .A2(G233gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535));
  INV_X1    g334(.A(G1gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT16), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(G1gat), .B2(new_n535), .ZN(new_n539));
  INV_X1    g338(.A(G8gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT21), .ZN(new_n542));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT9), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G71gat), .B(G78gat), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n543), .A2(KEYINPUT97), .ZN(new_n548));
  INV_X1    g347(.A(G71gat), .ZN(new_n549));
  INV_X1    g348(.A(G78gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n544), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G57gat), .ZN(new_n552));
  OR3_X1    g351(.A1(new_n552), .A2(KEYINPUT97), .A3(G64gat), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n548), .A2(new_n546), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n541), .B1(new_n542), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(new_n208), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n542), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(new_n298), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n559), .B2(new_n560), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n534), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n565), .ZN(new_n567));
  INV_X1    g366(.A(new_n534), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n567), .A2(new_n568), .A3(new_n563), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n530), .A2(new_n531), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g370(.A1(new_n449), .A2(new_n571), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n541), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n520), .A2(new_n541), .ZN(new_n574));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(KEYINPUT18), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n484), .B(new_n541), .Z(new_n580));
  XOR2_X1   g379(.A(new_n575), .B(KEYINPUT13), .Z(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n578), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n573), .A2(new_n574), .A3(new_n575), .A4(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n579), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT92), .B(KEYINPUT11), .Z(new_n586));
  XNOR2_X1  g385(.A(G113gat), .B(G141gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G169gat), .B(G197gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(KEYINPUT12), .Z(new_n591));
  NAND2_X1  g390(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n591), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n579), .A2(new_n593), .A3(new_n582), .A4(new_n584), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n555), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n596), .B1(new_n499), .B2(new_n501), .ZN(new_n597));
  INV_X1    g396(.A(G230gat), .ZN(new_n598));
  INV_X1    g397(.A(G233gat), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n555), .B1(new_n498), .B2(new_n496), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G120gat), .B(G148gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(G176gat), .B(G204gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  OAI211_X1 g407(.A(KEYINPUT10), .B(new_n596), .C1(new_n502), .C2(new_n503), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT10), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n597), .B2(new_n602), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n600), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n612), .A2(KEYINPUT102), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT102), .ZN(new_n614));
  AOI211_X1 g413(.A(new_n614), .B(new_n600), .C1(new_n609), .C2(new_n611), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n604), .B(new_n608), .C1(new_n613), .C2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n607), .B1(new_n612), .B2(new_n603), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n595), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n572), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n621), .A2(new_n375), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT103), .B(G1gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(G1324gat));
  INV_X1    g423(.A(new_n621), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n411), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT42), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT104), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT16), .Z(new_n629));
  NOR3_X1   g428(.A1(new_n626), .A2(new_n540), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(G8gat), .B1(new_n626), .B2(new_n627), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n626), .A2(new_n629), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(G1325gat));
  AOI21_X1  g432(.A(G15gat), .B1(new_n625), .B2(new_n283), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n418), .A2(new_n421), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n634), .B1(G15gat), .B2(new_n637), .ZN(G1326gat));
  NOR2_X1   g437(.A1(new_n621), .A2(new_n404), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT43), .B(G22gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(G1327gat));
  NAND2_X1  g440(.A1(new_n515), .A2(new_n526), .ZN(new_n642));
  INV_X1    g441(.A(new_n529), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n515), .A2(new_n526), .A3(new_n529), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR4_X1   g446(.A1(new_n411), .A2(new_n281), .A3(new_n282), .A4(new_n403), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n408), .B1(new_n648), .B2(new_n375), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n649), .A2(new_n447), .B1(new_n422), .B2(new_n445), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n647), .B1(new_n650), .B2(new_n410), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n570), .A3(new_n620), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n652), .A2(G29gat), .A3(new_n375), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT45), .Z(new_n654));
  OR2_X1    g453(.A1(new_n566), .A2(new_n569), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT105), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n620), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT106), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n449), .A2(new_n646), .ZN(new_n661));
  NOR2_X1   g460(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n662));
  NAND2_X1  g461(.A1(KEYINPUT107), .A2(KEYINPUT44), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n661), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n449), .A2(new_n646), .A3(new_n663), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n660), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n412), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(G29gat), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n669), .ZN(G1328gat));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n411), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT108), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n667), .A2(KEYINPUT108), .A3(new_n411), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(G36gat), .A3(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n323), .A2(G36gat), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT46), .B1(new_n652), .B2(new_n676), .ZN(new_n677));
  OR3_X1    g476(.A1(new_n652), .A2(KEYINPUT46), .A3(new_n676), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(G1329gat));
  NAND4_X1  g478(.A1(new_n651), .A2(new_n570), .A3(new_n283), .A4(new_n620), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n680), .A2(G43gat), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT110), .B1(new_n667), .B2(new_n635), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n664), .A2(new_n662), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n666), .B1(new_n651), .B2(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n684), .A2(KEYINPUT110), .A3(new_n635), .A4(new_n659), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G43gat), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n681), .B(KEYINPUT47), .C1(new_n682), .C2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n652), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n688), .A2(KEYINPUT109), .A3(new_n456), .A4(new_n283), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n680), .B2(G43gat), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n456), .B1(new_n667), .B2(new_n635), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n687), .B1(new_n694), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g494(.A1(new_n684), .A2(new_n403), .A3(new_n659), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G50gat), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT48), .B1(new_n697), .B2(KEYINPUT111), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n688), .A2(new_n454), .A3(new_n403), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n697), .B(new_n699), .C1(KEYINPUT111), .C2(KEYINPUT48), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(G1331gat));
  NAND3_X1  g502(.A1(new_n572), .A2(new_n595), .A3(new_n619), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n375), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(new_n552), .ZN(G1332gat));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n323), .ZN(new_n707));
  NOR2_X1   g506(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n708));
  AND2_X1   g507(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(new_n707), .B2(new_n708), .ZN(G1333gat));
  INV_X1    g510(.A(new_n704), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n549), .A3(new_n283), .ZN(new_n713));
  OAI21_X1  g512(.A(G71gat), .B1(new_n704), .B2(new_n636), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1334gat));
  NOR2_X1   g516(.A1(new_n704), .A2(new_n404), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(new_n550), .ZN(G1335gat));
  INV_X1    g518(.A(KEYINPUT51), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n651), .A2(new_n720), .A3(new_n570), .A4(new_n595), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n449), .A2(new_n570), .A3(new_n646), .A4(new_n595), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT51), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n721), .A2(new_n723), .A3(KEYINPUT112), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT112), .B1(new_n721), .B2(new_n723), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n369), .B(new_n412), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n592), .A2(new_n594), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n655), .A2(new_n727), .ZN(new_n728));
  AND4_X1   g527(.A1(new_n412), .A2(new_n684), .A3(new_n619), .A4(new_n728), .ZN(new_n729));
  OAI22_X1  g528(.A1(new_n726), .A2(new_n618), .B1(new_n369), .B2(new_n729), .ZN(G1336gat));
  AOI22_X1  g529(.A1(new_n721), .A2(new_n723), .B1(KEYINPUT113), .B2(new_n722), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n722), .A2(KEYINPUT113), .A3(new_n720), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n323), .A2(G92gat), .A3(new_n618), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n684), .A2(new_n411), .A3(new_n619), .A4(new_n728), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n736), .A2(G92gat), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT52), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(G92gat), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n721), .A2(new_n723), .A3(new_n733), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n742), .ZN(G1337gat));
  OAI211_X1 g542(.A(new_n267), .B(new_n283), .C1(new_n724), .C2(new_n725), .ZN(new_n744));
  AND4_X1   g543(.A1(new_n635), .A2(new_n684), .A3(new_n619), .A4(new_n728), .ZN(new_n745));
  OAI22_X1  g544(.A1(new_n744), .A2(new_n618), .B1(new_n267), .B2(new_n745), .ZN(G1338gat));
  NOR3_X1   g545(.A1(new_n404), .A2(G106gat), .A3(new_n618), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n731), .A2(new_n732), .A3(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n684), .A2(new_n403), .A3(new_n619), .A4(new_n728), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n750), .A2(G106gat), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT53), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT53), .B1(new_n750), .B2(G106gat), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n721), .A2(new_n723), .A3(new_n747), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n752), .A2(new_n758), .ZN(G1339gat));
  NAND3_X1  g558(.A1(new_n609), .A2(new_n611), .A3(new_n600), .ZN(new_n760));
  OAI211_X1 g559(.A(KEYINPUT54), .B(new_n760), .C1(new_n613), .C2(new_n615), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n608), .B1(new_n612), .B2(new_n762), .ZN(new_n763));
  AND3_X1   g562(.A1(new_n761), .A2(KEYINPUT55), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(KEYINPUT55), .B1(new_n761), .B2(new_n763), .ZN(new_n765));
  INV_X1    g564(.A(new_n616), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n575), .B1(new_n573), .B2(new_n574), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n580), .A2(new_n581), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n590), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n594), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n767), .B(new_n772), .C1(new_n530), .C2(new_n531), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n646), .A2(KEYINPUT116), .A3(new_n767), .A4(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n767), .A2(new_n727), .B1(new_n619), .B2(new_n772), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n778), .A2(new_n646), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n656), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n644), .A2(new_n655), .A3(new_n595), .A4(new_n645), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n781), .B1(new_n782), .B2(new_n619), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n571), .A2(KEYINPUT115), .A3(new_n595), .A4(new_n618), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n375), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n648), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n788), .B(KEYINPUT117), .Z(new_n789));
  OAI21_X1  g588(.A(G113gat), .B1(new_n789), .B2(new_n595), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n788), .A2(G113gat), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n595), .B2(new_n791), .ZN(G1340gat));
  OAI21_X1  g591(.A(G120gat), .B1(new_n789), .B2(new_n618), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n788), .A2(G120gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n618), .B2(new_n794), .ZN(G1341gat));
  INV_X1    g594(.A(G127gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n789), .A2(new_n796), .A3(new_n657), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n787), .A2(new_n655), .A3(new_n648), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n797), .B1(new_n796), .B2(new_n798), .ZN(G1342gat));
  OAI21_X1  g598(.A(G134gat), .B1(new_n789), .B2(new_n647), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n788), .A2(G134gat), .A3(new_n647), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT56), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1343gat));
  INV_X1    g602(.A(KEYINPUT121), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n771), .B1(new_n644), .B2(new_n645), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT116), .B1(new_n806), .B2(new_n767), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n773), .A2(new_n774), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n779), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n785), .B1(new_n809), .B2(new_n570), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT57), .B1(new_n810), .B2(new_n404), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n403), .C1(new_n780), .C2(new_n785), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n635), .A2(new_n375), .A3(new_n411), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n811), .A2(new_n727), .A3(new_n813), .A4(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT118), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n815), .A2(new_n816), .A3(new_n327), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n815), .B2(new_n327), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT119), .B1(new_n786), .B2(new_n375), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n778), .A2(new_n646), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n775), .B2(new_n776), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n783), .B(new_n784), .C1(new_n822), .C2(new_n656), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n823), .A2(new_n824), .A3(new_n412), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n635), .A2(new_n404), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n820), .A2(new_n323), .A3(new_n825), .A4(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(G141gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n829), .A3(new_n727), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n805), .B1(new_n819), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n327), .ZN(new_n832));
  XNOR2_X1  g631(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n804), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n827), .A2(G141gat), .A3(new_n595), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n837), .A2(new_n817), .A3(new_n818), .ZN(new_n838));
  OAI211_X1 g637(.A(KEYINPUT121), .B(new_n836), .C1(new_n838), .C2(new_n805), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n835), .A2(new_n839), .ZN(G1344gat));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n841), .B(G148gat), .C1(new_n842), .C2(new_n618), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n823), .A2(KEYINPUT57), .A3(new_n403), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n655), .B1(new_n779), .B2(new_n773), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n782), .A2(new_n619), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n403), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n812), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n823), .A2(KEYINPUT122), .A3(KEYINPUT57), .A4(new_n403), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n846), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n619), .A3(new_n814), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(G148gat), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT123), .B1(new_n854), .B2(KEYINPUT59), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n856));
  AOI211_X1 g655(.A(new_n856), .B(new_n841), .C1(new_n853), .C2(G148gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n843), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n828), .A2(new_n325), .A3(new_n619), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1345gat));
  NOR3_X1   g659(.A1(new_n842), .A2(new_n331), .A3(new_n657), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n828), .A2(new_n655), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n862), .B2(new_n331), .ZN(G1346gat));
  NOR3_X1   g662(.A1(new_n842), .A2(new_n332), .A3(new_n647), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n828), .A2(new_n646), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n332), .ZN(G1347gat));
  NOR2_X1   g665(.A1(new_n786), .A2(new_n412), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n407), .A2(new_n411), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT124), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n233), .A3(new_n727), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n867), .A2(new_n868), .ZN(new_n872));
  OAI21_X1  g671(.A(G169gat), .B1(new_n872), .B2(new_n595), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1348gat));
  AOI21_X1  g673(.A(G176gat), .B1(new_n870), .B2(new_n619), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n872), .A2(new_n232), .A3(new_n618), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(G1349gat));
  NAND3_X1  g676(.A1(new_n870), .A2(new_n655), .A3(new_n241), .ZN(new_n878));
  OAI21_X1  g677(.A(G183gat), .B1(new_n872), .B2(new_n657), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g680(.A1(new_n870), .A2(new_n646), .A3(new_n240), .ZN(new_n882));
  OAI21_X1  g681(.A(G190gat), .B1(new_n872), .B2(new_n647), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n883), .A2(KEYINPUT61), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(KEYINPUT61), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT125), .ZN(G1351gat));
  NOR3_X1   g686(.A1(new_n635), .A2(new_n412), .A3(new_n323), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT126), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n852), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G197gat), .B1(new_n890), .B2(new_n595), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n786), .A2(new_n404), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n888), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n893), .A2(G197gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n891), .B1(new_n595), .B2(new_n894), .ZN(G1352gat));
  AOI21_X1  g694(.A(new_n893), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n896));
  INV_X1    g695(.A(G204gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n897), .A3(new_n619), .ZN(new_n898));
  NOR2_X1   g697(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n899));
  XNOR2_X1  g698(.A(new_n898), .B(new_n899), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n852), .A2(new_n619), .A3(new_n889), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n897), .B2(new_n901), .ZN(G1353gat));
  NAND3_X1  g701(.A1(new_n852), .A2(new_n655), .A3(new_n889), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n903), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT63), .B1(new_n903), .B2(G211gat), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n655), .A2(new_n298), .ZN(new_n906));
  OAI22_X1  g705(.A1(new_n904), .A2(new_n905), .B1(new_n893), .B2(new_n906), .ZN(G1354gat));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n299), .A3(new_n647), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n646), .A3(new_n888), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n299), .B2(new_n909), .ZN(G1355gat));
endmodule


