

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X1 U322 ( .A(n430), .B(n429), .Z(n290) );
  INV_X1 U323 ( .A(KEYINPUT54), .ZN(n450) );
  XNOR2_X1 U324 ( .A(n450), .B(KEYINPUT120), .ZN(n451) );
  XNOR2_X1 U325 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U326 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U327 ( .A(n407), .B(n406), .ZN(n577) );
  NOR2_X1 U328 ( .A1(n456), .A2(n455), .ZN(n566) );
  XNOR2_X1 U329 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U330 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(G127GAT), .B(G120GAT), .Z(n292) );
  XNOR2_X1 U332 ( .A(G15GAT), .B(KEYINPUT84), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n308) );
  XOR2_X1 U334 ( .A(G190GAT), .B(G134GAT), .Z(n294) );
  XNOR2_X1 U335 ( .A(G43GAT), .B(G99GAT), .ZN(n293) );
  XNOR2_X1 U336 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U337 ( .A(n295), .B(G71GAT), .Z(n297) );
  XOR2_X1 U338 ( .A(G113GAT), .B(KEYINPUT0), .Z(n340) );
  XNOR2_X1 U339 ( .A(G169GAT), .B(n340), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U341 ( .A(KEYINPUT20), .B(G176GAT), .Z(n299) );
  NAND2_X1 U342 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U344 ( .A(n301), .B(n300), .Z(n306) );
  XOR2_X1 U345 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n303) );
  XNOR2_X1 U346 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n302) );
  XNOR2_X1 U347 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U348 ( .A(KEYINPUT19), .B(n304), .Z(n446) );
  XNOR2_X1 U349 ( .A(n446), .B(KEYINPUT83), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X2 U351 ( .A(n308), .B(n307), .Z(n528) );
  INV_X1 U352 ( .A(n528), .ZN(n456) );
  XOR2_X1 U353 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n310) );
  XNOR2_X1 U354 ( .A(G148GAT), .B(G204GAT), .ZN(n309) );
  XNOR2_X1 U355 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U356 ( .A(G106GAT), .B(G78GAT), .Z(n402) );
  XOR2_X1 U357 ( .A(n311), .B(n402), .Z(n317) );
  XNOR2_X1 U358 ( .A(G211GAT), .B(KEYINPUT88), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n312), .B(KEYINPUT21), .ZN(n313) );
  XOR2_X1 U360 ( .A(n313), .B(KEYINPUT87), .Z(n315) );
  XNOR2_X1 U361 ( .A(G197GAT), .B(G218GAT), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n445) );
  XOR2_X1 U363 ( .A(G50GAT), .B(G162GAT), .Z(n353) );
  XNOR2_X1 U364 ( .A(n445), .B(n353), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U366 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n319) );
  NAND2_X1 U367 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U369 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U370 ( .A(KEYINPUT3), .B(KEYINPUT89), .Z(n323) );
  XNOR2_X1 U371 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U373 ( .A(G141GAT), .B(n324), .ZN(n348) );
  XOR2_X1 U374 ( .A(G22GAT), .B(n348), .Z(n325) );
  XNOR2_X1 U375 ( .A(n326), .B(n325), .ZN(n470) );
  XOR2_X1 U376 ( .A(KEYINPUT90), .B(KEYINPUT94), .Z(n328) );
  XNOR2_X1 U377 ( .A(G162GAT), .B(KEYINPUT4), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U379 ( .A(KEYINPUT92), .B(KEYINPUT6), .Z(n330) );
  XNOR2_X1 U380 ( .A(KEYINPUT1), .B(KEYINPUT91), .ZN(n329) );
  XNOR2_X1 U381 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U382 ( .A(n332), .B(n331), .Z(n342) );
  INV_X1 U383 ( .A(G134GAT), .ZN(n333) );
  NAND2_X1 U384 ( .A1(G29GAT), .A2(n333), .ZN(n336) );
  INV_X1 U385 ( .A(G29GAT), .ZN(n334) );
  NAND2_X1 U386 ( .A1(n334), .A2(G134GAT), .ZN(n335) );
  NAND2_X1 U387 ( .A1(n336), .A2(n335), .ZN(n350) );
  XOR2_X1 U388 ( .A(G1GAT), .B(G127GAT), .Z(n372) );
  XOR2_X1 U389 ( .A(n350), .B(n372), .Z(n338) );
  NAND2_X1 U390 ( .A1(G225GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U394 ( .A(n343), .B(KEYINPUT5), .Z(n347) );
  XOR2_X1 U395 ( .A(G57GAT), .B(G85GAT), .Z(n345) );
  XNOR2_X1 U396 ( .A(G120GAT), .B(G148GAT), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n345), .B(n344), .ZN(n394) );
  XNOR2_X1 U398 ( .A(n394), .B(KEYINPUT93), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n349) );
  XNOR2_X1 U400 ( .A(n349), .B(n348), .ZN(n468) );
  XNOR2_X1 U401 ( .A(KEYINPUT95), .B(n468), .ZN(n514) );
  XOR2_X1 U402 ( .A(KEYINPUT71), .B(G99GAT), .Z(n401) );
  XNOR2_X1 U403 ( .A(n401), .B(n350), .ZN(n352) );
  AND2_X1 U404 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n352), .B(n351), .ZN(n354) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n362) );
  XOR2_X1 U407 ( .A(KEYINPUT76), .B(G92GAT), .Z(n356) );
  XNOR2_X1 U408 ( .A(G218GAT), .B(G85GAT), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U410 ( .A(KEYINPUT74), .B(KEYINPUT10), .Z(n358) );
  XNOR2_X1 U411 ( .A(G106GAT), .B(KEYINPUT78), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U413 ( .A(n360), .B(n359), .Z(n361) );
  XNOR2_X1 U414 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U415 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n364) );
  XNOR2_X1 U416 ( .A(KEYINPUT75), .B(KEYINPUT77), .ZN(n363) );
  XNOR2_X1 U417 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n366), .B(n365), .ZN(n370) );
  XNOR2_X1 U419 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n367) );
  XNOR2_X1 U420 ( .A(n367), .B(KEYINPUT7), .ZN(n414) );
  XNOR2_X1 U421 ( .A(G36GAT), .B(G190GAT), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n368), .B(KEYINPUT79), .ZN(n440) );
  XNOR2_X1 U423 ( .A(n414), .B(n440), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n541) );
  XNOR2_X1 U425 ( .A(n541), .B(KEYINPUT104), .ZN(n371) );
  XNOR2_X1 U426 ( .A(n371), .B(KEYINPUT36), .ZN(n488) );
  XOR2_X1 U427 ( .A(G71GAT), .B(KEYINPUT13), .Z(n403) );
  XOR2_X1 U428 ( .A(n403), .B(n372), .Z(n374) );
  XNOR2_X1 U429 ( .A(G183GAT), .B(G78GAT), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U431 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n376) );
  NAND2_X1 U432 ( .A1(G231GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U433 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U434 ( .A(n378), .B(n377), .Z(n380) );
  XOR2_X1 U435 ( .A(G15GAT), .B(G22GAT), .Z(n411) );
  XNOR2_X1 U436 ( .A(n411), .B(KEYINPUT12), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n388) );
  XOR2_X1 U438 ( .A(G57GAT), .B(G211GAT), .Z(n382) );
  XNOR2_X1 U439 ( .A(G8GAT), .B(G155GAT), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n386) );
  XOR2_X1 U441 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n384) );
  XNOR2_X1 U442 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U444 ( .A(n386), .B(n385), .Z(n387) );
  XOR2_X1 U445 ( .A(n388), .B(n387), .Z(n580) );
  NAND2_X1 U446 ( .A1(n488), .A2(n580), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n389), .B(KEYINPUT45), .ZN(n391) );
  INV_X1 U448 ( .A(KEYINPUT64), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n391), .B(n390), .ZN(n428) );
  XOR2_X1 U450 ( .A(G64GAT), .B(G92GAT), .Z(n393) );
  XNOR2_X1 U451 ( .A(G176GAT), .B(G204GAT), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n436) );
  XNOR2_X1 U453 ( .A(n394), .B(n436), .ZN(n399) );
  XOR2_X1 U454 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n396) );
  NAND2_X1 U455 ( .A1(G230GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U457 ( .A(n397), .B(KEYINPUT72), .Z(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U459 ( .A(n400), .B(KEYINPUT33), .Z(n407) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n403), .B(KEYINPUT31), .ZN(n404) );
  XOR2_X1 U462 ( .A(G197GAT), .B(G141GAT), .Z(n409) );
  XNOR2_X1 U463 ( .A(G36GAT), .B(G113GAT), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U465 ( .A(n410), .B(G29GAT), .Z(n413) );
  XNOR2_X1 U466 ( .A(n411), .B(G50GAT), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n418) );
  XOR2_X1 U468 ( .A(G169GAT), .B(G8GAT), .Z(n437) );
  XOR2_X1 U469 ( .A(n414), .B(n437), .Z(n416) );
  NAND2_X1 U470 ( .A1(G229GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U471 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U472 ( .A(n418), .B(n417), .Z(n426) );
  XOR2_X1 U473 ( .A(KEYINPUT70), .B(KEYINPUT68), .Z(n420) );
  XNOR2_X1 U474 ( .A(G1GAT), .B(KEYINPUT69), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U476 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n422) );
  XNOR2_X1 U477 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U480 ( .A(n426), .B(n425), .Z(n574) );
  NOR2_X1 U481 ( .A1(n577), .A2(n574), .ZN(n427) );
  NAND2_X1 U482 ( .A1(n428), .A2(n427), .ZN(n434) );
  INV_X1 U483 ( .A(n541), .ZN(n557) );
  INV_X1 U484 ( .A(n580), .ZN(n554) );
  NAND2_X1 U485 ( .A1(n557), .A2(n554), .ZN(n431) );
  XNOR2_X1 U486 ( .A(KEYINPUT46), .B(KEYINPUT111), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n577), .B(KEYINPUT41), .ZN(n550) );
  INV_X1 U488 ( .A(n574), .ZN(n547) );
  NOR2_X1 U489 ( .A1(n550), .A2(n547), .ZN(n429) );
  NOR2_X1 U490 ( .A1(n431), .A2(n290), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n432), .B(KEYINPUT47), .ZN(n433) );
  NAND2_X1 U492 ( .A1(n434), .A2(n433), .ZN(n435) );
  XOR2_X1 U493 ( .A(KEYINPUT48), .B(n435), .Z(n527) );
  XOR2_X1 U494 ( .A(KEYINPUT96), .B(KEYINPUT98), .Z(n439) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U496 ( .A(n439), .B(n438), .ZN(n444) );
  XOR2_X1 U497 ( .A(n440), .B(KEYINPUT97), .Z(n442) );
  NAND2_X1 U498 ( .A1(G226GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U500 ( .A(n444), .B(n443), .Z(n448) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U502 ( .A(n448), .B(n447), .ZN(n516) );
  XNOR2_X1 U503 ( .A(n516), .B(KEYINPUT119), .ZN(n449) );
  NOR2_X1 U504 ( .A1(n527), .A2(n449), .ZN(n452) );
  NOR2_X1 U505 ( .A1(n514), .A2(n453), .ZN(n571) );
  AND2_X1 U506 ( .A1(n470), .A2(n571), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n454), .B(KEYINPUT55), .ZN(n455) );
  NAND2_X1 U508 ( .A1(n566), .A2(n541), .ZN(n460) );
  XOR2_X1 U509 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n458) );
  INV_X1 U510 ( .A(G190GAT), .ZN(n457) );
  XOR2_X1 U511 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n480) );
  NOR2_X1 U512 ( .A1(n547), .A2(n577), .ZN(n492) );
  NOR2_X1 U513 ( .A1(n470), .A2(n528), .ZN(n461) );
  XNOR2_X1 U514 ( .A(n461), .B(KEYINPUT26), .ZN(n572) );
  XNOR2_X1 U515 ( .A(n516), .B(KEYINPUT27), .ZN(n472) );
  NAND2_X1 U516 ( .A1(n572), .A2(n472), .ZN(n462) );
  XNOR2_X1 U517 ( .A(KEYINPUT100), .B(n462), .ZN(n466) );
  NAND2_X1 U518 ( .A1(n528), .A2(n516), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n470), .A2(n463), .ZN(n464) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n464), .Z(n465) );
  NAND2_X1 U521 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U523 ( .A(n469), .B(KEYINPUT101), .ZN(n476) );
  XNOR2_X1 U524 ( .A(n470), .B(KEYINPUT65), .ZN(n471) );
  XNOR2_X1 U525 ( .A(n471), .B(KEYINPUT28), .ZN(n531) );
  NAND2_X1 U526 ( .A1(n514), .A2(n472), .ZN(n526) );
  NOR2_X1 U527 ( .A1(n531), .A2(n526), .ZN(n473) );
  XNOR2_X1 U528 ( .A(KEYINPUT99), .B(n473), .ZN(n474) );
  NOR2_X1 U529 ( .A1(n474), .A2(n528), .ZN(n475) );
  NOR2_X1 U530 ( .A1(n476), .A2(n475), .ZN(n489) );
  NOR2_X1 U531 ( .A1(n541), .A2(n554), .ZN(n477) );
  XOR2_X1 U532 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  NOR2_X1 U533 ( .A1(n489), .A2(n478), .ZN(n502) );
  AND2_X1 U534 ( .A1(n492), .A2(n502), .ZN(n486) );
  NAND2_X1 U535 ( .A1(n486), .A2(n514), .ZN(n479) );
  XNOR2_X1 U536 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U537 ( .A(G1GAT), .B(n481), .Z(G1324GAT) );
  XOR2_X1 U538 ( .A(G8GAT), .B(KEYINPUT103), .Z(n483) );
  NAND2_X1 U539 ( .A1(n486), .A2(n516), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(G1325GAT) );
  XOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT35), .Z(n485) );
  NAND2_X1 U542 ( .A1(n486), .A2(n528), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NAND2_X1 U544 ( .A1(n486), .A2(n531), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U546 ( .A1(n580), .A2(n489), .ZN(n490) );
  NAND2_X1 U547 ( .A1(n488), .A2(n490), .ZN(n491) );
  XOR2_X1 U548 ( .A(n491), .B(KEYINPUT37), .Z(n513) );
  INV_X1 U549 ( .A(n513), .ZN(n493) );
  NAND2_X1 U550 ( .A1(n493), .A2(n492), .ZN(n494) );
  XOR2_X1 U551 ( .A(KEYINPUT38), .B(n494), .Z(n500) );
  NAND2_X1 U552 ( .A1(n514), .A2(n500), .ZN(n496) );
  XOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .Z(n495) );
  XNOR2_X1 U554 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NAND2_X1 U555 ( .A1(n500), .A2(n516), .ZN(n497) );
  XNOR2_X1 U556 ( .A(n497), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U557 ( .A1(n500), .A2(n528), .ZN(n498) );
  XNOR2_X1 U558 ( .A(n498), .B(KEYINPUT40), .ZN(n499) );
  XNOR2_X1 U559 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n500), .A2(n531), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n501), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U562 ( .A(KEYINPUT105), .B(n550), .ZN(n563) );
  NAND2_X1 U563 ( .A1(n547), .A2(n563), .ZN(n512) );
  INV_X1 U564 ( .A(n502), .ZN(n503) );
  NOR2_X1 U565 ( .A1(n512), .A2(n503), .ZN(n509) );
  NAND2_X1 U566 ( .A1(n509), .A2(n514), .ZN(n504) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(n504), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n509), .A2(n516), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U571 ( .A1(n509), .A2(n528), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(KEYINPUT106), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U575 ( .A1(n509), .A2(n531), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  NOR2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n521), .A2(n514), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n515), .ZN(G1336GAT) );
  XOR2_X1 U580 ( .A(G92GAT), .B(KEYINPUT107), .Z(n518) );
  NAND2_X1 U581 ( .A1(n521), .A2(n516), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n521), .A2(n528), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(KEYINPUT108), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(n520), .ZN(G1338GAT) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(KEYINPUT109), .ZN(n525) );
  XOR2_X1 U587 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n523) );
  NAND2_X1 U588 ( .A1(n521), .A2(n531), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1339GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n533) );
  NOR2_X1 U592 ( .A1(n527), .A2(n526), .ZN(n546) );
  NAND2_X1 U593 ( .A1(n528), .A2(n546), .ZN(n529) );
  XNOR2_X1 U594 ( .A(KEYINPUT112), .B(n529), .ZN(n530) );
  NOR2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n542), .A2(n574), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U600 ( .A1(n542), .A2(n563), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n538) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT115), .Z(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  NAND2_X1 U604 ( .A1(n542), .A2(n580), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n539), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT51), .B(KEYINPUT117), .Z(n544) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U610 ( .A(G134GAT), .B(n545), .Z(G1343GAT) );
  NAND2_X1 U611 ( .A1(n546), .A2(n572), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n547), .A2(n556), .ZN(n548) );
  XOR2_X1 U613 ( .A(G141GAT), .B(n548), .Z(n549) );
  XNOR2_X1 U614 ( .A(KEYINPUT118), .B(n549), .ZN(G1344GAT) );
  NOR2_X1 U615 ( .A1(n550), .A2(n556), .ZN(n552) );
  XNOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U619 ( .A1(n554), .A2(n556), .ZN(n555) );
  XOR2_X1 U620 ( .A(G155GAT), .B(n555), .Z(G1346GAT) );
  NOR2_X1 U621 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  NAND2_X1 U623 ( .A1(n566), .A2(n574), .ZN(n559) );
  XNOR2_X1 U624 ( .A(G169GAT), .B(n559), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n561) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(KEYINPUT56), .B(n562), .Z(n565) );
  NAND2_X1 U629 ( .A1(n563), .A2(n566), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1349GAT) );
  XOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT123), .Z(n568) );
  NAND2_X1 U632 ( .A1(n566), .A2(n580), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1350GAT) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT126), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT60), .B(n570), .Z(n576) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(KEYINPUT125), .ZN(n582) );
  NAND2_X1 U639 ( .A1(n582), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  NAND2_X1 U642 ( .A1(n582), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n582), .A2(n580), .ZN(n581) );
  XNOR2_X1 U645 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U646 ( .A1(n488), .A2(n582), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

