//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n202));
  XNOR2_X1  g001(.A(G113gat), .B(G141gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT11), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n203), .A2(KEYINPUT11), .ZN(new_n206));
  OAI21_X1  g005(.A(G169gat), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n203), .A2(KEYINPUT11), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(new_n204), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n207), .A2(G197gat), .A3(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(G197gat), .B1(new_n207), .B2(new_n210), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n202), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G197gat), .ZN(new_n214));
  NOR3_X1   g013(.A1(new_n205), .A2(G169gat), .A3(new_n206), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n209), .B1(new_n208), .B2(new_n204), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n207), .A2(G197gat), .A3(new_n210), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(KEYINPUT12), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G43gat), .A2(G50gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(G43gat), .A2(G50gat), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT15), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G29gat), .ZN(new_n226));
  INV_X1    g025(.A(G36gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT14), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT14), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G29gat), .B2(G36gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n230), .A3(KEYINPUT87), .ZN(new_n231));
  NAND2_X1  g030(.A1(G29gat), .A2(G36gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT87), .B1(new_n228), .B2(new_n230), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n225), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT88), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT88), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n237), .B(new_n225), .C1(new_n233), .C2(new_n234), .ZN(new_n238));
  INV_X1    g037(.A(new_n223), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT15), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(new_n221), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n224), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n232), .A2(KEYINPUT89), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT89), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(G29gat), .A3(G36gat), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n228), .A2(new_n243), .A3(new_n230), .A4(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n236), .A2(new_n238), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G8gat), .ZN(new_n250));
  INV_X1    g049(.A(G22gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G15gat), .ZN(new_n252));
  INV_X1    g051(.A(G15gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(G22gat), .ZN(new_n254));
  INV_X1    g053(.A(G1gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT16), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n252), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT90), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n254), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(new_n255), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT90), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n252), .A2(new_n254), .A3(new_n256), .A4(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT92), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n259), .A2(new_n255), .B1(new_n264), .B2(G8gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT91), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n257), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n252), .A2(new_n254), .A3(new_n256), .A4(KEYINPUT91), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n250), .B1(new_n263), .B2(new_n269), .ZN(new_n270));
  AND4_X1   g069(.A1(new_n264), .A2(new_n265), .A3(new_n267), .A4(new_n268), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n249), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n260), .A3(new_n262), .ZN(new_n274));
  OAI21_X1  g073(.A(G8gat), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n247), .B1(new_n235), .B2(KEYINPUT88), .ZN(new_n276));
  INV_X1    g075(.A(new_n271), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .A4(new_n238), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G229gat), .A2(G233gat), .ZN(new_n280));
  XOR2_X1   g079(.A(new_n280), .B(KEYINPUT13), .Z(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n275), .A2(new_n277), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT17), .B1(new_n276), .B2(new_n238), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n236), .A2(KEYINPUT17), .A3(new_n238), .A4(new_n248), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT93), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n276), .A2(KEYINPUT93), .A3(KEYINPUT17), .A4(new_n238), .ZN(new_n288));
  AOI211_X1 g087(.A(new_n283), .B(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n236), .A2(new_n238), .A3(new_n248), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n263), .A2(new_n269), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n271), .B1(new_n291), .B2(G8gat), .ZN(new_n292));
  OAI211_X1 g091(.A(KEYINPUT18), .B(new_n280), .C1(new_n290), .C2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n282), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n287), .A2(new_n288), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n284), .A2(new_n283), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n272), .A2(new_n280), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT18), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n220), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n220), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n282), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT18), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(new_n289), .B2(new_n298), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT94), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n220), .B1(new_n279), .B2(new_n281), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n289), .B2(new_n293), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT94), .ZN(new_n311));
  NOR3_X1   g110(.A1(new_n310), .A2(new_n300), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n301), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT95), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n305), .A2(KEYINPUT94), .A3(new_n307), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n311), .B1(new_n310), .B2(new_n300), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT95), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n318), .A3(new_n301), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n321));
  INV_X1    g120(.A(G183gat), .ZN(new_n322));
  INV_X1    g121(.A(G190gat), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G176gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n209), .A2(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n329));
  NOR2_X1   g128(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT23), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n333), .A2(KEYINPUT25), .ZN(new_n334));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT67), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n326), .A2(new_n331), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n331), .A2(new_n333), .A3(new_n335), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT65), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n325), .B(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n324), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n342));
  OAI21_X1  g141(.A(new_n337), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT26), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n335), .B1(new_n332), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT68), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n345), .A2(new_n346), .B1(new_n344), .B2(new_n332), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(new_n346), .B2(new_n345), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT27), .B(G183gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n323), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n350), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n348), .B(new_n351), .C1(KEYINPUT28), .C2(new_n350), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G226gat), .ZN(new_n354));
  INV_X1    g153(.A(G233gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT29), .B1(new_n343), .B2(new_n352), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n357), .B1(new_n358), .B2(new_n356), .ZN(new_n359));
  XNOR2_X1  g158(.A(G211gat), .B(G218gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT75), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT74), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G197gat), .B(G204gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(new_n363), .B2(new_n362), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n361), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT75), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n360), .B(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n366), .A2(new_n364), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(KEYINPUT76), .A3(new_n371), .ZN(new_n372));
  OR3_X1    g171(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT76), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n359), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n357), .ZN(new_n376));
  XOR2_X1   g175(.A(KEYINPUT77), .B(KEYINPUT29), .Z(new_n377));
  AOI21_X1  g176(.A(new_n356), .B1(new_n353), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n374), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(G36gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT78), .B(G8gat), .ZN(new_n382));
  XOR2_X1   g181(.A(new_n381), .B(new_n382), .Z(new_n383));
  NAND3_X1  g182(.A1(new_n375), .A2(new_n379), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n375), .A2(new_n379), .A3(KEYINPUT79), .A4(new_n383), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT30), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n375), .A2(new_n379), .ZN(new_n389));
  INV_X1    g188(.A(new_n383), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT30), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(new_n384), .ZN(new_n393));
  OR2_X1    g192(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT70), .B(G120gat), .ZN(new_n395));
  MUX2_X1   g194(.A(G120gat), .B(new_n395), .S(G113gat), .Z(new_n396));
  INV_X1    g195(.A(G127gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G134gat), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n397), .A2(G134gat), .ZN(new_n399));
  OR2_X1    g198(.A1(KEYINPUT71), .A2(KEYINPUT1), .ZN(new_n400));
  NAND2_X1  g199(.A1(KEYINPUT71), .A2(KEYINPUT1), .ZN(new_n401));
  AND4_X1   g200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(KEYINPUT69), .B(G134gat), .Z(new_n403));
  OAI21_X1  g202(.A(new_n398), .B1(new_n403), .B2(new_n397), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT1), .ZN(new_n405));
  INV_X1    g204(.A(G113gat), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n406), .A2(G120gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(G120gat), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI22_X1  g208(.A1(new_n396), .A2(new_n402), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n353), .A2(new_n410), .ZN(new_n411));
  AND2_X1   g210(.A1(G227gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n410), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n343), .A2(new_n413), .A3(new_n352), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT32), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(G71gat), .B(G99gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT72), .ZN(new_n420));
  XOR2_X1   g219(.A(G15gat), .B(G43gat), .Z(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n422), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n415), .B(KEYINPUT32), .C1(new_n417), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n412), .B1(new_n411), .B2(new_n414), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n427), .A2(KEYINPUT34), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(KEYINPUT34), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT73), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n426), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n423), .A2(new_n428), .A3(new_n429), .A4(new_n425), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n426), .A2(new_n430), .A3(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n374), .ZN(new_n438));
  INV_X1    g237(.A(new_n377), .ZN(new_n439));
  XNOR2_X1  g238(.A(G141gat), .B(G148gat), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT2), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n441), .B1(G155gat), .B2(G162gat), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT80), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(G155gat), .B(G162gat), .Z(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XOR2_X1   g244(.A(KEYINPUT81), .B(KEYINPUT3), .Z(new_n446));
  AOI21_X1  g245(.A(new_n439), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n438), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT29), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n372), .A2(new_n373), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT3), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n445), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g251(.A(G228gat), .B(G233gat), .C1(new_n448), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G228gat), .A2(G233gat), .ZN(new_n454));
  INV_X1    g253(.A(new_n446), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n367), .A2(new_n371), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(new_n377), .ZN(new_n457));
  OAI221_X1 g256(.A(new_n454), .B1(new_n457), .B2(new_n445), .C1(new_n438), .C2(new_n447), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G78gat), .B(G106gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(KEYINPUT31), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n461), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n453), .A2(new_n458), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(G22gat), .B(G50gat), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n462), .A2(new_n466), .A3(new_n464), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n394), .A2(new_n437), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G1gat), .B(G29gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT0), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(G57gat), .ZN(new_n474));
  INV_X1    g273(.A(G85gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n445), .B(new_n410), .ZN(new_n477));
  NAND2_X1  g276(.A1(G225gat), .A2(G233gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(KEYINPUT83), .B(KEYINPUT5), .Z(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n445), .A2(new_n410), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n445), .A2(new_n446), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n485), .B(new_n413), .C1(new_n451), .C2(new_n445), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n478), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n484), .A2(new_n478), .A3(new_n486), .A4(new_n488), .ZN(new_n491));
  AOI211_X1 g290(.A(new_n476), .B(new_n482), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n482), .B1(new_n490), .B2(new_n491), .ZN(new_n494));
  INV_X1    g293(.A(new_n476), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(KEYINPUT84), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n498), .A2(new_n499), .B1(KEYINPUT6), .B2(new_n492), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT35), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n470), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n431), .A2(new_n434), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n388), .A2(new_n393), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n492), .A2(KEYINPUT6), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(new_n496), .B2(new_n492), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n503), .A2(new_n504), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n471), .A2(new_n502), .B1(new_n508), .B2(new_n501), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n470), .B1(new_n500), .B2(new_n394), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT40), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n478), .B1(new_n484), .B2(new_n486), .ZN(new_n512));
  XOR2_X1   g311(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n513));
  AOI21_X1  g312(.A(new_n495), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT39), .B1(new_n477), .B2(new_n479), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n492), .B1(new_n511), .B2(new_n516), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n516), .A2(new_n511), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n517), .B(new_n518), .C1(new_n388), .C2(new_n393), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT37), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n389), .A2(new_n520), .ZN(new_n521));
  OR3_X1    g320(.A1(new_n376), .A2(new_n378), .A3(new_n374), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT86), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n359), .A2(new_n374), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT37), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n522), .A2(KEYINPUT86), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n521), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n383), .A2(KEYINPUT38), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND3_X1   g328(.A1(new_n375), .A2(new_n379), .A3(KEYINPUT37), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT37), .B1(new_n375), .B2(new_n379), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n390), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT38), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n386), .A2(new_n387), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n506), .B(new_n535), .C1(new_n492), .C2(new_n496), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n519), .B(new_n503), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT36), .B1(new_n431), .B2(new_n434), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n538), .B1(new_n437), .B2(KEYINPUT36), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n510), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n320), .B1(new_n509), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT21), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(G57gat), .B2(G64gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(G71gat), .B(G78gat), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G57gat), .ZN(new_n547));
  OAI21_X1  g346(.A(G64gat), .B1(new_n547), .B2(KEYINPUT96), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT96), .ZN(new_n549));
  INV_X1    g348(.A(G64gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n550), .A3(G57gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G71gat), .ZN(new_n553));
  INV_X1    g352(.A(G78gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT97), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n552), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n552), .B2(new_n557), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n546), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n292), .B1(new_n542), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G183gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n564));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n563), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n542), .ZN(new_n568));
  XOR2_X1   g367(.A(G127gat), .B(G155gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G211gat), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n567), .A2(new_n571), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(KEYINPUT41), .ZN(new_n576));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(G99gat), .A2(G106gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT100), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT7), .ZN(new_n584));
  NAND3_X1  g383(.A1(KEYINPUT98), .A2(G85gat), .A3(G92gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n582), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n475), .ZN(new_n588));
  INV_X1    g387(.A(G92gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT8), .ZN(new_n593));
  NAND4_X1  g392(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT100), .B1(new_n580), .B2(new_n581), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n586), .A2(new_n591), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n596), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n599));
  INV_X1    g398(.A(G99gat), .ZN(new_n600));
  INV_X1    g399(.A(G106gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(new_n583), .A3(new_n592), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n585), .A2(new_n584), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n598), .B1(new_n599), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n597), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n284), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n295), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n249), .A2(new_n607), .B1(KEYINPUT41), .B2(new_n575), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n611), .A2(new_n612), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n579), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(new_n578), .A3(new_n613), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n574), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n544), .A2(new_n545), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n552), .A2(new_n557), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT97), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n552), .A2(new_n557), .A3(new_n558), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n622), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n607), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n561), .A2(new_n606), .A3(new_n597), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n607), .A2(KEYINPUT10), .A3(new_n626), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n631), .B1(new_n630), .B2(new_n632), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n621), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n627), .A2(new_n628), .ZN(new_n637));
  INV_X1    g436(.A(new_n621), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G176gat), .ZN(new_n641));
  INV_X1    g440(.A(G204gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n636), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n630), .A2(new_n632), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n621), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n639), .ZN(new_n647));
  INV_X1    g446(.A(new_n643), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n620), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n541), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n498), .A2(new_n499), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n506), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n255), .ZN(G1324gat));
  NOR2_X1   g455(.A1(new_n652), .A2(new_n505), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT102), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT16), .B(G8gat), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n658), .A2(G8gat), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n658), .B2(new_n659), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(G1325gat));
  OAI21_X1  g463(.A(G15gat), .B1(new_n652), .B2(new_n539), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n504), .A2(new_n253), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n665), .B1(new_n652), .B2(new_n666), .ZN(G1326gat));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n503), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT43), .B(G22gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  INV_X1    g469(.A(new_n574), .ZN(new_n671));
  INV_X1    g470(.A(new_n619), .ZN(new_n672));
  INV_X1    g471(.A(new_n650), .ZN(new_n673));
  AND4_X1   g472(.A1(new_n541), .A2(new_n671), .A3(new_n672), .A4(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n226), .A3(new_n500), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT45), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n619), .B1(new_n509), .B2(new_n540), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n313), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n574), .A2(new_n682), .A3(new_n650), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G29gat), .B1(new_n684), .B2(new_n654), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n676), .A2(new_n685), .ZN(G1328gat));
  NAND3_X1  g485(.A1(new_n674), .A2(new_n227), .A3(new_n394), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT46), .Z(new_n688));
  OAI21_X1  g487(.A(G36gat), .B1(new_n684), .B2(new_n505), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1329gat));
  INV_X1    g489(.A(new_n539), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n677), .A2(new_n678), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n678), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n691), .B(new_n683), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G43gat), .ZN(new_n695));
  NOR2_X1   g494(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n696));
  INV_X1    g495(.A(new_n504), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(G43gat), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n696), .B1(new_n674), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(KEYINPUT103), .A2(KEYINPUT47), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1330gat));
  INV_X1    g501(.A(G50gat), .ZN(new_n703));
  OAI211_X1 g502(.A(new_n470), .B(new_n683), .C1(new_n692), .C2(new_n693), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n705), .B2(new_n704), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n674), .A2(new_n703), .A3(new_n470), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n704), .A2(G50gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n709), .B1(new_n712), .B2(new_n708), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(G1331gat));
  NAND2_X1  g513(.A1(new_n682), .A2(new_n650), .ZN(new_n715));
  AOI211_X1 g514(.A(new_n620), .B(new_n715), .C1(new_n509), .C2(new_n540), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n500), .B(KEYINPUT105), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n394), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT49), .B(G64gat), .Z(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n720), .B2(new_n722), .ZN(G1333gat));
  AOI21_X1  g522(.A(new_n553), .B1(new_n716), .B2(new_n691), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n697), .A2(G71gat), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n716), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n716), .A2(new_n470), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g528(.A1(new_n588), .A2(new_n590), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n574), .A2(new_n313), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n650), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n732), .B1(new_n679), .B2(new_n680), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n730), .B1(new_n734), .B2(new_n654), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n510), .A2(new_n537), .A3(new_n539), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n505), .A2(new_n507), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n468), .A2(new_n504), .A3(new_n469), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n501), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n654), .A2(KEYINPUT35), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n503), .A2(new_n436), .A3(new_n505), .A4(new_n435), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n672), .B(new_n731), .C1(new_n736), .C2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n677), .A2(KEYINPUT51), .A3(new_n731), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n677), .A2(KEYINPUT106), .A3(KEYINPUT51), .A4(new_n731), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n654), .A2(new_n730), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n748), .A2(new_n650), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n751), .ZN(G1336gat));
  AOI21_X1  g551(.A(new_n589), .B1(new_n733), .B2(new_n394), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n745), .A2(new_n746), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n505), .A2(G92gat), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n754), .A2(new_n650), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT52), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n732), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n394), .B(new_n758), .C1(new_n692), .C2(new_n693), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT52), .B1(new_n759), .B2(G92gat), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n748), .A2(new_n650), .A3(new_n749), .A4(new_n755), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n760), .A2(KEYINPUT107), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT107), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(G1337gat));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n504), .A3(new_n650), .A4(new_n749), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n600), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n733), .A2(G99gat), .A3(new_n691), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT108), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n766), .A2(new_n770), .A3(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1338gat));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n733), .A2(new_n470), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n775), .B2(new_n601), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n503), .A2(G106gat), .A3(new_n673), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n748), .A2(new_n749), .A3(new_n777), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n774), .A2(G106gat), .B1(new_n754), .B2(new_n777), .ZN(new_n779));
  OAI22_X1  g578(.A1(new_n776), .A2(new_n778), .B1(new_n779), .B2(new_n773), .ZN(G1339gat));
  NAND2_X1  g579(.A1(new_n651), .A2(new_n682), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n279), .A2(new_n281), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT110), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n782), .B(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n280), .B1(new_n297), .B2(new_n272), .ZN(new_n785));
  OAI22_X1  g584(.A1(new_n784), .A2(new_n785), .B1(new_n211), .B2(new_n212), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n317), .A2(new_n786), .A3(new_n650), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n645), .A2(KEYINPUT101), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n638), .B1(new_n789), .B2(new_n633), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n630), .A2(new_n638), .A3(new_n632), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT54), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n788), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n792), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n636), .A2(KEYINPUT109), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n646), .A2(KEYINPUT54), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n643), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n793), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n793), .A2(new_n795), .A3(KEYINPUT55), .A4(new_n797), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n800), .A2(new_n644), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n787), .B1(new_n802), .B2(new_n682), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n317), .A2(new_n786), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT111), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n317), .A2(new_n786), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n802), .A2(new_n619), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n619), .A2(new_n803), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n781), .B1(new_n810), .B2(new_n574), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n717), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n741), .ZN(new_n813));
  AOI21_X1  g612(.A(G113gat), .B1(new_n813), .B2(new_n313), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n808), .A2(new_n809), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n801), .A2(new_n644), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n817), .A2(new_n313), .A3(new_n800), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n672), .B1(new_n818), .B2(new_n787), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n671), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n738), .B1(new_n820), .B2(new_n781), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n500), .A2(new_n505), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n320), .A2(new_n406), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n814), .B1(new_n824), .B2(new_n825), .ZN(G1340gat));
  INV_X1    g625(.A(new_n824), .ZN(new_n827));
  OAI21_X1  g626(.A(G120gat), .B1(new_n827), .B2(new_n673), .ZN(new_n828));
  INV_X1    g627(.A(new_n813), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n650), .A2(new_n395), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT112), .Z(new_n831));
  OAI21_X1  g630(.A(new_n828), .B1(new_n829), .B2(new_n831), .ZN(G1341gat));
  OAI21_X1  g631(.A(G127gat), .B1(new_n827), .B2(new_n671), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n397), .A3(new_n574), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1342gat));
  INV_X1    g634(.A(new_n403), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n813), .A2(new_n836), .A3(new_n672), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(KEYINPUT56), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT113), .Z(new_n839));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n672), .ZN(new_n840));
  AOI22_X1  g639(.A1(G134gat), .A2(new_n840), .B1(new_n837), .B2(KEYINPUT56), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(G1343gat));
  NAND2_X1  g641(.A1(new_n314), .A2(new_n319), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n691), .A2(new_n822), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n503), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT114), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n800), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n798), .A2(KEYINPUT114), .A3(new_n799), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n816), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n843), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n672), .B1(new_n852), .B2(new_n787), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n671), .B1(new_n853), .B2(new_n815), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n847), .B1(new_n854), .B2(new_n781), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT57), .B1(new_n811), .B2(new_n470), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n843), .B(new_n844), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT116), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n503), .B1(new_n820), .B2(new_n781), .ZN(new_n859));
  INV_X1    g658(.A(new_n781), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n808), .A2(new_n809), .ZN(new_n861));
  INV_X1    g660(.A(new_n787), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n862), .B1(new_n851), .B2(new_n843), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n863), .B2(new_n672), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n860), .B1(new_n864), .B2(new_n671), .ZN(new_n865));
  OAI22_X1  g664(.A1(new_n859), .A2(KEYINPUT57), .B1(new_n865), .B2(new_n847), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n843), .A4(new_n844), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n858), .A2(G141gat), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n812), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n811), .A2(KEYINPUT115), .A3(new_n717), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n691), .A2(new_n503), .A3(new_n394), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n320), .A2(G141gat), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n871), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n869), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(G141gat), .ZN(new_n880));
  INV_X1    g679(.A(new_n844), .ZN(new_n881));
  INV_X1    g680(.A(new_n850), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT114), .B1(new_n798), .B2(new_n799), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n817), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n787), .B1(new_n320), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n619), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n574), .B1(new_n886), .B2(new_n861), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n846), .B1(new_n887), .B2(new_n860), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n811), .A2(new_n470), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n845), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n881), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n880), .B1(new_n891), .B2(new_n313), .ZN(new_n892));
  INV_X1    g691(.A(new_n875), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT58), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT117), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n880), .B1(new_n857), .B2(KEYINPUT116), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n877), .B1(new_n897), .B2(new_n868), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n844), .B1(new_n855), .B2(new_n856), .ZN(new_n899));
  OAI21_X1  g698(.A(G141gat), .B1(new_n899), .B2(new_n682), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n876), .B1(new_n900), .B2(new_n875), .ZN(new_n901));
  OAI21_X1  g700(.A(KEYINPUT117), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n896), .A2(new_n902), .ZN(G1344gat));
  INV_X1    g702(.A(G148gat), .ZN(new_n904));
  AOI211_X1 g703(.A(KEYINPUT59), .B(new_n904), .C1(new_n891), .C2(new_n650), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n843), .A2(new_n620), .A3(new_n650), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n845), .B(new_n470), .C1(new_n887), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n889), .A2(KEYINPUT57), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n908), .A2(new_n650), .A3(new_n844), .A4(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n906), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n871), .A2(new_n873), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n872), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n650), .A2(new_n904), .ZN(new_n914));
  OAI22_X1  g713(.A1(new_n905), .A2(new_n911), .B1(new_n913), .B2(new_n914), .ZN(G1345gat));
  NAND3_X1  g714(.A1(new_n912), .A2(new_n574), .A3(new_n872), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(G155gat), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n574), .A2(G155gat), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n918), .A2(new_n919), .B1(new_n891), .B2(new_n920), .ZN(G1346gat));
  NOR2_X1   g720(.A1(new_n619), .A2(G162gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n912), .A2(new_n872), .A3(new_n922), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT119), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n891), .A2(KEYINPUT120), .A3(new_n672), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n899), .B2(new_n619), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n925), .A2(new_n927), .A3(G162gat), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n924), .A2(new_n928), .ZN(G1347gat));
  AOI21_X1  g728(.A(new_n500), .B1(new_n820), .B2(new_n781), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n437), .A2(new_n470), .A3(new_n505), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n209), .A3(new_n313), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT121), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n717), .A2(new_n505), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n821), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(G169gat), .B1(new_n936), .B2(new_n320), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(G1348gat));
  NAND3_X1  g737(.A1(new_n932), .A2(new_n327), .A3(new_n650), .ZN(new_n939));
  OAI21_X1  g738(.A(G176gat), .B1(new_n936), .B2(new_n673), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1349gat));
  AND2_X1   g740(.A1(new_n574), .A2(new_n349), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n943));
  AOI22_X1  g742(.A1(new_n932), .A2(new_n942), .B1(new_n943), .B2(KEYINPUT60), .ZN(new_n944));
  OAI21_X1  g743(.A(KEYINPUT122), .B1(new_n936), .B2(new_n671), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(G183gat), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n936), .A2(KEYINPUT122), .A3(new_n671), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n944), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OR2_X1    g747(.A1(new_n943), .A2(KEYINPUT60), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n948), .B(new_n949), .ZN(G1350gat));
  OAI21_X1  g749(.A(G190gat), .B1(new_n936), .B2(new_n619), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT61), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n932), .A2(new_n323), .A3(new_n672), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(G1351gat));
  NAND3_X1  g753(.A1(new_n539), .A2(new_n470), .A3(new_n394), .ZN(new_n955));
  XOR2_X1   g754(.A(new_n955), .B(KEYINPUT124), .Z(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n930), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n956), .A2(new_n930), .A3(KEYINPUT125), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g760(.A(G197gat), .B1(new_n961), .B2(new_n313), .ZN(new_n962));
  NOR3_X1   g761(.A1(new_n717), .A2(new_n691), .A3(new_n505), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n908), .A2(new_n909), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n320), .A2(new_n214), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G1352gat));
  NAND4_X1  g765(.A1(new_n956), .A2(new_n930), .A3(new_n642), .A4(new_n650), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT62), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n967), .A2(KEYINPUT62), .ZN(new_n969));
  AND4_X1   g768(.A1(new_n650), .A2(new_n908), .A3(new_n909), .A4(new_n963), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n968), .B(new_n969), .C1(new_n970), .C2(new_n642), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n971), .B(new_n972), .ZN(G1353gat));
  NAND2_X1  g772(.A1(new_n964), .A2(new_n574), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G211gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT63), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n671), .A2(G211gat), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n960), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT127), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT63), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n974), .A2(new_n980), .A3(G211gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n976), .A2(new_n979), .A3(new_n981), .ZN(G1354gat));
  AOI21_X1  g781(.A(G218gat), .B1(new_n961), .B2(new_n672), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n672), .A2(G218gat), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(new_n964), .B2(new_n984), .ZN(G1355gat));
endmodule


