//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n525, new_n526, new_n527, new_n528,
    new_n531, new_n532, new_n533, new_n534, new_n537, new_n538, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n584, new_n585, new_n588, new_n590, new_n591,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1125;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G219), .A3(G220), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  XOR2_X1   g029(.A(G325), .B(KEYINPUT67), .Z(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(new_n452), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n463), .A2(G137), .B1(G101), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n462), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n463), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n462), .A2(new_n464), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  INV_X1    g054(.A(G138), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n481), .B(new_n482), .C1(new_n461), .C2(new_n460), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  XNOR2_X1  g059(.A(KEYINPUT3), .B(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n482), .B1(new_n485), .B2(new_n481), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n464), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  OAI22_X1  g066(.A1(new_n488), .A2(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n487), .A2(new_n492), .ZN(G164));
  INV_X1    g068(.A(G543), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT5), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(KEYINPUT69), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(KEYINPUT5), .A3(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT6), .B(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G88), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G50), .ZN(new_n504));
  OAI22_X1  g079(.A1(new_n501), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  XNOR2_X1  g081(.A(new_n505), .B(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n499), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(G303));
  INV_X1    g086(.A(G303), .ZN(G166));
  OR2_X1    g087(.A1(new_n503), .A2(KEYINPUT71), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n503), .A2(KEYINPUT71), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G51), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT72), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  INV_X1    g094(.A(new_n501), .ZN(new_n520));
  AND2_X1   g095(.A1(G63), .A2(G651), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n520), .A2(G89), .B1(new_n499), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n516), .A2(new_n519), .A3(new_n522), .ZN(G286));
  INV_X1    g098(.A(G286), .ZN(G168));
  AND2_X1   g099(.A1(new_n515), .A2(G52), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n520), .A2(G90), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n499), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n509), .B2(new_n527), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n525), .A2(new_n528), .ZN(G301));
  INV_X1    g104(.A(G301), .ZN(G171));
  AOI22_X1  g105(.A1(new_n499), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G81), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n531), .A2(new_n509), .B1(new_n532), .B2(new_n501), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(G43), .B2(new_n515), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G860), .ZN(G153));
  NAND4_X1  g110(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g111(.A1(G1), .A2(G3), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT8), .ZN(new_n538));
  NAND4_X1  g113(.A1(G319), .A2(G483), .A3(G661), .A4(new_n538), .ZN(G188));
  NAND3_X1  g114(.A1(new_n500), .A2(G53), .A3(G543), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT9), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n541), .A2(KEYINPUT73), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n499), .A2(G91), .A3(new_n500), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n499), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n544), .B2(new_n509), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n541), .B2(KEYINPUT73), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(G299));
  INV_X1    g122(.A(new_n503), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n520), .A2(G87), .B1(new_n548), .B2(G49), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n499), .B2(G74), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(KEYINPUT74), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(KEYINPUT74), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(G288));
  AOI22_X1  g128(.A1(new_n499), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n554), .A2(new_n509), .ZN(new_n555));
  INV_X1    g130(.A(G86), .ZN(new_n556));
  INV_X1    g131(.A(G48), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n501), .A2(new_n556), .B1(new_n503), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(G305));
  AND2_X1   g135(.A1(new_n515), .A2(G47), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n499), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(KEYINPUT75), .B(G85), .ZN(new_n563));
  OAI22_X1  g138(.A1(new_n562), .A2(new_n509), .B1(new_n501), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G290));
  NAND2_X1  g141(.A1(G301), .A2(G868), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n520), .A2(G92), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT10), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n499), .ZN(new_n571));
  INV_X1    g146(.A(G66), .ZN(new_n572));
  INV_X1    g147(.A(G79), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n571), .A2(new_n572), .B1(new_n573), .B2(new_n494), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(KEYINPUT76), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  OAI221_X1 g151(.A(new_n576), .B1(new_n573), .B2(new_n494), .C1(new_n571), .C2(new_n572), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(G651), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n515), .A2(G54), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n570), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n567), .B1(new_n581), .B2(G868), .ZN(G284));
  OAI21_X1  g157(.A(new_n567), .B1(new_n581), .B2(G868), .ZN(G321));
  NAND2_X1  g158(.A1(G286), .A2(G868), .ZN(new_n584));
  INV_X1    g159(.A(G299), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(G868), .ZN(G297));
  OAI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(G868), .ZN(G280));
  INV_X1    g162(.A(G559), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n581), .B1(new_n588), .B2(G860), .ZN(G148));
  NAND2_X1  g164(.A1(new_n581), .A2(new_n588), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G868), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n591), .B1(G868), .B2(new_n534), .ZN(G323));
  XNOR2_X1  g167(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g168(.A1(new_n485), .A2(new_n465), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT12), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT13), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(G2100), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n474), .A2(G123), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n463), .A2(G135), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n600));
  NOR3_X1   g175(.A1(new_n600), .A2(new_n464), .A3(G111), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n464), .B2(G111), .ZN(new_n602));
  OR2_X1    g177(.A1(G99), .A2(G2105), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n602), .A2(G2104), .A3(new_n603), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n598), .B(new_n599), .C1(new_n601), .C2(new_n604), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT78), .B(G2096), .Z(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n597), .A2(new_n607), .ZN(G156));
  XNOR2_X1  g183(.A(KEYINPUT79), .B(KEYINPUT14), .ZN(new_n609));
  XOR2_X1   g184(.A(KEYINPUT15), .B(G2435), .Z(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(G2438), .ZN(new_n611));
  XOR2_X1   g186(.A(G2427), .B(G2430), .Z(new_n612));
  AOI21_X1  g187(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n611), .B2(new_n612), .ZN(new_n614));
  XNOR2_X1  g189(.A(G1341), .B(G1348), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT80), .Z(new_n616));
  XOR2_X1   g191(.A(G2451), .B(G2454), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT16), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n616), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n614), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2443), .B(G2446), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  AND3_X1   g198(.A1(new_n622), .A2(G14), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT81), .Z(G401));
  INV_X1    g200(.A(KEYINPUT18), .ZN(new_n626));
  XOR2_X1   g201(.A(G2084), .B(G2090), .Z(new_n627));
  XNOR2_X1  g202(.A(G2067), .B(G2678), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT17), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n626), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  XOR2_X1   g208(.A(G2072), .B(G2078), .Z(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n629), .B2(KEYINPUT18), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n633), .B(new_n636), .ZN(G227));
  XOR2_X1   g212(.A(G1971), .B(G1976), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT19), .ZN(new_n639));
  XOR2_X1   g214(.A(G1956), .B(G2474), .Z(new_n640));
  XOR2_X1   g215(.A(G1961), .B(G1966), .Z(new_n641));
  AND2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT20), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n640), .A2(new_n641), .ZN(new_n645));
  NOR3_X1   g220(.A1(new_n639), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n639), .B2(new_n645), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1991), .B(G1996), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT82), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1981), .B(G1986), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G229));
  NOR2_X1   g230(.A1(G5), .A2(G16), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT90), .ZN(new_n657));
  INV_X1    g232(.A(G16), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n657), .B1(G301), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT91), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G1961), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(G20), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT94), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT23), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n664), .B1(new_n585), .B2(new_n658), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT95), .B(G1956), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n581), .A2(G16), .ZN(new_n668));
  OR2_X1    g243(.A1(G4), .A2(G16), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n667), .B1(new_n671), .B2(G1348), .ZN(new_n672));
  INV_X1    g247(.A(G1348), .ZN(new_n673));
  AOI22_X1  g248(.A1(new_n670), .A2(new_n673), .B1(new_n666), .B2(new_n665), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n661), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n658), .A2(G19), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(new_n534), .B2(new_n658), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1341), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n658), .A2(G21), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(G168), .B2(new_n658), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G1966), .ZN(new_n681));
  NOR2_X1   g256(.A1(G29), .A2(G35), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(G162), .B2(G29), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G2090), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n685));
  XOR2_X1   g260(.A(new_n684), .B(new_n685), .Z(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G33), .ZN(new_n688));
  AOI22_X1  g263(.A1(new_n485), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n689), .A2(new_n464), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT25), .ZN(new_n691));
  NAND2_X1  g266(.A1(G103), .A2(G2104), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(G2105), .ZN(new_n693));
  NAND4_X1  g268(.A1(new_n464), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n694));
  AOI22_X1  g269(.A1(new_n463), .A2(G139), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT87), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n688), .B1(new_n697), .B2(new_n687), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(G2072), .Z(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g276(.A(G29), .B1(new_n701), .B2(G34), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G34), .B2(new_n701), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G160), .B2(new_n687), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT89), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G2084), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n687), .A2(G32), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n463), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n474), .A2(G129), .ZN(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT26), .Z(new_n711));
  NAND3_X1  g286(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n707), .B1(new_n712), .B2(G29), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT27), .B(G1996), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n687), .A2(G26), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  NAND2_X1  g291(.A1(new_n463), .A2(G140), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n474), .A2(G128), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n464), .A2(G116), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n716), .B1(new_n721), .B2(G29), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT86), .B(G2067), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n713), .A2(new_n714), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n687), .A2(G27), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT92), .Z(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G164), .B2(new_n687), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G2078), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n605), .A2(new_n687), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT30), .B(G28), .ZN(new_n730));
  OR2_X1    g305(.A1(KEYINPUT31), .A2(G11), .ZN(new_n731));
  NAND2_X1  g306(.A1(KEYINPUT31), .A2(G11), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n730), .A2(new_n687), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n724), .A2(new_n728), .A3(new_n729), .A4(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n727), .A2(G2078), .ZN(new_n735));
  OAI22_X1  g310(.A1(new_n713), .A2(new_n714), .B1(new_n722), .B2(new_n723), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n686), .A2(new_n699), .A3(new_n706), .A4(new_n737), .ZN(new_n738));
  NOR4_X1   g313(.A1(new_n675), .A2(new_n678), .A3(new_n681), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT96), .ZN(new_n740));
  NOR2_X1   g315(.A1(G16), .A2(G22), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G166), .B2(G16), .ZN(new_n742));
  INV_X1    g317(.A(G1971), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(G16), .A2(G23), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT84), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G288), .B2(new_n658), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT33), .B(G1976), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n658), .A2(G6), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n559), .B2(new_n658), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT32), .B(G1981), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT83), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n751), .B(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n744), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(KEYINPUT34), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(KEYINPUT34), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n565), .A2(G16), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G16), .B2(G24), .ZN(new_n759));
  INV_X1    g334(.A(G1986), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n463), .A2(G131), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n474), .A2(G119), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n464), .A2(G107), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n763), .B(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G25), .B(new_n767), .S(G29), .Z(new_n768));
  XOR2_X1   g343(.A(KEYINPUT35), .B(G1991), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  AND4_X1   g345(.A1(KEYINPUT85), .A2(new_n761), .A3(new_n762), .A4(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n756), .A2(new_n757), .A3(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT36), .ZN(new_n773));
  OR2_X1    g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n740), .A2(new_n774), .A3(new_n775), .ZN(G150));
  INV_X1    g351(.A(G150), .ZN(G311));
  NOR2_X1   g352(.A1(new_n580), .A2(new_n588), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n499), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n781));
  INV_X1    g356(.A(G93), .ZN(new_n782));
  OAI22_X1  g357(.A1(new_n781), .A2(new_n509), .B1(new_n782), .B2(new_n501), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G55), .B2(new_n515), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n533), .ZN(new_n786));
  INV_X1    g361(.A(new_n515), .ZN(new_n787));
  INV_X1    g362(.A(G43), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n534), .A2(new_n784), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n780), .B(new_n792), .Z(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT39), .ZN(new_n794));
  INV_X1    g369(.A(G860), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(KEYINPUT39), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n784), .A2(new_n795), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT37), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n799), .ZN(G145));
  INV_X1    g375(.A(KEYINPUT100), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n767), .B(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(new_n595), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n804));
  INV_X1    g379(.A(G118), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(G2105), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n474), .A2(G130), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT99), .ZN(new_n808));
  AOI211_X1 g383(.A(new_n806), .B(new_n808), .C1(G142), .C2(new_n463), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n803), .B(new_n809), .Z(new_n810));
  OAI21_X1  g385(.A(KEYINPUT98), .B1(new_n484), .B2(new_n486), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n481), .B1(new_n460), .B2(new_n461), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT4), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n813), .A2(new_n814), .A3(new_n483), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n492), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(new_n721), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(new_n712), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n818), .A2(new_n697), .ZN(new_n819));
  INV_X1    g394(.A(new_n696), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n818), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n810), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n810), .A2(new_n821), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n471), .B(new_n478), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(new_n605), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT102), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n822), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT103), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT101), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n822), .A2(new_n829), .A3(new_n823), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n810), .A2(new_n821), .A3(KEYINPUT101), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n831), .A2(new_n825), .ZN(new_n832));
  AOI21_X1  g407(.A(G37), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g410(.A(new_n585), .B(new_n580), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT41), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n590), .B(new_n792), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n836), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n838), .A2(KEYINPUT104), .A3(new_n839), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n842), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(G303), .B(new_n565), .ZN(new_n847));
  XNOR2_X1  g422(.A(G288), .B(new_n559), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT107), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n849), .A2(new_n850), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT42), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(KEYINPUT105), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT105), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n860), .A3(KEYINPUT42), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n846), .A2(new_n863), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n855), .A2(new_n854), .B1(new_n859), .B2(new_n861), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n842), .A2(new_n844), .A3(new_n845), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(G868), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n784), .A2(G868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(G295));
  NAND2_X1  g446(.A1(new_n846), .A2(new_n863), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n865), .A2(new_n866), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI211_X1 g449(.A(KEYINPUT108), .B(new_n869), .C1(new_n874), .C2(G868), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT108), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(new_n868), .B2(new_n870), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n875), .A2(new_n877), .ZN(G331));
  XNOR2_X1  g453(.A(new_n792), .B(G301), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(G286), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n838), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n879), .A2(G168), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n879), .A2(G168), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n836), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n857), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT109), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT109), .ZN(new_n887));
  NAND4_X1  g462(.A1(new_n881), .A2(new_n884), .A3(new_n887), .A4(new_n857), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n857), .B1(new_n881), .B2(new_n884), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(G37), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n890), .B1(new_n889), .B2(new_n892), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  OAI22_X1  g470(.A1(new_n893), .A2(new_n894), .B1(KEYINPUT110), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n889), .A2(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT43), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n899));
  XOR2_X1   g474(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n896), .A2(new_n901), .ZN(G397));
  OAI21_X1  g477(.A(KEYINPUT111), .B1(new_n816), .B2(G1384), .ZN(new_n903));
  INV_X1    g478(.A(new_n492), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n813), .A2(new_n814), .A3(new_n483), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n814), .B1(new_n813), .B2(new_n483), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT111), .ZN(new_n908));
  INV_X1    g483(.A(G1384), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT50), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n903), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT112), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n909), .B1(new_n487), .B2(new_n492), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n913), .B1(new_n915), .B2(new_n911), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(G40), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n471), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n903), .A2(new_n910), .A3(new_n913), .A4(new_n911), .ZN(new_n920));
  XNOR2_X1  g495(.A(KEYINPUT115), .B(G2084), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n917), .A2(new_n919), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(G1966), .ZN(new_n923));
  AOI21_X1  g498(.A(KEYINPUT45), .B1(new_n903), .B2(new_n910), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n919), .B1(new_n914), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n923), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(G168), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(G8), .ZN(new_n929));
  AOI21_X1  g504(.A(G168), .B1(new_n922), .B2(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(KEYINPUT51), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT62), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT51), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(new_n933), .A3(G8), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G1981), .ZN(new_n936));
  INV_X1    g511(.A(new_n555), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n937), .B2(KEYINPUT113), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT49), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n559), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(KEYINPUT49), .B1(new_n555), .B2(new_n558), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n938), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n903), .A2(new_n910), .A3(new_n919), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(G8), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(KEYINPUT114), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n945), .A2(G8), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT114), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n944), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1976), .ZN(new_n952));
  OR2_X1    g527(.A1(G288), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n945), .A2(G8), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT52), .B1(G288), .B2(new_n952), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n957), .B1(KEYINPUT52), .B2(new_n954), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n951), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(G160), .A2(G40), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n914), .B2(new_n925), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n816), .A2(G1384), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G2078), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT53), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n960), .B1(new_n912), .B2(new_n916), .ZN(new_n968));
  AOI21_X1  g543(.A(G1961), .B1(new_n968), .B2(new_n920), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n971));
  OR4_X1    g546(.A1(new_n971), .A2(new_n924), .A3(G2078), .A4(new_n926), .ZN(new_n972));
  AOI21_X1  g547(.A(G301), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n964), .A2(new_n743), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n816), .A2(KEYINPUT111), .A3(G1384), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n908), .B1(new_n907), .B2(new_n909), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT50), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n919), .B1(new_n914), .B2(KEYINPUT50), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n974), .B1(new_n980), .B2(G2090), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(G8), .ZN(new_n982));
  NAND2_X1  g557(.A1(G303), .A2(G8), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT55), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n974), .B1(new_n986), .B2(G2090), .ZN(new_n987));
  INV_X1    g562(.A(new_n984), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(G8), .A3(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n959), .A2(new_n973), .A3(new_n985), .A4(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT127), .B1(new_n935), .B2(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n959), .A2(new_n985), .A3(new_n989), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT127), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n973), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n931), .A2(new_n934), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT62), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n991), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  AOI211_X1 g573(.A(G1976), .B(G288), .C1(new_n947), .C2(new_n950), .ZN(new_n999));
  NOR2_X1   g574(.A1(G305), .A2(G1981), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n948), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n951), .A2(new_n958), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n1001), .B1(new_n989), .B2(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n959), .A2(KEYINPUT63), .A3(new_n989), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n987), .A2(G8), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n988), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1007), .B1(new_n1006), .B2(new_n1005), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n922), .A2(new_n927), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1009), .A2(G8), .A3(G168), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT116), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1004), .A2(new_n1008), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT63), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1010), .B(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n959), .A2(new_n985), .A3(new_n989), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1003), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n545), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT118), .B(new_n543), .C1(new_n544), .C2(new_n509), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(new_n541), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n542), .A2(new_n546), .A3(KEYINPUT57), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(KEYINPUT119), .A3(new_n1023), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1026), .A2(KEYINPUT122), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT122), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1027), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT119), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1956), .B1(new_n977), .B2(new_n979), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT56), .B(G2072), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n961), .A2(new_n963), .A3(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1029), .B(new_n1033), .C1(new_n1034), .C2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n986), .A2(new_n673), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n945), .A2(KEYINPUT120), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n903), .A2(new_n910), .A3(new_n1040), .A4(new_n919), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1038), .B(KEYINPUT121), .C1(G2067), .C2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT121), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1348), .B1(new_n968), .B2(new_n920), .ZN(new_n1045));
  AOI21_X1  g620(.A(G2067), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1956), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n911), .B1(new_n903), .B2(new_n910), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1049), .B1(new_n1050), .B2(new_n978), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n961), .A2(new_n963), .A3(new_n1035), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n581), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1037), .B1(new_n1048), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT61), .ZN(new_n1057));
  AND3_X1   g632(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1052), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1037), .A2(KEYINPUT61), .A3(new_n1054), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT58), .B(G1341), .Z(new_n1063));
  NAND3_X1  g638(.A1(new_n1039), .A2(new_n1041), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1996), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n961), .A2(new_n1065), .A3(new_n963), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1062), .B1(new_n1067), .B2(new_n534), .ZN(new_n1068));
  AOI211_X1 g643(.A(KEYINPUT59), .B(new_n789), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1060), .B(new_n1061), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT123), .ZN(new_n1071));
  XNOR2_X1  g646(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n580), .B1(new_n1048), .B2(KEYINPUT60), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT60), .ZN(new_n1074));
  AOI211_X1 g649(.A(new_n1074), .B(new_n581), .C1(new_n1043), .C2(new_n1047), .ZN(new_n1075));
  OAI22_X1  g650(.A1(new_n1073), .A2(new_n1075), .B1(KEYINPUT60), .B2(new_n1048), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1056), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n1078));
  INV_X1    g653(.A(new_n970), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n962), .A2(KEYINPUT45), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n464), .B1(new_n469), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1082), .B1(new_n1081), .B2(new_n469), .ZN(new_n1083));
  OR2_X1    g658(.A1(new_n966), .A2(KEYINPUT125), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n966), .A2(KEYINPUT125), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n971), .B(new_n918), .C1(new_n1084), .C2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n466), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1080), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n963), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(KEYINPUT126), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1079), .A2(new_n1090), .A3(G171), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1078), .B1(new_n1091), .B2(new_n973), .ZN(new_n1092));
  OAI21_X1  g667(.A(G171), .B1(new_n1079), .B2(new_n1090), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n970), .A2(G301), .A3(new_n972), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(KEYINPUT54), .A3(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1092), .A2(new_n992), .A3(new_n996), .A4(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n998), .B(new_n1018), .C1(new_n1077), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1080), .A2(new_n919), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n565), .B(new_n760), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n712), .B(new_n1065), .ZN(new_n1101));
  INV_X1    g676(.A(G2067), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n721), .B(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n769), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n767), .A2(new_n1104), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n767), .A2(new_n1104), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1101), .A2(new_n1103), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1099), .B1(new_n1100), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1097), .A2(new_n1108), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1098), .A2(G1986), .A3(G290), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(KEYINPUT48), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1110), .A2(KEYINPUT48), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n1111), .B(new_n1112), .C1(new_n1099), .C2(new_n1107), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1099), .A2(new_n1065), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT46), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1103), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1099), .B1(new_n712), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  XOR2_X1   g693(.A(new_n1118), .B(KEYINPUT47), .Z(new_n1119));
  NAND2_X1  g694(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1120), .A2(new_n1106), .B1(G2067), .B2(new_n721), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1113), .B(new_n1119), .C1(new_n1099), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1109), .A2(new_n1122), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g698(.A1(G229), .A2(new_n458), .A3(new_n624), .A4(G227), .ZN(new_n1125));
  OAI211_X1 g699(.A(new_n834), .B(new_n1125), .C1(new_n893), .C2(new_n894), .ZN(G225));
  INV_X1    g700(.A(G225), .ZN(G308));
endmodule


