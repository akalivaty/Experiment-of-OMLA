//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G137), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  AOI21_X1  g008(.A(KEYINPUT65), .B1(new_n194), .B2(G134), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n198), .B(new_n196), .C1(new_n192), .C2(G137), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(G131), .B1(new_n197), .B2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n198), .B1(new_n192), .B2(G137), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT11), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n203), .A2(new_n204), .A3(new_n199), .A4(new_n193), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(KEYINPUT66), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n207), .B(G131), .C1(new_n197), .C2(new_n200), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT12), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT1), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n213), .A2(new_n215), .A3(new_n216), .A4(G128), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n212), .A2(G143), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n213), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n214), .A2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(G128), .B1(new_n222), .B2(new_n216), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n218), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n227));
  INV_X1    g041(.A(G107), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT79), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G107), .ZN(new_n231));
  AOI21_X1  g045(.A(G104), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(G104), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n227), .B(G101), .C1(new_n232), .C2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n228), .B2(G104), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n233), .ZN(new_n238));
  INV_X1    g052(.A(G101), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n229), .A2(new_n231), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n236), .A2(G104), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n238), .B(new_n239), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n235), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(KEYINPUT79), .B(G107), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n233), .B1(new_n244), .B2(G104), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n227), .B1(new_n245), .B2(G101), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n226), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G104), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n234), .B1(new_n240), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT80), .B1(new_n249), .B2(new_n239), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n213), .A2(new_n215), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n225), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n217), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n250), .A2(new_n253), .A3(new_n242), .A4(new_n235), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n211), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n209), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n247), .A2(KEYINPUT82), .A3(new_n254), .ZN(new_n259));
  AOI211_X1 g073(.A(KEYINPUT83), .B(KEYINPUT12), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT83), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n255), .A2(new_n257), .ZN(new_n262));
  INV_X1    g076(.A(new_n209), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n263), .A3(new_n259), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n261), .B1(new_n264), .B2(new_n210), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n256), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n243), .A2(new_n246), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n213), .A2(new_n220), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n268), .B1(new_n213), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n225), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n217), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n267), .A2(KEYINPUT10), .A3(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n254), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n240), .A2(new_n241), .ZN(new_n276));
  INV_X1    g090(.A(new_n238), .ZN(new_n277));
  OAI21_X1  g091(.A(G101), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT4), .A3(new_n242), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT0), .B(G128), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n221), .B2(new_n223), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT0), .ZN(new_n282));
  INV_X1    g096(.A(G128), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n251), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT4), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n286), .B(G101), .C1(new_n276), .C2(new_n277), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n279), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n273), .A2(new_n275), .A3(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n289), .A2(new_n263), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n266), .A2(new_n291), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G140), .ZN(new_n293));
  INV_X1    g107(.A(G953), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n294), .A2(G227), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n293), .B(new_n295), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n296), .B(KEYINPUT78), .Z(new_n297));
  NOR2_X1   g111(.A1(new_n290), .A2(new_n296), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n289), .A2(new_n263), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n292), .A2(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G469), .B1(new_n300), .B2(G902), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT84), .B(G469), .Z(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n298), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n247), .A2(KEYINPUT82), .A3(new_n254), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT82), .B1(new_n247), .B2(new_n254), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n305), .A2(new_n306), .A3(new_n209), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT83), .B1(new_n307), .B2(KEYINPUT12), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n264), .A2(new_n261), .A3(new_n210), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n304), .B1(new_n310), .B2(new_n256), .ZN(new_n311));
  INV_X1    g125(.A(new_n296), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(new_n291), .B2(new_n299), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n190), .B(new_n303), .C1(new_n311), .C2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n191), .B1(new_n301), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT94), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT93), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n283), .B2(G143), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n214), .A2(KEYINPUT93), .A3(G128), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT13), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n283), .A2(G143), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n321), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n320), .A2(new_n316), .A3(new_n321), .ZN(new_n326));
  OAI21_X1  g140(.A(G134), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT95), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n320), .A2(new_n328), .A3(new_n323), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n328), .B1(new_n320), .B2(new_n323), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n192), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT92), .B(G122), .ZN(new_n333));
  INV_X1    g147(.A(G116), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(G122), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n240), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n244), .B(new_n336), .C1(new_n333), .C2(new_n334), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n327), .A2(new_n332), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n336), .B(KEYINPUT14), .ZN(new_n342));
  OAI21_X1  g156(.A(G107), .B1(new_n342), .B2(new_n335), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n330), .A2(new_n192), .A3(new_n331), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n320), .A2(new_n323), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT95), .ZN(new_n346));
  AOI21_X1  g160(.A(G134), .B1(new_n346), .B2(new_n329), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n339), .B(new_n343), .C1(new_n344), .C2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n189), .A2(G217), .A3(new_n294), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n341), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n350), .B1(new_n341), .B2(new_n348), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n190), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT96), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n341), .A2(new_n348), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n349), .ZN(new_n357));
  AOI21_X1  g171(.A(G902), .B1(new_n357), .B2(new_n351), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT96), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT15), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G478), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT16), .ZN(new_n365));
  INV_X1    g179(.A(G140), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n365), .A2(new_n366), .A3(G125), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(G125), .ZN(new_n368));
  INV_X1    g182(.A(G125), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G140), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(G146), .B(new_n367), .C1(new_n371), .C2(new_n365), .ZN(new_n372));
  INV_X1    g186(.A(G237), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(new_n294), .A3(G214), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(new_n214), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G131), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n374), .B(G143), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n204), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n368), .A2(new_n370), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT91), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n371), .A2(KEYINPUT91), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(KEYINPUT19), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n384), .B1(KEYINPUT19), .B2(new_n371), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n372), .B(new_n379), .C1(new_n385), .C2(G146), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(G146), .A3(new_n383), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n380), .A2(new_n212), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT18), .A2(G131), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n377), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n375), .A2(KEYINPUT18), .A3(G131), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(G113), .B(G122), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(new_n248), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n375), .A2(KEYINPUT17), .A3(G131), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n379), .B2(KEYINPUT17), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT73), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n372), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n367), .B1(new_n371), .B2(new_n365), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n212), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n402), .B(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n396), .B(new_n393), .C1(new_n400), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n398), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(G475), .A2(G902), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n407), .A2(new_n413), .A3(new_n408), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n393), .B1(new_n400), .B2(new_n405), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n397), .ZN(new_n416));
  AOI21_X1  g230(.A(G902), .B1(new_n416), .B2(new_n406), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n412), .A2(new_n414), .B1(new_n418), .B2(G475), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n363), .B1(new_n358), .B2(new_n359), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G234), .ZN(new_n422));
  OAI211_X1 g236(.A(G952), .B(new_n294), .C1(new_n422), .C2(new_n373), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(KEYINPUT97), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(G898), .ZN(new_n426));
  AOI211_X1 g240(.A(new_n190), .B(new_n294), .C1(G234), .C2(G237), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n364), .A2(new_n419), .A3(new_n421), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT98), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n420), .B1(new_n361), .B2(new_n363), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT98), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n432), .A2(new_n433), .A3(new_n429), .A4(new_n419), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G214), .B1(G237), .B2(G902), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G122), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT85), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n334), .A2(G119), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT67), .ZN(new_n442));
  INV_X1    g256(.A(G119), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(G116), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n334), .A2(KEYINPUT67), .A3(G119), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n441), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT2), .B(G113), .Z(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(KEYINPUT68), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT68), .B1(new_n446), .B2(new_n447), .ZN(new_n450));
  OAI22_X1  g264(.A1(new_n449), .A2(new_n450), .B1(new_n446), .B2(new_n447), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n287), .A3(new_n279), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n443), .A2(G116), .ZN(new_n453));
  OAI21_X1  g267(.A(G113), .B1(new_n453), .B2(KEYINPUT5), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n446), .B2(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n446), .A2(new_n447), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT68), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n455), .B1(new_n458), .B2(new_n448), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n267), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n440), .B1(new_n452), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n462));
  AOI21_X1  g276(.A(KEYINPUT86), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n452), .A2(new_n460), .A3(new_n440), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT6), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n463), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n461), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n467), .A2(KEYINPUT86), .A3(KEYINPUT6), .A4(new_n464), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n285), .A2(G125), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n470), .B1(G125), .B2(new_n226), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n294), .A2(G224), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(G210), .B1(G237), .B2(G902), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n250), .A2(KEYINPUT87), .A3(new_n242), .A4(new_n235), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n476), .A2(new_n459), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n459), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n439), .B(KEYINPUT8), .Z(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(KEYINPUT88), .A2(KEYINPUT7), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n226), .A2(G125), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n281), .A2(new_n284), .A3(new_n369), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n472), .A2(KEYINPUT7), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n471), .A2(KEYINPUT7), .A3(new_n472), .A4(new_n481), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n480), .A2(new_n464), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(KEYINPUT89), .A3(new_n190), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n190), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT89), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n474), .A2(new_n475), .A3(new_n489), .A4(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n475), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n489), .ZN(new_n495));
  INV_X1    g309(.A(new_n473), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n496), .B1(new_n466), .B2(new_n468), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n494), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n437), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n315), .A2(new_n435), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n206), .A2(new_n285), .A3(new_n208), .ZN(new_n501));
  INV_X1    g315(.A(new_n193), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n192), .A2(G137), .ZN(new_n503));
  OAI21_X1  g317(.A(G131), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n205), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n272), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n508), .B1(new_n505), .B2(new_n272), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n510), .A2(new_n501), .A3(KEYINPUT69), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT69), .B1(new_n510), .B2(new_n501), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n451), .B(new_n509), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n446), .A2(new_n447), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n458), .B2(new_n448), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n501), .A2(new_n506), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n373), .A2(new_n294), .A3(G210), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT26), .B(G101), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n501), .A2(new_n506), .A3(new_n515), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n515), .B1(new_n501), .B2(new_n506), .ZN(new_n525));
  OAI21_X1  g339(.A(KEYINPUT28), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT28), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n516), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n520), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n523), .A2(KEYINPUT31), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT70), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n510), .A2(new_n501), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT69), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n510), .A2(new_n501), .A3(KEYINPUT69), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n515), .B1(new_n507), .B2(new_n508), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n521), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT31), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n532), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND4_X1   g355(.A1(new_n532), .A2(new_n513), .A3(new_n540), .A4(new_n522), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n531), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT71), .ZN(new_n544));
  NOR2_X1   g358(.A1(G472), .A2(G902), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n545), .B(KEYINPUT72), .Z(new_n546));
  INV_X1    g360(.A(KEYINPUT71), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n531), .B(new_n547), .C1(new_n541), .C2(new_n542), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT32), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g365(.A1(new_n544), .A2(new_n548), .A3(KEYINPUT32), .A4(new_n546), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n513), .A2(new_n516), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n530), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT29), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n526), .A2(new_n520), .A3(new_n528), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n190), .B1(new_n556), .B2(new_n555), .ZN(new_n558));
  OAI21_X1  g372(.A(G472), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n551), .A2(new_n552), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT23), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n443), .B2(G128), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n283), .A2(KEYINPUT23), .A3(G119), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n562), .B(new_n563), .C1(G119), .C2(new_n283), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n564), .A2(G110), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT74), .ZN(new_n566));
  XNOR2_X1  g380(.A(G119), .B(G128), .ZN(new_n567));
  XOR2_X1   g381(.A(KEYINPUT24), .B(G110), .Z(new_n568));
  OAI22_X1  g382(.A1(new_n565), .A2(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n565), .A2(new_n566), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n372), .B(new_n388), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n564), .A2(G110), .B1(new_n567), .B2(new_n568), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n405), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT22), .B(G137), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n187), .A2(new_n422), .A3(G953), .ZN(new_n576));
  XOR2_X1   g390(.A(new_n575), .B(new_n576), .Z(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n571), .A2(new_n573), .A3(new_n577), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT25), .ZN(new_n581));
  AOI21_X1  g395(.A(G902), .B1(new_n581), .B2(KEYINPUT75), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n581), .A2(KEYINPUT75), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G217), .B1(new_n422), .B2(G902), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n583), .B2(new_n584), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n579), .A2(new_n580), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n190), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT76), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT77), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n560), .A2(new_n594), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n500), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(G101), .ZN(G3));
  INV_X1    g411(.A(G478), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n349), .B2(KEYINPUT99), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n352), .A2(new_n353), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n601), .B1(new_n352), .B2(new_n353), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n598), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n598), .A2(new_n190), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n606), .B1(new_n358), .B2(new_n598), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n419), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n499), .A2(new_n429), .A3(new_n609), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n544), .A2(new_n548), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n544), .A2(new_n190), .A3(new_n548), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n611), .A2(new_n546), .B1(new_n612), .B2(G472), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n610), .A2(new_n315), .A3(new_n613), .A4(new_n594), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT34), .B(G104), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NAND2_X1  g430(.A1(new_n493), .A2(new_n498), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n436), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n409), .A2(new_n411), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n410), .B1(new_n407), .B2(new_n408), .ZN(new_n620));
  INV_X1    g434(.A(G475), .ZN(new_n621));
  OAI22_X1  g435(.A1(new_n619), .A2(new_n620), .B1(new_n621), .B2(new_n417), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n432), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n618), .A2(new_n428), .A3(new_n623), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n624), .A2(new_n594), .A3(new_n315), .A4(new_n613), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT35), .B(G107), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NOR2_X1   g441(.A1(new_n578), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n574), .B(new_n628), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n585), .A2(new_n587), .B1(new_n591), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n431), .B2(new_n434), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n315), .A2(new_n613), .A3(new_n631), .A4(new_n499), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT37), .B(G110), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT100), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n632), .B(new_n634), .ZN(G12));
  INV_X1    g449(.A(new_n630), .ZN(new_n636));
  INV_X1    g450(.A(G900), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n425), .B1(new_n637), .B2(new_n427), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n432), .A2(new_n622), .A3(new_n638), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n499), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n560), .A2(new_n640), .A3(new_n315), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G128), .ZN(G30));
  XOR2_X1   g456(.A(KEYINPUT101), .B(KEYINPUT39), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n638), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n315), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n645), .B(KEYINPUT40), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n617), .B(KEYINPUT38), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n432), .A2(new_n419), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n647), .A2(new_n436), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n553), .A2(new_n520), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n524), .A2(new_n525), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n190), .B1(new_n653), .B2(new_n520), .ZN(new_n654));
  OAI21_X1  g468(.A(G472), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n551), .A2(new_n552), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n649), .A2(new_n636), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n646), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G143), .ZN(G45));
  INV_X1    g474(.A(new_n414), .ZN(new_n661));
  OAI22_X1  g475(.A1(new_n661), .A2(new_n620), .B1(new_n621), .B2(new_n417), .ZN(new_n662));
  INV_X1    g476(.A(new_n604), .ZN(new_n663));
  OAI21_X1  g477(.A(G478), .B1(new_n663), .B2(new_n602), .ZN(new_n664));
  INV_X1    g478(.A(new_n638), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n662), .A2(new_n664), .A3(new_n607), .A4(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n630), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n667), .A2(new_n499), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n560), .A2(new_n315), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n560), .A2(new_n315), .A3(new_n668), .A4(KEYINPUT102), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n313), .B1(new_n266), .B2(new_n298), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n675), .B1(new_n676), .B2(G902), .ZN(new_n677));
  OAI211_X1 g491(.A(KEYINPUT103), .B(new_n190), .C1(new_n311), .C2(new_n313), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n677), .A2(new_n678), .A3(G469), .ZN(new_n679));
  INV_X1    g493(.A(new_n191), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n680), .A3(new_n314), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT104), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n679), .A2(new_n683), .A3(new_n680), .A4(new_n314), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n560), .A2(new_n610), .A3(new_n594), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT41), .B(G113), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  AND3_X1   g503(.A1(new_n624), .A2(new_n594), .A3(new_n560), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n690), .A2(new_n691), .A3(new_n682), .A4(new_n684), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n624), .A2(new_n560), .A3(new_n594), .ZN(new_n693));
  OAI21_X1  g507(.A(KEYINPUT105), .B1(new_n685), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  AND3_X1   g510(.A1(new_n679), .A2(new_n680), .A3(new_n314), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(new_n560), .A3(new_n499), .A4(new_n631), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT106), .B(G119), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G21));
  AND2_X1   g514(.A1(new_n543), .A2(new_n546), .ZN(new_n701));
  AOI211_X1 g515(.A(new_n593), .B(new_n701), .C1(new_n612), .C2(G472), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n499), .A2(new_n429), .A3(new_n648), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n682), .A2(new_n684), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  AOI21_X1  g519(.A(new_n701), .B1(new_n612), .B2(G472), .ZN(new_n706));
  INV_X1    g520(.A(new_n666), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n706), .A2(new_n636), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n679), .A2(new_n680), .A3(new_n499), .A4(new_n314), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n369), .ZN(G27));
  NAND3_X1  g525(.A1(new_n549), .A2(KEYINPUT109), .A3(new_n550), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n712), .A2(new_n552), .A3(new_n559), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT109), .B1(new_n549), .B2(new_n550), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n593), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  AND4_X1   g530(.A1(new_n680), .A2(new_n493), .A3(new_n498), .A4(new_n436), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n308), .A2(new_n309), .B1(new_n255), .B2(new_n211), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n297), .B1(new_n718), .B2(new_n290), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n298), .A2(new_n299), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n719), .A2(KEYINPUT107), .A3(G469), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(G469), .A2(G902), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n314), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT107), .B1(new_n300), .B2(G469), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n717), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n717), .B(KEYINPUT108), .C1(new_n723), .C2(new_n724), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n716), .A2(new_n707), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n595), .B1(new_n727), .B2(new_n728), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n730), .A2(KEYINPUT42), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  INV_X1    g548(.A(new_n595), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n729), .A2(new_n735), .A3(new_n639), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT110), .B(G134), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G36));
  NOR2_X1   g552(.A1(new_n617), .A2(new_n437), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n605), .A2(new_n608), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n419), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n636), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n613), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n739), .B1(new_n745), .B2(KEYINPUT44), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(KEYINPUT44), .B2(new_n745), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n300), .A2(KEYINPUT45), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n300), .A2(KEYINPUT45), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(G469), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT46), .B1(new_n750), .B2(new_n722), .ZN(new_n751));
  INV_X1    g565(.A(new_n314), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n750), .A2(KEYINPUT46), .A3(new_n722), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n191), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n755), .A2(KEYINPUT111), .A3(new_n644), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT111), .B1(new_n755), .B2(new_n644), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n747), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G137), .ZN(G39));
  INV_X1    g573(.A(new_n739), .ZN(new_n760));
  NOR4_X1   g574(.A1(new_n560), .A2(new_n760), .A3(new_n594), .A4(new_n666), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(KEYINPUT112), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n755), .A2(KEYINPUT47), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n755), .A2(KEYINPUT47), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G140), .ZN(G42));
  NAND2_X1  g581(.A1(new_n679), .A2(new_n314), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT49), .Z(new_n769));
  INV_X1    g583(.A(new_n647), .ZN(new_n770));
  NOR4_X1   g584(.A1(new_n741), .A2(new_n593), .A3(new_n191), .A4(new_n437), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n769), .A2(new_n657), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n704), .B(new_n698), .C1(new_n685), .C2(new_n686), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n774), .B1(new_n692), .B2(new_n694), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n432), .A2(new_n662), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n499), .A2(new_n429), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n315), .A3(new_n613), .A4(new_n594), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n632), .A3(KEYINPUT113), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT113), .B1(new_n778), .B2(new_n632), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n614), .B1(new_n595), .B2(new_n500), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  AOI211_X1 g597(.A(new_n630), .B(new_n701), .C1(new_n612), .C2(G472), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n729), .A2(new_n707), .A3(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n636), .A2(new_n432), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n786), .A2(new_n622), .A3(new_n638), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n560), .A2(new_n315), .A3(new_n739), .A4(new_n787), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n736), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n775), .A2(new_n783), .A3(new_n789), .A4(new_n733), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n697), .A2(new_n784), .A3(new_n499), .A4(new_n707), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n638), .A2(new_n191), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n499), .A2(new_n648), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n719), .A2(G469), .A3(new_n720), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT107), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n314), .A3(new_n721), .A4(new_n722), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n656), .A2(new_n793), .A3(new_n630), .A4(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n791), .A2(new_n641), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(new_n799), .B2(new_n673), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n801));
  INV_X1    g615(.A(new_n641), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n801), .B1(new_n802), .B2(new_n710), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n791), .A2(KEYINPUT114), .A3(new_n641), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n803), .A2(new_n673), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n798), .A2(KEYINPUT52), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n800), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n773), .B1(new_n790), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT115), .ZN(new_n809));
  INV_X1    g623(.A(new_n790), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n799), .A2(KEYINPUT52), .A3(new_n673), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT116), .B1(new_n811), .B2(new_n800), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n671), .A2(new_n672), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n791), .A2(new_n798), .A3(new_n641), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n799), .A2(KEYINPUT52), .A3(new_n673), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n810), .A2(KEYINPUT53), .A3(new_n812), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n821), .B(new_n773), .C1(new_n790), .C2(new_n807), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n809), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT54), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n698), .B1(new_n685), .B2(new_n686), .ZN(new_n825));
  INV_X1    g639(.A(new_n704), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n728), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT108), .B1(new_n797), .B2(new_n717), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n707), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n712), .A2(new_n552), .A3(new_n559), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n592), .B(new_n588), .C1(new_n831), .C2(new_n714), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT42), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n731), .A2(new_n732), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n695), .A2(new_n827), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n778), .A2(new_n632), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(new_n596), .A3(new_n614), .A4(new_n779), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n736), .A2(new_n785), .A3(new_n788), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n812), .A2(new_n835), .A3(new_n819), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n775), .A2(KEYINPUT53), .A3(new_n733), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n807), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT117), .B1(new_n783), .B2(new_n789), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n839), .A2(new_n840), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n773), .A2(new_n842), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n765), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n679), .A2(new_n191), .A3(new_n314), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n763), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n702), .A2(new_n425), .A3(new_n743), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n739), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n854), .A2(KEYINPUT119), .A3(new_n857), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n855), .A2(new_n437), .A3(new_n770), .A4(new_n697), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT50), .Z(new_n863));
  NAND2_X1  g677(.A1(new_n697), .A2(new_n739), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT120), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n657), .A2(new_n594), .A3(new_n425), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n740), .A2(new_n662), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n743), .A2(new_n425), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n784), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n863), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n860), .A2(new_n861), .A3(new_n873), .ZN(new_n874));
  XOR2_X1   g688(.A(KEYINPUT118), .B(KEYINPUT51), .Z(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n873), .A2(new_n858), .A3(KEYINPUT51), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n871), .A2(KEYINPUT48), .A3(new_n716), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n866), .A2(new_n609), .A3(new_n867), .ZN(new_n879));
  INV_X1    g693(.A(G952), .ZN(new_n880));
  INV_X1    g694(.A(new_n709), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n880), .B(G953), .C1(new_n855), .C2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT48), .B1(new_n871), .B2(new_n716), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n877), .A2(new_n878), .A3(new_n885), .ZN(new_n886));
  AND4_X1   g700(.A1(new_n824), .A2(new_n851), .A3(new_n876), .A4(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(G952), .A2(G953), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n772), .B1(new_n887), .B2(new_n888), .ZN(G75));
  XNOR2_X1  g703(.A(new_n469), .B(new_n473), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT55), .ZN(new_n891));
  INV_X1    g705(.A(G210), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n849), .A2(new_n892), .A3(new_n190), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n891), .B1(new_n893), .B2(KEYINPUT56), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT56), .ZN(new_n895));
  INV_X1    g709(.A(new_n891), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n842), .A2(new_n773), .ZN(new_n897));
  INV_X1    g711(.A(new_n843), .ZN(new_n898));
  INV_X1    g712(.A(new_n847), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n805), .A2(new_n806), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(new_n816), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n846), .B1(new_n839), .B2(new_n840), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n898), .A2(new_n899), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(G902), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n895), .B(new_n896), .C1(new_n905), .C2(new_n892), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n294), .A2(G952), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n894), .A2(new_n906), .A3(new_n908), .ZN(G51));
  XOR2_X1   g723(.A(new_n722), .B(KEYINPUT57), .Z(new_n910));
  AND3_X1   g724(.A1(new_n897), .A2(new_n850), .A3(new_n903), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n850), .B1(new_n897), .B2(new_n903), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n676), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OR2_X1    g729(.A1(new_n905), .A2(new_n750), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n907), .B1(new_n915), .B2(new_n916), .ZN(G54));
  INV_X1    g731(.A(new_n905), .ZN(new_n918));
  NAND2_X1  g732(.A1(KEYINPUT58), .A2(G475), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT121), .Z(new_n920));
  AOI21_X1  g734(.A(new_n407), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  AND4_X1   g735(.A1(G902), .A2(new_n904), .A3(new_n407), .A4(new_n920), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n921), .A2(new_n922), .A3(new_n907), .ZN(G60));
  NAND2_X1  g737(.A1(new_n603), .A2(new_n604), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n606), .B(KEYINPUT59), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n911), .B2(new_n912), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n908), .ZN(new_n928));
  INV_X1    g742(.A(new_n925), .ZN(new_n929));
  INV_X1    g743(.A(new_n842), .ZN(new_n930));
  AOI22_X1  g744(.A1(new_n930), .A2(KEYINPUT53), .B1(new_n808), .B2(KEYINPUT115), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n850), .B1(new_n931), .B2(new_n822), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n929), .B1(new_n932), .B2(new_n911), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n928), .B1(new_n924), .B2(new_n933), .ZN(G63));
  NAND2_X1  g748(.A1(G217), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT60), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n904), .A2(new_n629), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n936), .B1(new_n897), .B2(new_n903), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n938), .B(new_n908), .C1(new_n589), .C2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT122), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT61), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n939), .A2(new_n589), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n907), .B1(new_n939), .B2(new_n629), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT122), .B1(new_n939), .B2(new_n629), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n944), .B(new_n945), .C1(new_n946), .C2(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n943), .A2(new_n947), .ZN(G66));
  INV_X1    g762(.A(G224), .ZN(new_n949));
  OAI21_X1  g763(.A(G953), .B1(new_n426), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n775), .A2(new_n783), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n951), .B2(G953), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n466), .B(new_n468), .C1(G898), .C2(new_n294), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G69));
  NAND2_X1  g768(.A1(new_n537), .A2(new_n509), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(new_n385), .ZN(new_n956));
  OAI211_X1 g770(.A(G900), .B(G953), .C1(new_n956), .C2(G227), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(G227), .B2(new_n956), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n499), .A2(new_n648), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n716), .B(new_n959), .C1(new_n756), .C2(new_n757), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(new_n758), .A3(new_n766), .A4(new_n805), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n733), .A2(new_n736), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT124), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(G953), .B1(new_n964), .B2(new_n956), .ZN(new_n965));
  INV_X1    g779(.A(new_n956), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n967), .B1(new_n805), .B2(new_n659), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT123), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n805), .A2(new_n967), .A3(new_n659), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n739), .B1(new_n609), .B2(new_n776), .ZN(new_n972));
  OR3_X1    g786(.A1(new_n595), .A2(new_n645), .A3(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n758), .A2(new_n766), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n966), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n958), .B1(new_n965), .B2(new_n975), .ZN(G72));
  NOR3_X1   g790(.A1(new_n970), .A2(new_n974), .A3(new_n650), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n513), .A2(new_n516), .A3(new_n530), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n961), .A2(new_n963), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n951), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n650), .A2(new_n978), .ZN(new_n981));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT63), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT125), .Z(new_n984));
  AOI21_X1  g798(.A(new_n907), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  OR2_X1    g800(.A1(new_n554), .A2(KEYINPUT126), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n539), .B1(new_n554), .B2(KEYINPUT126), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n983), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n823), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n823), .A2(KEYINPUT127), .A3(new_n989), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n986), .B1(new_n992), .B2(new_n993), .ZN(G57));
endmodule


