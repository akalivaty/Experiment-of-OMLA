//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:34:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355, new_n1356;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G116), .ZN(new_n211));
  INV_X1    g0011(.A(G270), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n213), .B(new_n219), .C1(G107), .C2(G264), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT66), .B(G68), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G238), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n208), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT67), .Z(new_n226));
  INV_X1    g0026(.A(G13), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n208), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G20), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n215), .B1(new_n203), .B2(KEYINPUT65), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n235), .B1(KEYINPUT65), .B2(new_n203), .ZN(new_n236));
  OAI221_X1 g0036(.A(new_n231), .B1(new_n234), .B2(new_n236), .C1(new_n223), .C2(new_n224), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n226), .A2(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT69), .ZN(new_n245));
  XOR2_X1   g0045(.A(G264), .B(G270), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n243), .B(new_n247), .Z(G358));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G223), .A3(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G222), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n257), .B1(new_n258), .B2(new_n256), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G41), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n233), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT70), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(KEYINPUT70), .A2(G33), .A3(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(new_n233), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(G274), .A3(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n273), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G226), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n266), .A2(new_n274), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G200), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n266), .A2(G190), .A3(new_n274), .A4(new_n277), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n232), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n217), .A2(KEYINPUT8), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n283), .B(KEYINPUT71), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT8), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G58), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT72), .ZN(new_n287));
  XNOR2_X1  g0087(.A(new_n286), .B(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n207), .A2(G33), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n292));
  INV_X1    g0092(.A(G150), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n282), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(G50), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n282), .B1(new_n206), .B2(G20), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n299), .B1(new_n300), .B2(G50), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(KEYINPUT9), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n297), .B2(new_n301), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n279), .B(new_n280), .C1(new_n303), .C2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n279), .A2(new_n280), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(KEYINPUT75), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n306), .B(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT73), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n286), .A2(new_n283), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n294), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT15), .B(G87), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n313), .B1(new_n207), .B2(new_n258), .C1(new_n290), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n282), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n300), .A2(G77), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(new_n317), .C1(G77), .C2(new_n298), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n256), .A2(G238), .A3(G1698), .ZN(new_n319));
  INV_X1    g0119(.A(G107), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n319), .B1(new_n320), .B2(new_n256), .C1(new_n260), .C2(new_n218), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n265), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n270), .A2(G274), .ZN(new_n323));
  AOI22_X1  g0123(.A1(G244), .A2(new_n276), .B1(new_n323), .B2(new_n273), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n311), .B(new_n318), .C1(new_n325), .C2(G169), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(G169), .B1(new_n322), .B2(new_n324), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n317), .B1(G77), .B2(new_n298), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n282), .B2(new_n315), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT73), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n326), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n325), .A2(G190), .ZN(new_n334));
  INV_X1    g0134(.A(G200), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n334), .B(new_n331), .C1(new_n335), .C2(new_n325), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT74), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n278), .A2(G179), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n278), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n302), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n310), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n289), .A2(new_n300), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n345), .B1(new_n298), .B2(new_n289), .ZN(new_n346));
  INV_X1    g0146(.A(G33), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT3), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT3), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n349), .A2(KEYINPUT79), .A3(G33), .ZN(new_n350));
  AOI21_X1  g0150(.A(KEYINPUT79), .B1(new_n349), .B2(G33), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n353), .A3(new_n207), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n349), .A2(G33), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT79), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n347), .B2(KEYINPUT3), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n349), .A2(KEYINPUT79), .A3(G33), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT7), .B1(new_n359), .B2(G20), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(new_n360), .A3(G68), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT80), .ZN(new_n362));
  INV_X1    g0162(.A(G159), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n295), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n202), .B1(new_n221), .B2(G58), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n362), .B(new_n365), .C1(new_n366), .C2(new_n207), .ZN(new_n367));
  AND2_X1   g0167(.A1(KEYINPUT66), .A2(G68), .ZN(new_n368));
  NOR2_X1   g0168(.A1(KEYINPUT66), .A2(G68), .ZN(new_n369));
  OAI21_X1  g0169(.A(G58), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n207), .B1(new_n370), .B2(new_n203), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT80), .B1(new_n371), .B2(new_n364), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n361), .A2(KEYINPUT16), .A3(new_n367), .A4(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n373), .A2(new_n282), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n372), .A2(new_n367), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT81), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n349), .B2(G33), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n347), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n349), .A2(G33), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n353), .B1(new_n381), .B2(new_n207), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n368), .A2(new_n369), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n256), .A2(KEYINPUT7), .A3(G20), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n375), .B1(new_n376), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n346), .B1(new_n374), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n270), .A2(new_n275), .A3(G232), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n274), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n347), .A2(new_n209), .ZN(new_n390));
  NOR2_X1   g0190(.A1(G223), .A2(G1698), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n216), .B2(G1698), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n359), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n265), .B1(new_n393), .B2(KEYINPUT82), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT82), .ZN(new_n395));
  AOI211_X1 g0195(.A(new_n395), .B(new_n390), .C1(new_n359), .C2(new_n392), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n389), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G169), .ZN(new_n398));
  OAI211_X1 g0198(.A(G179), .B(new_n389), .C1(new_n394), .C2(new_n396), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT18), .B1(new_n387), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n397), .A2(new_n335), .ZN(new_n403));
  INV_X1    g0203(.A(G190), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n404), .B(new_n389), .C1(new_n394), .C2(new_n396), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n386), .A2(new_n282), .A3(new_n373), .ZN(new_n407));
  INV_X1    g0207(.A(new_n346), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n387), .A2(KEYINPUT17), .A3(new_n406), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n407), .A2(new_n408), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT18), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n400), .A3(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n402), .A2(new_n411), .A3(new_n412), .A4(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n348), .A2(new_n380), .A3(G232), .A4(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT76), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT76), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n256), .A2(new_n419), .A3(G232), .A4(G1698), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n348), .A2(new_n380), .A3(G226), .A4(new_n259), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G97), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n264), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n270), .A2(new_n275), .A3(G238), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n274), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT13), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n274), .A2(new_n427), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT13), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n424), .B1(new_n420), .B2(new_n418), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n430), .B(new_n431), .C1(new_n432), .C2(new_n264), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G200), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT12), .ZN(new_n436));
  INV_X1    g0236(.A(new_n298), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n436), .B1(new_n383), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT77), .ZN(new_n439));
  INV_X1    g0239(.A(G68), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n439), .A2(new_n441), .B1(G68), .B2(new_n300), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n221), .A2(new_n207), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n295), .A2(new_n215), .B1(new_n290), .B2(new_n258), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n282), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT11), .ZN(new_n446));
  AND2_X1   g0246(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n429), .A2(G190), .A3(new_n433), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n435), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n434), .A2(G169), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT14), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n429), .A2(G179), .A3(new_n433), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT14), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n434), .A2(new_n453), .A3(G169), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT78), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n442), .A2(new_n456), .A3(new_n446), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n456), .B1(new_n442), .B2(new_n446), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n449), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n337), .A2(new_n338), .ZN(new_n462));
  NOR4_X1   g0262(.A1(new_n344), .A2(new_n416), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n272), .A2(G1), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(G41), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT84), .B1(new_n465), .B2(G41), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT84), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(new_n271), .A3(KEYINPUT5), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n467), .A2(new_n270), .A3(new_n471), .A4(G274), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n271), .A2(KEYINPUT5), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n464), .A2(new_n473), .A3(new_n466), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n270), .A2(new_n474), .A3(G270), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G257), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n477), .A2(G1698), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n359), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT88), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT88), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n359), .A2(new_n481), .A3(new_n478), .ZN(new_n482));
  AND2_X1   g0282(.A1(G264), .A2(G1698), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n348), .A2(new_n380), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n359), .A2(new_n483), .B1(G303), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n480), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n476), .B1(new_n486), .B2(new_n265), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n281), .A2(new_n232), .B1(G20), .B2(new_n211), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G33), .A2(G283), .ZN(new_n489));
  INV_X1    g0289(.A(G97), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n489), .B(new_n207), .C1(G33), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n492), .B(KEYINPUT20), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n437), .A2(new_n211), .ZN(new_n494));
  INV_X1    g0294(.A(new_n282), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n495), .B(new_n298), .C1(G1), .C2(new_n347), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n494), .B1(new_n496), .B2(new_n211), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n487), .B(G179), .C1(new_n493), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT21), .ZN(new_n499));
  OAI21_X1  g0299(.A(G169), .B1(new_n493), .B2(new_n497), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n487), .B2(new_n500), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n487), .A2(new_n500), .A3(new_n499), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n498), .B(new_n501), .C1(new_n502), .C2(KEYINPUT89), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT89), .ZN(new_n505));
  NOR4_X1   g0305(.A1(new_n487), .A2(new_n500), .A3(new_n505), .A4(new_n499), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n487), .A2(G190), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n493), .A2(new_n497), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n487), .B2(new_n335), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT24), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n359), .A2(new_n207), .A3(G87), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT22), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n484), .A2(G20), .A3(new_n209), .ZN(new_n517));
  XOR2_X1   g0317(.A(KEYINPUT90), .B(KEYINPUT22), .Z(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT23), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n207), .B2(G107), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n320), .A2(KEYINPUT23), .A3(G20), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n347), .A2(new_n211), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n207), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n514), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n515), .A2(KEYINPUT22), .B1(new_n517), .B2(new_n518), .ZN(new_n527));
  INV_X1    g0327(.A(new_n525), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n527), .A2(KEYINPUT24), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n282), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n437), .A2(KEYINPUT25), .A3(new_n320), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT25), .B1(new_n437), .B2(new_n320), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n496), .A2(new_n320), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n270), .A2(new_n474), .A3(G264), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G250), .A2(G1698), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n477), .B2(G1698), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n359), .A2(new_n538), .B1(G33), .B2(G294), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n472), .B(new_n536), .C1(new_n539), .C2(new_n264), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n335), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(G190), .B2(new_n540), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n530), .A2(new_n535), .A3(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n270), .A2(new_n474), .A3(G264), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G294), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n477), .A2(G1698), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(G250), .B2(G1698), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n545), .B1(new_n352), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n544), .B1(new_n548), .B2(new_n265), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(new_n327), .A3(new_n472), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n540), .A2(new_n341), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n520), .A2(new_n514), .A3(new_n525), .ZN(new_n553));
  OAI21_X1  g0353(.A(KEYINPUT24), .B1(new_n527), .B2(new_n528), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n495), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n552), .B1(new_n555), .B2(new_n534), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n543), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n270), .A2(new_n474), .A3(G257), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n472), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G244), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n561), .A2(G1698), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT4), .B1(new_n359), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n348), .A2(new_n380), .A3(G250), .A4(G1698), .ZN(new_n564));
  AND2_X1   g0364(.A1(KEYINPUT4), .A2(G244), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n348), .A2(new_n380), .A3(new_n565), .A4(new_n259), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n566), .A3(new_n489), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n265), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n560), .A2(new_n568), .A3(new_n404), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n359), .A2(new_n562), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT4), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n567), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n559), .B1(new_n574), .B2(new_n265), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n569), .B1(new_n575), .B2(G200), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n437), .A2(new_n490), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n496), .B2(new_n490), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n384), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n381), .A2(new_n207), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(G107), .C1(new_n581), .C2(new_n353), .ZN(new_n582));
  XNOR2_X1  g0382(.A(G97), .B(G107), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT6), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n584), .A2(new_n490), .A3(G107), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n589));
  AOI211_X1 g0389(.A(KEYINPUT83), .B(new_n495), .C1(new_n582), .C2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT83), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n582), .A2(new_n589), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(new_n282), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n576), .B(new_n579), .C1(new_n590), .C2(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n382), .A2(new_n320), .A3(new_n384), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n586), .B1(new_n584), .B2(new_n583), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n596), .A2(new_n207), .B1(new_n258), .B2(new_n295), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT83), .B1(new_n598), .B2(new_n495), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n592), .A2(new_n591), .A3(new_n282), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n578), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n575), .A2(new_n327), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n560), .A2(new_n568), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n341), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n594), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n314), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n298), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n496), .A2(new_n209), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n359), .A2(new_n207), .A3(G68), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT19), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n290), .B2(new_n490), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT86), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n207), .B1(new_n423), .B2(new_n611), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n209), .A2(new_n490), .A3(new_n320), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AND3_X1   g0416(.A1(new_n614), .A2(new_n613), .A3(new_n615), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n610), .B(new_n612), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT87), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n495), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n616), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n614), .A2(new_n613), .A3(new_n615), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n623), .A2(KEYINPUT87), .A3(new_n610), .A4(new_n612), .ZN(new_n624));
  AOI211_X1 g0424(.A(new_n608), .B(new_n609), .C1(new_n620), .C2(new_n624), .ZN(new_n625));
  OR3_X1    g0425(.A1(new_n272), .A2(G1), .A3(G274), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n270), .B(new_n626), .C1(G250), .C2(new_n464), .ZN(new_n627));
  NOR2_X1   g0427(.A1(G238), .A2(G1698), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n561), .B2(G1698), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n524), .B1(new_n359), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT85), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n265), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI211_X1 g0432(.A(KEYINPUT85), .B(new_n524), .C1(new_n359), .C2(new_n629), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n627), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n335), .ZN(new_n635));
  INV_X1    g0435(.A(new_n524), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n561), .A2(G1698), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(G238), .B2(G1698), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n352), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT85), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n630), .A2(new_n631), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n641), .A3(new_n265), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n404), .A3(new_n627), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n635), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n625), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n612), .B1(new_n617), .B2(new_n616), .ZN(new_n646));
  INV_X1    g0446(.A(new_n610), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n619), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(new_n624), .A3(new_n282), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n496), .A2(new_n314), .ZN(new_n650));
  INV_X1    g0450(.A(new_n608), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n642), .A2(new_n327), .A3(new_n627), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n634), .A2(new_n341), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n645), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n606), .A2(new_n656), .ZN(new_n657));
  AND4_X1   g0457(.A1(new_n463), .A2(new_n513), .A3(new_n557), .A4(new_n657), .ZN(G372));
  INV_X1    g0458(.A(new_n343), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n449), .A2(new_n333), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n454), .A2(new_n452), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n453), .B1(new_n434), .B2(G169), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n459), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n411), .A2(new_n412), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n660), .A2(KEYINPUT91), .A3(new_n663), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n415), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n414), .B1(new_n413), .B2(new_n400), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n659), .B1(new_n673), .B2(new_n310), .ZN(new_n674));
  INV_X1    g0474(.A(new_n655), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n579), .B1(new_n593), .B2(new_n590), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n602), .A3(new_n604), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n676), .B1(new_n656), .B2(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n654), .A2(new_n653), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n680), .A2(new_n652), .B1(new_n625), .B2(new_n644), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n601), .A2(new_n605), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(KEYINPUT26), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n675), .B1(new_n679), .B2(new_n683), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n502), .A2(KEYINPUT89), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n498), .A2(new_n501), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n685), .A2(new_n687), .A3(new_n507), .A4(new_n556), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n657), .A2(new_n543), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n463), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n674), .A2(new_n691), .ZN(G369));
  NAND3_X1  g0492(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n510), .A2(new_n699), .ZN(new_n700));
  MUX2_X1   g0500(.A(new_n513), .B(new_n508), .S(new_n700), .Z(new_n701));
  XNOR2_X1  g0501(.A(KEYINPUT92), .B(G330), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n698), .B1(new_n555), .B2(new_n534), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n557), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n556), .B2(new_n699), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n698), .B1(new_n504), .B2(new_n507), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n550), .A2(new_n551), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n530), .B2(new_n535), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n708), .A2(new_n557), .B1(new_n710), .B2(new_n699), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n711), .ZN(G399));
  NOR2_X1   g0512(.A1(new_n228), .A2(G41), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n615), .A2(G116), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(G1), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n716), .B1(new_n236), .B2(new_n714), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT28), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT96), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n681), .A2(new_n543), .A3(new_n678), .A4(new_n594), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n503), .A2(new_n710), .A3(new_n506), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n657), .A2(KEYINPUT96), .A3(new_n543), .A4(new_n688), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n684), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n719), .B1(new_n725), .B2(new_n699), .ZN(new_n726));
  AOI211_X1 g0526(.A(KEYINPUT29), .B(new_n698), .C1(new_n684), .C2(new_n689), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  AND3_X1   g0529(.A1(new_n487), .A2(G179), .A3(new_n575), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT93), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n642), .A2(new_n731), .A3(new_n549), .A4(new_n627), .ZN(new_n732));
  INV_X1    g0532(.A(new_n549), .ZN(new_n733));
  OAI21_X1  g0533(.A(KEYINPUT93), .B1(new_n634), .B2(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n730), .A2(KEYINPUT30), .A3(new_n732), .A4(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n487), .B1(new_n642), .B2(new_n627), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n327), .A3(new_n540), .A4(new_n603), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n327), .B(new_n476), .C1(new_n486), .C2(new_n265), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n734), .A2(new_n739), .A3(new_n575), .A4(new_n732), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT94), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(KEYINPUT94), .A3(new_n741), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n738), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n729), .B1(new_n746), .B2(new_n699), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n557), .A2(new_n678), .A3(new_n681), .A4(new_n594), .ZN(new_n748));
  INV_X1    g0548(.A(new_n512), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n504), .A2(new_n507), .A3(new_n749), .A4(new_n699), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT95), .B1(new_n748), .B2(new_n750), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n735), .A2(new_n737), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n742), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n699), .A2(new_n729), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR4_X1   g0555(.A1(new_n503), .A2(new_n512), .A3(new_n506), .A4(new_n698), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT95), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n756), .A2(new_n657), .A3(new_n757), .A4(new_n557), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n747), .A2(new_n751), .A3(new_n755), .A4(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n702), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n728), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n718), .B1(new_n762), .B2(G1), .ZN(G364));
  NOR2_X1   g0563(.A1(new_n701), .A2(new_n702), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n227), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n206), .B1(new_n765), .B2(G45), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n713), .A2(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n703), .A2(new_n764), .A3(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n701), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n229), .A2(new_n256), .ZN(new_n775));
  INV_X1    g0575(.A(G355), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n775), .A2(new_n776), .B1(G116), .B2(new_n229), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n359), .A2(new_n228), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n236), .B2(G45), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT97), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n779), .A2(new_n780), .B1(new_n251), .B2(G45), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(G20), .B1(KEYINPUT98), .B2(G169), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(KEYINPUT98), .B2(G169), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(new_n232), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n772), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n768), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(G20), .A2(G179), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT99), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G190), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n335), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(new_n404), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n335), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI22_X1  g0597(.A1(new_n215), .A2(new_n794), .B1(new_n797), .B2(new_n440), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n792), .A2(G200), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n798), .B1(G58), .B2(new_n799), .ZN(new_n800));
  NOR4_X1   g0600(.A1(new_n207), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT100), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(KEYINPUT100), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n363), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT32), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n207), .A2(new_n335), .A3(G179), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G190), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n404), .A2(G179), .A3(G200), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n207), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n809), .A2(G87), .B1(new_n812), .B2(G97), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n807), .A2(new_n404), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(G107), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n813), .A2(new_n256), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n795), .A2(G200), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n817), .B1(G77), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n800), .A2(new_n806), .A3(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n793), .A2(G326), .B1(G294), .B2(new_n812), .ZN(new_n821));
  INV_X1    g0621(.A(G311), .ZN(new_n822));
  INV_X1    g0622(.A(new_n818), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT101), .ZN(new_n825));
  INV_X1    g0625(.A(G303), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n484), .B1(new_n808), .B2(new_n826), .C1(new_n827), .C2(new_n814), .ZN(new_n828));
  INV_X1    g0628(.A(new_n804), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n828), .B1(G329), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(KEYINPUT33), .B(G317), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G322), .A2(new_n799), .B1(new_n796), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n820), .B1(new_n825), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n789), .B1(new_n834), .B2(new_n786), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n769), .B1(new_n774), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  AOI21_X1  g0637(.A(new_n698), .B1(new_n684), .B2(new_n689), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n318), .A2(new_n698), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n333), .A2(new_n336), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(KEYINPUT103), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT103), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n333), .A2(new_n842), .A3(new_n336), .A4(new_n839), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n333), .A2(new_n839), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n838), .B(new_n846), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n768), .B1(new_n847), .B2(new_n760), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n760), .B2(new_n847), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n771), .B1(new_n785), .B2(new_n232), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n768), .B1(new_n850), .B2(G77), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G294), .A2(new_n799), .B1(new_n793), .B2(G303), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n852), .B1(new_n211), .B2(new_n823), .C1(new_n827), .C2(new_n797), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n804), .A2(new_n822), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n484), .B1(new_n811), .B2(new_n490), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n815), .A2(G87), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n320), .B2(new_n808), .ZN(new_n857));
  NOR4_X1   g0657(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT102), .Z(new_n859));
  AOI22_X1  g0659(.A1(G143), .A2(new_n799), .B1(new_n796), .B2(G150), .ZN(new_n860));
  INV_X1    g0660(.A(G137), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n860), .B1(new_n861), .B2(new_n794), .C1(new_n363), .C2(new_n823), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT34), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n352), .B1(new_n812), .B2(G58), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n815), .A2(G68), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n866), .B(new_n867), .C1(new_n215), .C2(new_n808), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(G132), .B2(new_n829), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n859), .B1(new_n864), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n851), .B1(new_n871), .B2(new_n786), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n771), .B2(new_n846), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n849), .A2(new_n873), .ZN(G384));
  AOI211_X1 g0674(.A(new_n211), .B(new_n234), .C1(new_n588), .C2(KEYINPUT35), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(KEYINPUT35), .B2(new_n588), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT36), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n370), .A2(G77), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n236), .A2(new_n878), .B1(new_n440), .B2(new_n201), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(G1), .A3(new_n227), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g0681(.A(new_n881), .B(KEYINPUT104), .Z(new_n882));
  NAND3_X1  g0682(.A1(new_n361), .A2(new_n367), .A3(new_n372), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n375), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n346), .B1(new_n374), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n409), .B1(new_n885), .B2(new_n696), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n401), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n413), .A2(new_n400), .ZN(new_n889));
  INV_X1    g0689(.A(new_n696), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n413), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT37), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n889), .A2(new_n891), .A3(new_n892), .A4(new_n409), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n885), .A2(new_n696), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n416), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n894), .A2(new_n896), .A3(KEYINPUT38), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT39), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n889), .A2(new_n891), .A3(new_n409), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  INV_X1    g0700(.A(new_n891), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n893), .A2(new_n900), .B1(new_n416), .B2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n897), .B(new_n898), .C1(KEYINPUT38), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT106), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n894), .A2(new_n896), .A3(KEYINPUT38), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT38), .B1(new_n894), .B2(new_n896), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT39), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n900), .A2(new_n893), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n891), .B1(new_n672), .B2(new_n667), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT106), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(new_n898), .A4(new_n897), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n904), .A2(new_n907), .A3(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n663), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n699), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT107), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n672), .A2(new_n890), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n333), .A2(new_n698), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n921), .B1(new_n838), .B2(new_n846), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n435), .A2(new_n447), .A3(new_n448), .ZN(new_n923));
  INV_X1    g0723(.A(new_n457), .ZN(new_n924));
  INV_X1    g0724(.A(new_n458), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(new_n925), .A3(new_n698), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n663), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  AOI211_X1 g0727(.A(KEYINPUT14), .B(new_n341), .C1(new_n429), .C2(new_n433), .ZN(new_n928));
  INV_X1    g0728(.A(new_n452), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n662), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n926), .B1(new_n930), .B2(new_n923), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n927), .B1(new_n931), .B2(KEYINPUT105), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n457), .A2(new_n458), .A3(new_n699), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n455), .B2(new_n449), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT105), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n922), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n905), .A2(new_n906), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n920), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n918), .A2(new_n919), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n919), .B1(new_n918), .B2(new_n941), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n463), .B1(new_n726), .B2(new_n727), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n674), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  INV_X1    g0748(.A(new_n745), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT94), .B1(new_n740), .B2(new_n741), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n752), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n754), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n747), .A2(new_n751), .A3(new_n758), .A4(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n935), .A2(new_n934), .B1(new_n460), .B2(new_n926), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n931), .A2(KEYINPUT105), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n845), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n948), .B1(new_n957), .B2(new_n939), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n897), .B1(new_n902), .B2(KEYINPUT38), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n959), .A2(new_n956), .A3(new_n953), .A4(KEYINPUT40), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n463), .A2(new_n953), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n963), .A2(new_n702), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n947), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n206), .B2(new_n765), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n947), .A2(new_n965), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n882), .B1(new_n967), .B2(new_n968), .ZN(G367));
  INV_X1    g0769(.A(new_n778), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n787), .B1(new_n229), .B2(new_n314), .C1(new_n247), .C2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT111), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n768), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n815), .A2(G97), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n976), .B(new_n352), .C1(new_n320), .C2(new_n811), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT46), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n808), .B2(new_n211), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n809), .A2(KEYINPUT46), .A3(G116), .ZN(new_n980));
  INV_X1    g0780(.A(G317), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n979), .B(new_n980), .C1(new_n804), .C2(new_n981), .ZN(new_n982));
  AOI211_X1 g0782(.A(new_n977), .B(new_n982), .C1(G303), .C2(new_n799), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G294), .A2(new_n796), .B1(new_n793), .B2(G311), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n983), .B(new_n984), .C1(new_n827), .C2(new_n823), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n812), .A2(G68), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n217), .B2(new_n808), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n484), .B(new_n987), .C1(G77), .C2(new_n815), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n861), .B2(new_n804), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G143), .A2(new_n793), .B1(new_n799), .B2(G150), .ZN(new_n990));
  INV_X1    g0790(.A(new_n201), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n990), .B1(new_n363), .B2(new_n797), .C1(new_n991), .C2(new_n823), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n985), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT47), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n973), .B(new_n975), .C1(new_n994), .C2(new_n786), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n681), .B1(new_n625), .B2(new_n699), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n655), .A2(new_n625), .A3(new_n699), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n995), .B1(new_n773), .B2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n713), .B(KEYINPUT41), .Z(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n708), .A2(new_n557), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n706), .B2(new_n708), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n703), .B(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n762), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n678), .B(new_n594), .C1(new_n601), .C2(new_n699), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n682), .A2(new_n698), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n711), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT45), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n707), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT110), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n711), .A2(new_n1009), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT109), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT44), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(KEYINPUT44), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1014), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1006), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1002), .B1(new_n1023), .B2(new_n761), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n766), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1009), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(new_n1003), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT42), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT42), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n678), .B1(new_n1007), .B2(new_n556), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1028), .A2(new_n1029), .B1(new_n699), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT43), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n998), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT108), .Z(new_n1035));
  XNOR2_X1  g0835(.A(new_n998), .B(KEYINPUT43), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n707), .B2(new_n1026), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1035), .A2(new_n1012), .A3(new_n1009), .A4(new_n1037), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1000), .B1(new_n1025), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(G387));
  OR2_X1    g0844(.A1(new_n706), .A2(new_n773), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n775), .A2(new_n715), .B1(G107), .B2(new_n229), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n243), .A2(G45), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n715), .ZN(new_n1048));
  AOI211_X1 g0848(.A(G45), .B(new_n1048), .C1(G68), .C2(G77), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n312), .A2(new_n215), .ZN(new_n1050));
  XOR2_X1   g0850(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n1051));
  XNOR2_X1  g0851(.A(new_n1050), .B(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n970), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1046), .B1(new_n1047), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n768), .B1(new_n1054), .B2(new_n788), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n809), .A2(G77), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n812), .A2(new_n607), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n976), .A2(new_n1056), .A3(new_n1057), .A4(new_n359), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G150), .B2(new_n829), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G50), .A2(new_n799), .B1(new_n793), .B2(G159), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n289), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1061), .A2(new_n796), .B1(new_n818), .B2(G68), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n829), .A2(G326), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n359), .B1(new_n815), .B2(G116), .ZN(new_n1065));
  INV_X1    g0865(.A(G294), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n808), .A2(new_n1066), .B1(new_n811), .B2(new_n827), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G303), .A2(new_n818), .B1(new_n793), .B2(G322), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n799), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1068), .B1(new_n822), .B2(new_n797), .C1(new_n981), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1067), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n1071), .B2(new_n1070), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT49), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1064), .B(new_n1065), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1063), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1055), .B1(new_n1077), .B2(new_n786), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1005), .A2(new_n767), .B1(new_n1045), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1006), .A2(KEYINPUT113), .A3(new_n713), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n762), .B2(new_n1005), .ZN(new_n1081));
  AOI21_X1  g0881(.A(KEYINPUT113), .B1(new_n1006), .B2(new_n713), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(G393));
  NOR2_X1   g0883(.A1(new_n1023), .A2(new_n714), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1006), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1026), .A2(new_n772), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n787), .B1(new_n490), .B2(new_n229), .C1(new_n254), .C2(new_n970), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n768), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G150), .A2(new_n793), .B1(new_n799), .B2(G159), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT51), .Z(new_n1092));
  NAND2_X1  g0892(.A1(new_n809), .A2(new_n221), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n812), .A2(G77), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n856), .A2(new_n1093), .A3(new_n1094), .A4(new_n359), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G143), .B2(new_n829), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n201), .A2(new_n796), .B1(new_n818), .B2(new_n312), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1092), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n809), .A2(G283), .B1(new_n812), .B2(G116), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(new_n484), .A3(new_n816), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1066), .A2(new_n823), .B1(new_n797), .B2(new_n826), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1100), .B(new_n1101), .C1(G322), .C2(new_n829), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G311), .A2(new_n799), .B1(new_n793), .B2(G317), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT114), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT52), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1104), .A2(KEYINPUT52), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1098), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1090), .B1(new_n1108), .B2(new_n786), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1086), .A2(new_n767), .B1(new_n1088), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1087), .A2(new_n1110), .ZN(G390));
  OAI21_X1  g0911(.A(new_n916), .B1(new_n922), .B2(new_n937), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1112), .A2(new_n904), .A3(new_n907), .A4(new_n913), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n959), .A2(new_n916), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n725), .A2(new_n699), .A3(new_n846), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n921), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT115), .B1(new_n932), .B2(new_n936), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n934), .A2(new_n935), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT115), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n955), .A2(new_n1120), .A3(new_n1121), .A4(new_n927), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1115), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n937), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1125), .A2(new_n759), .A3(new_n702), .A4(new_n846), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1113), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n953), .A2(new_n956), .A3(G330), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n1113), .B2(new_n1124), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n904), .A2(new_n907), .A3(new_n913), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n770), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n768), .B1(new_n1061), .B2(new_n850), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G97), .A2(new_n818), .B1(new_n796), .B2(G107), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1134), .B1(new_n211), .B2(new_n1069), .C1(new_n827), .C2(new_n794), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n829), .A2(G294), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n256), .B1(new_n809), .B2(G87), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1136), .A2(new_n867), .A3(new_n1094), .A4(new_n1137), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT54), .B(G143), .Z(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT117), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n818), .A2(new_n1140), .B1(new_n796), .B2(G137), .ZN(new_n1141));
  INV_X1    g0941(.A(G128), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n794), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n829), .A2(G125), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n808), .A2(new_n293), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n256), .B1(new_n991), .B2(new_n814), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(G159), .B2(new_n812), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n799), .A2(G132), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1135), .A2(new_n1138), .B1(new_n1143), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1133), .B1(new_n1151), .B2(new_n786), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1130), .A2(new_n767), .B1(new_n1132), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1113), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1119), .A2(new_n1122), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1114), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1131), .B2(new_n1112), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1154), .B1(new_n1158), .B2(new_n1128), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n953), .A2(G330), .A3(new_n846), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(new_n1123), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(new_n1118), .A3(new_n1126), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n953), .A2(G330), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n759), .A2(new_n702), .A3(new_n846), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1163), .A2(new_n956), .B1(new_n1164), .B2(new_n937), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1162), .B1(new_n1165), .B2(new_n922), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n463), .A2(G330), .A3(new_n953), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n945), .A2(new_n674), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n714), .B1(new_n1159), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n838), .A2(new_n846), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1117), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1164), .A2(new_n937), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1128), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1168), .B1(new_n1176), .B2(new_n1162), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1177), .B(new_n1154), .C1(new_n1158), .C2(new_n1128), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1171), .A2(KEYINPUT116), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT116), .B1(new_n1171), .B2(new_n1178), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1153), .B1(new_n1179), .B2(new_n1180), .ZN(G378));
  AND2_X1   g0981(.A1(new_n913), .A2(new_n907), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n916), .B1(new_n1182), .B2(new_n904), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1173), .A2(new_n1125), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n1184), .A2(new_n939), .B1(new_n672), .B2(new_n890), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT107), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n918), .A2(new_n941), .A3(new_n919), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n310), .A2(new_n343), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n302), .A3(new_n890), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n302), .A2(new_n890), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n310), .A2(new_n343), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1192), .B(new_n1194), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1195), .A2(G330), .A3(new_n958), .A4(new_n960), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n958), .A2(G330), .A3(new_n960), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1192), .B(new_n1193), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1186), .A2(new_n1187), .A3(new_n1196), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1196), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n942), .B2(new_n943), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1202), .A3(new_n767), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n768), .B1(new_n850), .B2(new_n201), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n1142), .A2(new_n1069), .B1(new_n823), .B2(new_n861), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1140), .A2(new_n809), .B1(G150), .B2(new_n812), .ZN(new_n1206));
  INV_X1    g1006(.A(G132), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n1207), .B2(new_n797), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1205), .B(new_n1208), .C1(G125), .C2(new_n793), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  OR2_X1    g1010(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(KEYINPUT59), .ZN(new_n1212));
  XOR2_X1   g1012(.A(KEYINPUT120), .B(G124), .Z(new_n1213));
  NAND2_X1  g1013(.A1(new_n829), .A2(new_n1213), .ZN(new_n1214));
  AOI211_X1 g1014(.A(G33), .B(G41), .C1(new_n815), .C2(G159), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1211), .A2(new_n1212), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n986), .B1(new_n827), .B2(new_n804), .C1(new_n1069), .C2(new_n320), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1056), .A2(new_n271), .A3(new_n352), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1217), .B1(KEYINPUT119), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(KEYINPUT119), .B2(new_n1218), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n490), .A2(new_n797), .B1(new_n794), .B2(new_n211), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n814), .A2(new_n217), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT118), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n314), .B2(new_n823), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1220), .A2(new_n1221), .A3(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(KEYINPUT58), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(KEYINPUT58), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G50), .B1(new_n347), .B2(new_n271), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n359), .B2(G41), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1216), .A2(new_n1226), .A3(new_n1227), .A4(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1204), .B1(new_n1230), .B2(new_n786), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1195), .B2(new_n771), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1203), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT121), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1233), .B(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT57), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1168), .B1(new_n1130), .B2(new_n1177), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1169), .B1(new_n1159), .B2(new_n1170), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1240), .A2(KEYINPUT57), .A3(new_n1200), .A4(new_n1202), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1239), .A2(new_n713), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1235), .A2(new_n1242), .ZN(G375));
  INV_X1    g1043(.A(KEYINPUT122), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n766), .B1(new_n1176), .B2(new_n1162), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1123), .A2(new_n770), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n768), .B1(new_n850), .B2(G68), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G107), .A2(new_n818), .B1(new_n796), .B2(G116), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n1248), .B1(new_n827), .B2(new_n1069), .C1(new_n1066), .C2(new_n794), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n829), .A2(G303), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n256), .B1(new_n815), .B2(G77), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n809), .A2(G97), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1250), .A2(new_n1057), .A3(new_n1251), .A4(new_n1252), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n796), .A2(new_n1140), .B1(new_n793), .B2(G132), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n293), .B2(new_n823), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n829), .A2(G128), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n359), .B1(new_n808), .B2(new_n363), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G50), .B2(new_n812), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n799), .A2(G137), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1256), .A2(new_n1223), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1249), .A2(new_n1253), .B1(new_n1255), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1247), .B1(new_n1261), .B2(new_n786), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1246), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1244), .B1(new_n1245), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1166), .A2(new_n767), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(KEYINPUT122), .A3(new_n1263), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1162), .B(new_n1168), .C1(new_n1165), .C2(new_n922), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1170), .A2(new_n1002), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1268), .A2(new_n1270), .ZN(G381));
  NAND2_X1  g1071(.A1(new_n1171), .A2(new_n1178), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1272), .A2(new_n1153), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(G387), .A2(G390), .A3(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G375), .ZN(new_n1276));
  NOR4_X1   g1076(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1278), .A2(KEYINPUT123), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(KEYINPUT123), .ZN(new_n1280));
  OR2_X1    g1080(.A1(new_n1279), .A2(new_n1280), .ZN(G407));
  NAND2_X1  g1081(.A1(new_n1273), .A2(new_n697), .ZN(new_n1282));
  OAI221_X1 g1082(.A(G213), .B1(G375), .B2(new_n1282), .C1(new_n1279), .C2(new_n1280), .ZN(G409));
  INV_X1    g1083(.A(KEYINPUT126), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1087), .A2(new_n1110), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1284), .B1(new_n1285), .B2(new_n1043), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(G393), .B(G396), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1041), .B1(new_n1024), .B2(new_n766), .ZN(new_n1288));
  OAI21_X1  g1088(.A(G390), .B1(new_n1288), .B2(new_n1000), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1286), .A2(new_n1287), .A3(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1287), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT121), .B1(new_n1203), .B2(new_n1232), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1242), .B(G378), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1240), .A2(new_n1002), .A3(new_n1200), .A4(new_n1202), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT124), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1299), .A2(KEYINPUT124), .A3(new_n1002), .A4(new_n1240), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1203), .A2(new_n1232), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1298), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1273), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1295), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(G213), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1305), .A2(G343), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1304), .A2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n714), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT60), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1269), .A2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1176), .A2(KEYINPUT60), .A3(new_n1168), .A4(new_n1162), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1309), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(KEYINPUT122), .B1(new_n1266), .B2(new_n1263), .ZN(new_n1314));
  AOI211_X1 g1114(.A(new_n1244), .B(new_n1264), .C1(new_n1166), .C2(new_n767), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1313), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(G384), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1268), .A2(G384), .A3(new_n1313), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(KEYINPUT125), .A3(new_n1319), .ZN(new_n1320));
  AND2_X1   g1120(.A1(new_n1306), .A2(G2897), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT125), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1319), .ZN(new_n1324));
  AOI21_X1  g1124(.A(G384), .B1(new_n1268), .B2(new_n1313), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1323), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1322), .A2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1323), .B(new_n1321), .C1(new_n1324), .C2(new_n1325), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT61), .B1(new_n1308), .B2(new_n1329), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1304), .A2(new_n1307), .A3(new_n1331), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1332), .A2(KEYINPUT63), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(KEYINPUT63), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1292), .B(new_n1330), .C1(new_n1333), .C2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(new_n1291), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1286), .A2(new_n1287), .A3(new_n1289), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT61), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1306), .B1(new_n1295), .B2(new_n1303), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1339), .B1(new_n1340), .B2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT62), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1332), .A2(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1340), .A2(KEYINPUT62), .A3(new_n1331), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1342), .B1(new_n1344), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT127), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1338), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1345), .ZN(new_n1349));
  AOI21_X1  g1149(.A(KEYINPUT62), .B1(new_n1340), .B2(new_n1331), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n1347), .B(new_n1330), .C1(new_n1349), .C2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1351), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1335), .B1(new_n1348), .B2(new_n1352), .ZN(G405));
  NAND2_X1  g1153(.A1(G375), .A2(new_n1273), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(new_n1295), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1355), .B(new_n1331), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(new_n1338), .B(new_n1356), .ZN(G402));
endmodule


