//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1120, new_n1121;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT67), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT70), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n468), .A2(new_n469), .A3(G125), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT69), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n460), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G101), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n468), .ZN(new_n481));
  INV_X1    g056(.A(G137), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G160));
  NOR2_X1   g061(.A1(new_n476), .A2(new_n464), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OAI221_X1 g063(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n476), .C2(G112), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n464), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n488), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  NAND3_X1  g068(.A1(new_n476), .A2(new_n468), .A3(G138), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n476), .A2(new_n468), .A3(new_n496), .A4(G138), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  INV_X1    g074(.A(G126), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n464), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G2105), .B1(G102), .B2(new_n479), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT71), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n498), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(G164));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT72), .A3(G50), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n519), .A2(new_n508), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n510), .A2(new_n514), .B1(G88), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n521), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n508), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G63), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n531), .B2(new_n523), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(new_n519), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n509), .A2(KEYINPUT73), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n512), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G51), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n533), .B(new_n535), .C1(new_n539), .C2(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  AND3_X1   g117(.A1(new_n536), .A2(G52), .A3(new_n538), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n519), .A2(new_n508), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n544), .A2(new_n523), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n543), .A2(new_n547), .ZN(G171));
  AND3_X1   g123(.A1(new_n536), .A2(G43), .A3(new_n538), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n550), .A2(new_n523), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n509), .A2(G53), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n520), .A2(G91), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n519), .B(KEYINPUT75), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n561), .B(new_n562), .C1(new_n564), .C2(new_n523), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  NAND3_X1  g141(.A1(new_n508), .A2(G49), .A3(G543), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT76), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n520), .A2(G87), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  NAND2_X1  g146(.A1(new_n520), .A2(G86), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n516), .A2(new_n518), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n509), .A2(G48), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n572), .A2(new_n577), .A3(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n580), .A2(new_n523), .B1(new_n581), .B2(new_n545), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n536), .A2(new_n538), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n582), .B1(new_n583), .B2(G47), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n583), .A2(KEYINPUT78), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n539), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(G54), .A3(new_n589), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n563), .A2(G66), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT79), .Z(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n520), .A2(G92), .ZN(new_n595));
  XOR2_X1   g170(.A(KEYINPUT77), .B(KEYINPUT10), .Z(new_n596));
  XNOR2_X1  g171(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n590), .A2(new_n594), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT80), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n586), .B1(new_n600), .B2(G868), .ZN(G284));
  XNOR2_X1  g176(.A(G284), .B(KEYINPUT81), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n600), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n490), .A2(G2104), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n487), .A2(G123), .ZN(new_n617));
  OAI221_X1 g192(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n476), .C2(G111), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n490), .A2(G135), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n616), .A2(new_n621), .ZN(G156));
  XNOR2_X1  g197(.A(G2451), .B(G2454), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT16), .ZN(new_n624));
  XNOR2_X1  g199(.A(G2443), .B(G2446), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n626), .B(new_n627), .Z(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2435), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2438), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n628), .B(new_n633), .ZN(new_n634));
  AND2_X1   g209(.A1(new_n634), .A2(G14), .ZN(G401));
  XOR2_X1   g210(.A(G2067), .B(G2678), .Z(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2084), .B(G2090), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n639), .A2(KEYINPUT17), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  AOI21_X1  g216(.A(KEYINPUT18), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2072), .B(G2078), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT82), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(KEYINPUT18), .B2(new_n639), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n642), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2096), .B(G2100), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(G227));
  XNOR2_X1  g223(.A(G1971), .B(G1976), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT19), .ZN(new_n650));
  XOR2_X1   g225(.A(G1956), .B(G2474), .Z(new_n651));
  XOR2_X1   g226(.A(G1961), .B(G1966), .Z(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n650), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n651), .A2(new_n652), .ZN(new_n656));
  AOI22_X1  g231(.A1(new_n654), .A2(KEYINPUT20), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n658), .A2(new_n650), .A3(new_n653), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n657), .B(new_n659), .C1(KEYINPUT20), .C2(new_n654), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT84), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1991), .B(G1996), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT83), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n661), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(G229));
  INV_X1    g243(.A(G16), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(G24), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(new_n584), .B2(new_n669), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n671), .A2(G1986), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(G1986), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT36), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n672), .B(new_n673), .C1(KEYINPUT86), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(G22), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(G166), .B2(new_n669), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1971), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n669), .A2(G23), .ZN(new_n679));
  INV_X1    g254(.A(G288), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n679), .B1(new_n680), .B2(new_n669), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT33), .Z(new_n682));
  AOI21_X1  g257(.A(new_n678), .B1(new_n682), .B2(G1976), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n669), .A2(G6), .ZN(new_n684));
  INV_X1    g259(.A(G305), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n669), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT32), .B(G1981), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n683), .B(new_n688), .C1(G1976), .C2(new_n682), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n675), .B1(new_n689), .B2(KEYINPUT34), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G25), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n487), .A2(G119), .ZN(new_n693));
  OAI221_X1 g268(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n476), .C2(G107), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n490), .A2(G131), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n692), .B1(new_n697), .B2(new_n691), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT35), .B(G1991), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT85), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n690), .B(new_n701), .C1(KEYINPUT34), .C2(new_n689), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n674), .A2(KEYINPUT86), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n691), .A2(G35), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G162), .B2(new_n691), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT29), .B(G2090), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n702), .A2(new_n703), .ZN(new_n709));
  NAND2_X1  g284(.A1(G168), .A2(G16), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G16), .B2(G21), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT92), .B(G1966), .Z(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(G171), .A2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G5), .B2(G16), .ZN(new_n715));
  INV_X1    g290(.A(G1961), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n711), .A2(new_n712), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n620), .A2(new_n691), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT93), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT30), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n691), .B1(new_n721), .B2(G28), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n721), .B2(G28), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n713), .A2(new_n717), .A3(new_n718), .A4(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT31), .B(G11), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n715), .A2(new_n716), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n669), .A2(G19), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(new_n553), .B2(new_n669), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(G1341), .ZN(new_n730));
  OR2_X1    g305(.A1(G29), .A2(G33), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT25), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n490), .A2(G139), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n733), .B(new_n734), .C1(new_n476), .C2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n731), .B1(new_n736), .B2(new_n691), .ZN(new_n737));
  INV_X1    g312(.A(G2072), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n729), .A2(G1341), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n727), .A2(new_n730), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n725), .A2(new_n726), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n669), .A2(G20), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT95), .Z(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT23), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G299), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1956), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n737), .A2(new_n738), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT88), .ZN(new_n749));
  AND2_X1   g324(.A1(KEYINPUT24), .A2(G34), .ZN(new_n750));
  NOR2_X1   g325(.A1(KEYINPUT24), .A2(G34), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n750), .A2(new_n751), .A3(G29), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n485), .B2(G29), .ZN(new_n753));
  INV_X1    g328(.A(G2084), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT28), .ZN(new_n756));
  INV_X1    g331(.A(G26), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G29), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(G29), .ZN(new_n759));
  AOI22_X1  g334(.A1(G128), .A2(new_n487), .B1(new_n490), .B2(G140), .ZN(new_n760));
  OAI221_X1 g335(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n476), .C2(G116), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n759), .B1(new_n762), .B2(G29), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n758), .B1(new_n763), .B2(new_n756), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n755), .B1(G2067), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G2067), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n753), .A2(new_n754), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT94), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n742), .A2(new_n747), .A3(new_n749), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G4), .A2(G16), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n600), .B2(G16), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT87), .B(G1348), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G27), .A2(G29), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(G164), .B2(G29), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2078), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n479), .A2(G105), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT89), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n487), .A2(G129), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT26), .Z(new_n782));
  NAND2_X1  g357(.A1(new_n490), .A2(G141), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n779), .A2(new_n780), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT90), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n785), .A2(KEYINPUT91), .A3(G29), .ZN(new_n786));
  AOI21_X1  g361(.A(KEYINPUT91), .B1(new_n785), .B2(G29), .ZN(new_n787));
  OAI22_X1  g362(.A1(new_n786), .A2(new_n787), .B1(G29), .B2(G32), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT27), .B(G1996), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n770), .A2(new_n774), .A3(new_n777), .A4(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n704), .A2(new_n708), .A3(new_n709), .A4(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(G311));
  XOR2_X1   g368(.A(new_n792), .B(KEYINPUT96), .Z(G150));
  AND2_X1   g369(.A1(new_n583), .A2(G55), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT97), .B(G93), .ZN(new_n797));
  OAI22_X1  g372(.A1(new_n796), .A2(new_n523), .B1(new_n545), .B2(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G860), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT37), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n553), .ZN(new_n802));
  OR3_X1    g377(.A1(new_n795), .A2(new_n553), .A3(new_n798), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT38), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n600), .A2(G559), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(KEYINPUT39), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT98), .ZN(new_n809));
  AOI21_X1  g384(.A(G860), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n809), .B2(new_n808), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n807), .A2(KEYINPUT39), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n801), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT99), .Z(G145));
  NAND2_X1  g389(.A1(new_n736), .A2(new_n784), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n785), .B(KEYINPUT101), .Z(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(new_n736), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(new_n620), .Z(new_n818));
  AOI22_X1  g393(.A1(G130), .A2(new_n487), .B1(new_n490), .B2(G142), .ZN(new_n819));
  OAI221_X1 g394(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n476), .C2(G118), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n614), .B(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n762), .B(KEYINPUT100), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n503), .B(new_n696), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n818), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n818), .A2(new_n826), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n485), .B(new_n492), .ZN(new_n829));
  OR3_X1    g404(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(G37), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n827), .B2(new_n828), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g409(.A1(new_n799), .A2(G868), .ZN(new_n835));
  INV_X1    g410(.A(new_n804), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n600), .A2(new_n607), .A3(new_n804), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n590), .A2(new_n594), .A3(new_n597), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(G299), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n598), .A2(new_n604), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT41), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n841), .A2(KEYINPUT41), .A3(new_n842), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT102), .B1(new_n839), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n839), .A2(new_n843), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n837), .A2(new_n847), .A3(new_n851), .A4(new_n838), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(G303), .B(new_n685), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n584), .B(G288), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n856), .B1(new_n857), .B2(KEYINPUT103), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(KEYINPUT103), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT42), .Z(new_n861));
  NAND4_X1  g436(.A1(new_n849), .A2(KEYINPUT104), .A3(new_n850), .A4(new_n852), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n855), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n861), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n864), .A2(new_n853), .A3(new_n854), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n835), .B1(new_n866), .B2(G868), .ZN(G331));
  XNOR2_X1  g442(.A(G331), .B(KEYINPUT105), .ZN(G295));
  INV_X1    g443(.A(KEYINPUT110), .ZN(new_n869));
  XNOR2_X1  g444(.A(G168), .B(G171), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n804), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT107), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n802), .A3(new_n803), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n836), .A2(KEYINPUT107), .A3(new_n870), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n875), .A2(new_n876), .B1(new_n842), .B2(new_n841), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT108), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n836), .A2(new_n880), .A3(new_n870), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n872), .A2(new_n880), .A3(new_n874), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n847), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n860), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n875), .A2(new_n876), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n843), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n878), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n877), .A2(KEYINPUT108), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n888), .A2(new_n860), .A3(new_n884), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n831), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT43), .B1(new_n885), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n883), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n843), .B1(new_n893), .B2(new_n881), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT109), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n847), .A2(new_n876), .A3(new_n875), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT109), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n897), .B(new_n843), .C1(new_n893), .C2(new_n881), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n860), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n831), .A4(new_n890), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n892), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n869), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI211_X1 g481(.A(KEYINPUT110), .B(KEYINPUT44), .C1(new_n892), .C2(new_n903), .ZN(new_n907));
  NOR3_X1   g482(.A1(new_n885), .A2(new_n891), .A3(KEYINPUT43), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n891), .B1(new_n900), .B2(new_n899), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT44), .B1(new_n909), .B2(new_n902), .ZN(new_n910));
  OAI22_X1  g485(.A1(new_n906), .A2(new_n907), .B1(new_n908), .B2(new_n910), .ZN(G397));
  NAND2_X1  g486(.A1(G305), .A2(G1981), .ZN(new_n912));
  INV_X1    g487(.A(G1981), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n572), .A2(new_n913), .A3(new_n577), .A4(new_n578), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(KEYINPUT49), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G8), .ZN(new_n916));
  INV_X1    g491(.A(G40), .ZN(new_n917));
  AOI211_X1 g492(.A(new_n917), .B(new_n483), .C1(new_n477), .C2(new_n471), .ZN(new_n918));
  AOI21_X1  g493(.A(G1384), .B1(new_n498), .B2(new_n502), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n912), .A2(new_n914), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT49), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT113), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT113), .ZN(new_n924));
  AOI211_X1 g499(.A(new_n924), .B(KEYINPUT49), .C1(new_n912), .C2(new_n914), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n915), .B(new_n920), .C1(new_n923), .C2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(G1976), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT52), .B1(G288), .B2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n920), .B(new_n928), .C1(new_n927), .C2(G288), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n920), .B1(new_n927), .B2(G288), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT52), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n926), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n498), .A2(new_n505), .A3(new_n502), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n505), .B1(new_n498), .B2(new_n502), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n934), .A2(new_n935), .A3(G1384), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT50), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G2090), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n478), .A2(G40), .A3(new_n484), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n937), .B2(new_n919), .ZN(new_n941));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n504), .A2(new_n942), .A3(new_n506), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n938), .A2(new_n939), .A3(new_n941), .A4(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n940), .B1(KEYINPUT45), .B2(new_n919), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(new_n936), .B2(KEYINPUT45), .ZN(new_n947));
  INV_X1    g522(.A(G1971), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n916), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n951));
  OR2_X1    g526(.A1(new_n951), .A2(KEYINPUT112), .ZN(new_n952));
  NAND3_X1  g527(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(KEYINPUT112), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n932), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n955), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n504), .A2(new_n937), .A3(new_n942), .A4(new_n506), .ZN(new_n958));
  INV_X1    g533(.A(new_n919), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT50), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n958), .A2(new_n960), .A3(new_n939), .A4(new_n918), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n918), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n943), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT116), .B(new_n961), .C1(new_n965), .C2(G1971), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(G8), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT116), .B1(new_n949), .B2(new_n961), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n957), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n938), .A2(new_n754), .A3(new_n941), .A4(new_n944), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n940), .B1(new_n959), .B2(new_n964), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n971), .B1(new_n943), .B2(new_n964), .ZN(new_n972));
  INV_X1    g547(.A(G1966), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n916), .B(G286), .C1(new_n970), .C2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n956), .A2(new_n969), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT117), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT63), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT117), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n956), .A2(new_n969), .A3(new_n979), .A4(new_n975), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n950), .A2(new_n955), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n970), .A2(new_n974), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(G8), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n982), .A2(G286), .A3(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(new_n932), .B(KEYINPUT114), .Z(new_n986));
  NAND2_X1  g561(.A1(new_n950), .A2(new_n955), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT63), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n981), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n926), .A2(new_n927), .A3(new_n680), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n914), .ZN(new_n991));
  XOR2_X1   g566(.A(new_n991), .B(KEYINPUT115), .Z(new_n992));
  INV_X1    g567(.A(new_n987), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n992), .A2(new_n920), .B1(new_n993), .B2(new_n986), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n971), .A2(KEYINPUT123), .B1(KEYINPUT45), .B2(new_n919), .ZN(new_n995));
  INV_X1    g570(.A(G2078), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT53), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n918), .B1(KEYINPUT45), .B2(new_n919), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT123), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AND3_X1   g575(.A1(new_n995), .A2(new_n1000), .A3(KEYINPUT124), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT124), .B1(new_n995), .B2(new_n1000), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n938), .A2(new_n941), .A3(new_n944), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n716), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n996), .B(new_n946), .C1(new_n936), .C2(KEYINPUT45), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT122), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT122), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1003), .A2(new_n1005), .A3(new_n1009), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(G171), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1005), .A2(new_n1011), .A3(new_n1009), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT125), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n972), .A2(new_n997), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1014), .A2(new_n1015), .A3(G301), .A4(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1005), .A2(new_n1011), .A3(new_n1016), .A4(new_n1009), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT125), .B1(new_n1018), .B2(G171), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1013), .A2(new_n1017), .A3(KEYINPUT54), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n918), .A2(new_n919), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(G2067), .ZN(new_n1022));
  INV_X1    g597(.A(G1348), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1004), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(new_n598), .ZN(new_n1025));
  AOI211_X1 g600(.A(new_n840), .B(new_n1022), .C1(new_n1004), .C2(new_n1023), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT60), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g602(.A(KEYINPUT60), .B(new_n1022), .C1(new_n1004), .C2(new_n1023), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT61), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n958), .A2(new_n918), .A3(new_n960), .ZN(new_n1030));
  INV_X1    g605(.A(G1956), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT56), .B(G2072), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n946), .B(new_n1033), .C1(new_n936), .C2(KEYINPUT45), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(G299), .B(KEYINPUT57), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1029), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n965), .A2(new_n1033), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1036), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1028), .A2(new_n840), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n553), .ZN(new_n1042));
  INV_X1    g617(.A(G1996), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n965), .A2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT58), .B(G1341), .Z(new_n1045));
  NAND2_X1  g620(.A1(new_n1021), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1042), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1027), .A2(new_n1041), .A3(new_n1049), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1035), .A2(KEYINPUT118), .A3(new_n1036), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT119), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n1025), .A2(new_n1055), .B1(new_n1036), .B2(new_n1035), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT119), .B1(new_n1024), .B2(new_n598), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1054), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1020), .B1(new_n1050), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1018), .A2(G171), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1060), .B1(new_n1012), .B2(G171), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(G286), .A2(G8), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT51), .B1(new_n1064), .B2(KEYINPUT120), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n984), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n983), .A2(G8), .A3(G286), .ZN(new_n1068));
  OAI211_X1 g643(.A(G8), .B(new_n1065), .C1(new_n983), .C2(G286), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1029), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1071), .A2(new_n956), .A3(new_n969), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1063), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n989), .B(new_n994), .C1(new_n1059), .C2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT126), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(new_n1060), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1077), .A2(new_n956), .A3(new_n969), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1025), .A2(new_n1055), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n1057), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1054), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1027), .A2(new_n1041), .A3(new_n1049), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AND4_X1   g661(.A1(new_n956), .A2(new_n1070), .A3(new_n969), .A4(new_n1071), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1086), .A2(new_n1087), .A3(new_n1020), .A4(new_n1063), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT126), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n994), .A4(new_n989), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1075), .A2(new_n1079), .A3(new_n1090), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n940), .A2(new_n919), .A3(KEYINPUT45), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n785), .A2(new_n1043), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n784), .A2(G1996), .ZN(new_n1094));
  XOR2_X1   g669(.A(new_n762), .B(G2067), .Z(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n697), .A2(new_n700), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n697), .A2(new_n700), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1986), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n584), .B(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1092), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1091), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1092), .A2(new_n1043), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1105), .A2(KEYINPUT46), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(KEYINPUT46), .ZN(new_n1107));
  INV_X1    g682(.A(new_n784), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1095), .A2(new_n1108), .ZN(new_n1109));
  AOI22_X1  g684(.A1(new_n1106), .A2(new_n1107), .B1(new_n1092), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(KEYINPUT47), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1092), .A2(new_n1101), .A3(new_n584), .ZN(new_n1112));
  XOR2_X1   g687(.A(new_n1112), .B(KEYINPUT127), .Z(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(KEYINPUT48), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1092), .B2(new_n1100), .ZN(new_n1115));
  OAI22_X1  g690(.A1(new_n1096), .A2(new_n1099), .B1(G2067), .B2(new_n762), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n1111), .B(new_n1115), .C1(new_n1092), .C2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1104), .A2(new_n1117), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g693(.A1(G227), .A2(new_n458), .ZN(new_n1120));
  NOR2_X1   g694(.A1(G229), .A2(G401), .ZN(new_n1121));
  NAND4_X1  g695(.A1(new_n904), .A2(new_n833), .A3(new_n1120), .A4(new_n1121), .ZN(G225));
  INV_X1    g696(.A(G225), .ZN(G308));
endmodule


