

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U549 ( .A1(n541), .A2(n540), .ZN(n542) );
  BUF_X2 U550 ( .A(n894), .Z(n515) );
  NAND2_X1 U551 ( .A1(n692), .A2(n785), .ZN(n748) );
  XNOR2_X1 U552 ( .A(n691), .B(KEYINPUT64), .ZN(n785) );
  BUF_X1 U553 ( .A(n608), .Z(n609) );
  AND2_X1 U554 ( .A1(n536), .A2(n535), .ZN(n894) );
  XNOR2_X1 U555 ( .A(KEYINPUT32), .B(KEYINPUT104), .ZN(n755) );
  NOR2_X1 U556 ( .A1(n762), .A2(n779), .ZN(n516) );
  NOR2_X2 U557 ( .A1(n536), .A2(n535), .ZN(n890) );
  XNOR2_X1 U558 ( .A(n704), .B(KEYINPUT31), .ZN(n705) );
  XNOR2_X1 U559 ( .A(n706), .B(n705), .ZN(n742) );
  NOR2_X1 U560 ( .A1(G651), .A2(n630), .ZN(n655) );
  NOR2_X1 U561 ( .A1(G543), .A2(G651), .ZN(n651) );
  NAND2_X1 U562 ( .A1(G89), .A2(n651), .ZN(n517) );
  XNOR2_X1 U563 ( .A(n517), .B(KEYINPUT74), .ZN(n518) );
  XNOR2_X1 U564 ( .A(n518), .B(KEYINPUT4), .ZN(n520) );
  XOR2_X1 U565 ( .A(G543), .B(KEYINPUT0), .Z(n630) );
  INV_X1 U566 ( .A(G651), .ZN(n522) );
  NOR2_X1 U567 ( .A1(n630), .A2(n522), .ZN(n649) );
  NAND2_X1 U568 ( .A1(G76), .A2(n649), .ZN(n519) );
  NAND2_X1 U569 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U570 ( .A(n521), .B(KEYINPUT5), .ZN(n528) );
  NAND2_X1 U571 ( .A1(G51), .A2(n655), .ZN(n525) );
  NOR2_X1 U572 ( .A1(G543), .A2(n522), .ZN(n523) );
  XOR2_X1 U573 ( .A(KEYINPUT1), .B(n523), .Z(n656) );
  NAND2_X1 U574 ( .A1(G63), .A2(n656), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U576 ( .A(KEYINPUT6), .B(n526), .Z(n527) );
  NAND2_X1 U577 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U578 ( .A(n529), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U579 ( .A(G168), .B(KEYINPUT8), .ZN(n530) );
  XNOR2_X1 U580 ( .A(n530), .B(KEYINPUT75), .ZN(G286) );
  XOR2_X1 U581 ( .A(KEYINPUT65), .B(G2104), .Z(n536) );
  INV_X1 U582 ( .A(G2105), .ZN(n535) );
  NAND2_X1 U583 ( .A1(G102), .A2(n894), .ZN(n533) );
  NOR2_X1 U584 ( .A1(G2105), .A2(G2104), .ZN(n531) );
  XOR2_X1 U585 ( .A(KEYINPUT17), .B(n531), .Z(n608) );
  NAND2_X1 U586 ( .A1(G138), .A2(n608), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U588 ( .A(n534), .B(KEYINPUT87), .ZN(n541) );
  NAND2_X1 U589 ( .A1(G126), .A2(n890), .ZN(n539) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  NAND2_X1 U591 ( .A1(n889), .A2(G114), .ZN(n537) );
  XNOR2_X1 U592 ( .A(KEYINPUT86), .B(n537), .ZN(n538) );
  AND2_X1 U593 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U594 ( .A(n542), .B(KEYINPUT88), .ZN(n690) );
  BUF_X1 U595 ( .A(n690), .Z(G164) );
  XNOR2_X1 U596 ( .A(G2427), .B(KEYINPUT109), .ZN(n552) );
  XOR2_X1 U597 ( .A(G2443), .B(G2438), .Z(n544) );
  XNOR2_X1 U598 ( .A(G2430), .B(G2454), .ZN(n543) );
  XNOR2_X1 U599 ( .A(n544), .B(n543), .ZN(n548) );
  XOR2_X1 U600 ( .A(KEYINPUT108), .B(G2435), .Z(n546) );
  INV_X1 U601 ( .A(G1341), .ZN(n994) );
  XOR2_X1 U602 ( .A(n994), .B(G1348), .Z(n545) );
  XNOR2_X1 U603 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U604 ( .A(n548), .B(n547), .Z(n550) );
  XNOR2_X1 U605 ( .A(G2451), .B(G2446), .ZN(n549) );
  XNOR2_X1 U606 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U607 ( .A(n552), .B(n551), .ZN(n553) );
  AND2_X1 U608 ( .A1(n553), .A2(G14), .ZN(G401) );
  AND2_X1 U609 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U610 ( .A(G57), .ZN(G237) );
  INV_X1 U611 ( .A(G108), .ZN(G238) );
  INV_X1 U612 ( .A(G120), .ZN(G236) );
  INV_X1 U613 ( .A(G132), .ZN(G219) );
  INV_X1 U614 ( .A(G82), .ZN(G220) );
  NAND2_X1 U615 ( .A1(G137), .A2(n608), .ZN(n554) );
  XNOR2_X1 U616 ( .A(n554), .B(KEYINPUT66), .ZN(n557) );
  NAND2_X1 U617 ( .A1(G101), .A2(n515), .ZN(n555) );
  XOR2_X1 U618 ( .A(KEYINPUT23), .B(n555), .Z(n556) );
  NAND2_X1 U619 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G113), .A2(n889), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G125), .A2(n890), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U623 ( .A1(n561), .A2(n560), .ZN(G160) );
  NAND2_X1 U624 ( .A1(G77), .A2(n649), .ZN(n563) );
  NAND2_X1 U625 ( .A1(G90), .A2(n651), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U627 ( .A(KEYINPUT9), .B(n564), .ZN(n568) );
  NAND2_X1 U628 ( .A1(G52), .A2(n655), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G64), .A2(n656), .ZN(n565) );
  AND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n568), .A2(n567), .ZN(G301) );
  INV_X1 U632 ( .A(G301), .ZN(G171) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n569) );
  XOR2_X1 U634 ( .A(n569), .B(KEYINPUT10), .Z(n837) );
  NAND2_X1 U635 ( .A1(n837), .A2(G567), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U637 ( .A1(n656), .A2(G56), .ZN(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT14), .B(n571), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n651), .A2(G81), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G68), .A2(n649), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U643 ( .A(KEYINPUT13), .B(n575), .ZN(n576) );
  NAND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n578), .B(KEYINPUT71), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n655), .A2(G43), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n975) );
  INV_X1 U648 ( .A(G860), .ZN(n624) );
  NOR2_X1 U649 ( .A1(n975), .A2(n624), .ZN(n581) );
  XOR2_X1 U650 ( .A(KEYINPUT72), .B(n581), .Z(G153) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U652 ( .A1(G79), .A2(n649), .ZN(n583) );
  NAND2_X1 U653 ( .A1(G54), .A2(n655), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n588) );
  NAND2_X1 U655 ( .A1(G66), .A2(n656), .ZN(n585) );
  NAND2_X1 U656 ( .A1(G92), .A2(n651), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U658 ( .A(KEYINPUT73), .B(n586), .Z(n587) );
  NOR2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U660 ( .A(KEYINPUT15), .B(n589), .Z(n970) );
  INV_X1 U661 ( .A(n970), .ZN(n730) );
  INV_X1 U662 ( .A(G868), .ZN(n670) );
  NAND2_X1 U663 ( .A1(n730), .A2(n670), .ZN(n590) );
  NAND2_X1 U664 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U665 ( .A1(G78), .A2(n649), .ZN(n592) );
  XNOR2_X1 U666 ( .A(n592), .B(KEYINPUT70), .ZN(n599) );
  NAND2_X1 U667 ( .A1(G53), .A2(n655), .ZN(n594) );
  NAND2_X1 U668 ( .A1(G65), .A2(n656), .ZN(n593) );
  NAND2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U670 ( .A1(G91), .A2(n651), .ZN(n595) );
  XNOR2_X1 U671 ( .A(KEYINPUT69), .B(n595), .ZN(n596) );
  NOR2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U673 ( .A1(n599), .A2(n598), .ZN(G299) );
  NOR2_X1 U674 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U675 ( .A1(G286), .A2(n670), .ZN(n600) );
  NOR2_X1 U676 ( .A1(n601), .A2(n600), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n624), .A2(G559), .ZN(n602) );
  NAND2_X1 U678 ( .A1(n602), .A2(n970), .ZN(n603) );
  XNOR2_X1 U679 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n975), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n970), .A2(G868), .ZN(n604) );
  NOR2_X1 U682 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U683 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U684 ( .A1(G123), .A2(n890), .ZN(n607) );
  XNOR2_X1 U685 ( .A(n607), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n609), .A2(G135), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U688 ( .A1(G99), .A2(n515), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G111), .A2(n889), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n925) );
  XNOR2_X1 U692 ( .A(n925), .B(G2096), .ZN(n616) );
  INV_X1 U693 ( .A(G2100), .ZN(n846) );
  NAND2_X1 U694 ( .A1(n616), .A2(n846), .ZN(G156) );
  NAND2_X1 U695 ( .A1(G55), .A2(n655), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G67), .A2(n656), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G80), .A2(n649), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G93), .A2(n651), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  OR2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n671) );
  XNOR2_X1 U702 ( .A(n671), .B(KEYINPUT76), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G559), .A2(n970), .ZN(n623) );
  XOR2_X1 U704 ( .A(n975), .B(n623), .Z(n667) );
  NAND2_X1 U705 ( .A1(n667), .A2(n624), .ZN(n625) );
  XNOR2_X1 U706 ( .A(n626), .B(n625), .ZN(G145) );
  NAND2_X1 U707 ( .A1(G49), .A2(n655), .ZN(n628) );
  NAND2_X1 U708 ( .A1(G74), .A2(G651), .ZN(n627) );
  NAND2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U710 ( .A1(n656), .A2(n629), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n630), .A2(G87), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U713 ( .A1(G48), .A2(n655), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G61), .A2(n656), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n638) );
  XOR2_X1 U716 ( .A(KEYINPUT2), .B(KEYINPUT77), .Z(n636) );
  NAND2_X1 U717 ( .A1(n649), .A2(G73), .ZN(n635) );
  XOR2_X1 U718 ( .A(n636), .B(n635), .Z(n637) );
  NOR2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n651), .A2(G86), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G88), .A2(n651), .ZN(n647) );
  NAND2_X1 U723 ( .A1(G75), .A2(n649), .ZN(n642) );
  NAND2_X1 U724 ( .A1(G50), .A2(n655), .ZN(n641) );
  NAND2_X1 U725 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n656), .A2(G62), .ZN(n643) );
  XOR2_X1 U727 ( .A(KEYINPUT78), .B(n643), .Z(n644) );
  NOR2_X1 U728 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U729 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U730 ( .A(n648), .B(KEYINPUT79), .ZN(G166) );
  NAND2_X1 U731 ( .A1(n649), .A2(G72), .ZN(n650) );
  XOR2_X1 U732 ( .A(KEYINPUT67), .B(n650), .Z(n653) );
  NAND2_X1 U733 ( .A1(n651), .A2(G85), .ZN(n652) );
  NAND2_X1 U734 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U735 ( .A(KEYINPUT68), .B(n654), .Z(n660) );
  NAND2_X1 U736 ( .A1(G47), .A2(n655), .ZN(n658) );
  NAND2_X1 U737 ( .A1(G60), .A2(n656), .ZN(n657) );
  AND2_X1 U738 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U739 ( .A1(n660), .A2(n659), .ZN(G290) );
  XNOR2_X1 U740 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n662) );
  XOR2_X1 U741 ( .A(G288), .B(G299), .Z(n661) );
  XNOR2_X1 U742 ( .A(n662), .B(n661), .ZN(n663) );
  XOR2_X1 U743 ( .A(n671), .B(n663), .Z(n665) );
  XNOR2_X1 U744 ( .A(G305), .B(G166), .ZN(n664) );
  XNOR2_X1 U745 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U746 ( .A(n666), .B(G290), .ZN(n911) );
  XNOR2_X1 U747 ( .A(n667), .B(n911), .ZN(n668) );
  XNOR2_X1 U748 ( .A(KEYINPUT81), .B(n668), .ZN(n669) );
  NOR2_X1 U749 ( .A1(n670), .A2(n669), .ZN(n673) );
  NOR2_X1 U750 ( .A1(G868), .A2(n671), .ZN(n672) );
  NOR2_X1 U751 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2084), .A2(G2078), .ZN(n674) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U754 ( .A1(n675), .A2(G2090), .ZN(n676) );
  XNOR2_X1 U755 ( .A(n676), .B(KEYINPUT21), .ZN(n677) );
  XNOR2_X1 U756 ( .A(KEYINPUT82), .B(n677), .ZN(n678) );
  NAND2_X1 U757 ( .A1(G2072), .A2(n678), .ZN(G158) );
  XOR2_X1 U758 ( .A(KEYINPUT83), .B(G44), .Z(n679) );
  XNOR2_X1 U759 ( .A(KEYINPUT3), .B(n679), .ZN(G218) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U761 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U762 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U763 ( .A1(G96), .A2(n682), .ZN(n842) );
  NAND2_X1 U764 ( .A1(G2106), .A2(n842), .ZN(n683) );
  XNOR2_X1 U765 ( .A(n683), .B(KEYINPUT84), .ZN(n688) );
  NOR2_X1 U766 ( .A1(G236), .A2(G238), .ZN(n684) );
  NAND2_X1 U767 ( .A1(G69), .A2(n684), .ZN(n685) );
  NOR2_X1 U768 ( .A1(n685), .A2(G237), .ZN(n686) );
  XNOR2_X1 U769 ( .A(n686), .B(KEYINPUT85), .ZN(n843) );
  NAND2_X1 U770 ( .A1(G567), .A2(n843), .ZN(n687) );
  NAND2_X1 U771 ( .A1(n688), .A2(n687), .ZN(n916) );
  NAND2_X1 U772 ( .A1(G483), .A2(G661), .ZN(n689) );
  NOR2_X1 U773 ( .A1(n916), .A2(n689), .ZN(n841) );
  NAND2_X1 U774 ( .A1(n841), .A2(G36), .ZN(G176) );
  XNOR2_X1 U775 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  XOR2_X1 U776 ( .A(G1981), .B(G305), .Z(n984) );
  NAND2_X1 U777 ( .A1(G160), .A2(G40), .ZN(n786) );
  INV_X1 U778 ( .A(n786), .ZN(n692) );
  NOR2_X1 U779 ( .A1(n690), .A2(G1384), .ZN(n691) );
  NOR2_X1 U780 ( .A1(G2084), .A2(n748), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n693), .A2(G8), .ZN(n746) );
  NAND2_X1 U782 ( .A1(G8), .A2(n748), .ZN(n779) );
  NOR2_X1 U783 ( .A1(G1966), .A2(n779), .ZN(n744) );
  NOR2_X1 U784 ( .A1(n744), .A2(n693), .ZN(n694) );
  XNOR2_X1 U785 ( .A(n694), .B(KEYINPUT100), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n695), .A2(G8), .ZN(n696) );
  XNOR2_X1 U787 ( .A(n696), .B(KEYINPUT30), .ZN(n697) );
  NOR2_X1 U788 ( .A1(G168), .A2(n697), .ZN(n703) );
  INV_X2 U789 ( .A(n748), .ZN(n724) );
  NOR2_X1 U790 ( .A1(n724), .A2(G1961), .ZN(n698) );
  XOR2_X1 U791 ( .A(KEYINPUT96), .B(n698), .Z(n700) );
  XNOR2_X1 U792 ( .A(KEYINPUT25), .B(G2078), .ZN(n949) );
  NAND2_X1 U793 ( .A1(n724), .A2(n949), .ZN(n699) );
  NAND2_X1 U794 ( .A1(n700), .A2(n699), .ZN(n707) );
  NOR2_X1 U795 ( .A1(G171), .A2(n707), .ZN(n701) );
  XOR2_X1 U796 ( .A(KEYINPUT101), .B(n701), .Z(n702) );
  NOR2_X1 U797 ( .A1(n703), .A2(n702), .ZN(n706) );
  INV_X1 U798 ( .A(KEYINPUT102), .ZN(n704) );
  NAND2_X1 U799 ( .A1(n707), .A2(G171), .ZN(n740) );
  INV_X1 U800 ( .A(KEYINPUT29), .ZN(n738) );
  INV_X1 U801 ( .A(G299), .ZN(n714) );
  NAND2_X1 U802 ( .A1(n724), .A2(G2072), .ZN(n708) );
  XNOR2_X1 U803 ( .A(n708), .B(KEYINPUT27), .ZN(n710) );
  XNOR2_X1 U804 ( .A(G1956), .B(KEYINPUT97), .ZN(n993) );
  NOR2_X1 U805 ( .A1(n993), .A2(n724), .ZN(n709) );
  NOR2_X1 U806 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U807 ( .A(KEYINPUT98), .B(n711), .ZN(n713) );
  NOR2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n712) );
  XOR2_X1 U809 ( .A(n712), .B(KEYINPUT28), .Z(n736) );
  NAND2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n734) );
  NOR2_X1 U811 ( .A1(n724), .A2(n994), .ZN(n715) );
  NAND2_X1 U812 ( .A1(KEYINPUT26), .A2(n715), .ZN(n717) );
  NAND2_X1 U813 ( .A1(n717), .A2(KEYINPUT99), .ZN(n722) );
  INV_X1 U814 ( .A(KEYINPUT99), .ZN(n720) );
  NAND2_X1 U815 ( .A1(G1996), .A2(n724), .ZN(n716) );
  XNOR2_X1 U816 ( .A(KEYINPUT26), .B(n716), .ZN(n718) );
  NAND2_X1 U817 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U818 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U819 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U820 ( .A1(n975), .A2(n723), .ZN(n728) );
  NAND2_X1 U821 ( .A1(G1348), .A2(n748), .ZN(n726) );
  NAND2_X1 U822 ( .A1(G2067), .A2(n724), .ZN(n725) );
  NAND2_X1 U823 ( .A1(n726), .A2(n725), .ZN(n729) );
  NOR2_X1 U824 ( .A1(n730), .A2(n729), .ZN(n727) );
  OR2_X1 U825 ( .A1(n728), .A2(n727), .ZN(n732) );
  NAND2_X1 U826 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U827 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U828 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U829 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U830 ( .A(n738), .B(n737), .ZN(n739) );
  NAND2_X1 U831 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n747) );
  XNOR2_X1 U833 ( .A(n747), .B(KEYINPUT103), .ZN(n743) );
  NOR2_X1 U834 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U835 ( .A1(n746), .A2(n745), .ZN(n758) );
  NAND2_X1 U836 ( .A1(n747), .A2(G286), .ZN(n753) );
  NOR2_X1 U837 ( .A1(G1971), .A2(n779), .ZN(n750) );
  NOR2_X1 U838 ( .A1(G2090), .A2(n748), .ZN(n749) );
  NOR2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n751), .A2(G303), .ZN(n752) );
  NAND2_X1 U841 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U842 ( .A1(n754), .A2(G8), .ZN(n756) );
  XNOR2_X1 U843 ( .A(n756), .B(n755), .ZN(n757) );
  NAND2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n772) );
  NOR2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n765) );
  NOR2_X1 U846 ( .A1(G1971), .A2(G303), .ZN(n759) );
  NOR2_X1 U847 ( .A1(n765), .A2(n759), .ZN(n972) );
  INV_X1 U848 ( .A(KEYINPUT33), .ZN(n760) );
  AND2_X1 U849 ( .A1(n972), .A2(n760), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n772), .A2(n761), .ZN(n764) );
  NAND2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n973) );
  INV_X1 U852 ( .A(n973), .ZN(n762) );
  OR2_X1 U853 ( .A1(KEYINPUT33), .A2(n516), .ZN(n763) );
  NAND2_X1 U854 ( .A1(n764), .A2(n763), .ZN(n768) );
  NAND2_X1 U855 ( .A1(n765), .A2(KEYINPUT33), .ZN(n766) );
  NOR2_X1 U856 ( .A1(n766), .A2(n779), .ZN(n767) );
  NOR2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U858 ( .A1(n984), .A2(n769), .ZN(n783) );
  NOR2_X1 U859 ( .A1(G2090), .A2(G303), .ZN(n770) );
  NAND2_X1 U860 ( .A1(G8), .A2(n770), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n773), .A2(n779), .ZN(n774) );
  XNOR2_X1 U863 ( .A(n774), .B(KEYINPUT105), .ZN(n781) );
  NOR2_X1 U864 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XNOR2_X1 U865 ( .A(KEYINPUT24), .B(KEYINPUT95), .ZN(n775) );
  XNOR2_X1 U866 ( .A(n775), .B(KEYINPUT94), .ZN(n776) );
  XNOR2_X1 U867 ( .A(n777), .B(n776), .ZN(n778) );
  NOR2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n784), .B(KEYINPUT106), .ZN(n820) );
  NOR2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n816) );
  XOR2_X1 U873 ( .A(G2067), .B(KEYINPUT37), .Z(n821) );
  NAND2_X1 U874 ( .A1(G104), .A2(n515), .ZN(n788) );
  NAND2_X1 U875 ( .A1(G140), .A2(n609), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U877 ( .A(KEYINPUT34), .B(n789), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G116), .A2(n889), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G128), .A2(n890), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U881 ( .A(n792), .B(KEYINPUT35), .Z(n793) );
  NOR2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U883 ( .A(KEYINPUT36), .B(n795), .Z(n796) );
  XNOR2_X1 U884 ( .A(KEYINPUT92), .B(n796), .ZN(n887) );
  AND2_X1 U885 ( .A1(n821), .A2(n887), .ZN(n923) );
  NAND2_X1 U886 ( .A1(n816), .A2(n923), .ZN(n822) );
  XNOR2_X1 U887 ( .A(KEYINPUT90), .B(G1986), .ZN(n797) );
  XNOR2_X1 U888 ( .A(n797), .B(G290), .ZN(n988) );
  NAND2_X1 U889 ( .A1(n988), .A2(n816), .ZN(n798) );
  XOR2_X1 U890 ( .A(KEYINPUT91), .B(n798), .Z(n799) );
  AND2_X1 U891 ( .A1(n822), .A2(n799), .ZN(n818) );
  NAND2_X1 U892 ( .A1(G107), .A2(n889), .ZN(n801) );
  NAND2_X1 U893 ( .A1(G119), .A2(n890), .ZN(n800) );
  NAND2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U895 ( .A1(G95), .A2(n515), .ZN(n802) );
  XNOR2_X1 U896 ( .A(KEYINPUT93), .B(n802), .ZN(n803) );
  NOR2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U898 ( .A1(n609), .A2(G131), .ZN(n805) );
  NAND2_X1 U899 ( .A1(n806), .A2(n805), .ZN(n903) );
  AND2_X1 U900 ( .A1(n903), .A2(G1991), .ZN(n815) );
  NAND2_X1 U901 ( .A1(G117), .A2(n889), .ZN(n808) );
  NAND2_X1 U902 ( .A1(G129), .A2(n890), .ZN(n807) );
  NAND2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n515), .A2(G105), .ZN(n809) );
  XOR2_X1 U905 ( .A(KEYINPUT38), .B(n809), .Z(n810) );
  NOR2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n609), .A2(G141), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n902) );
  AND2_X1 U909 ( .A1(n902), .A2(G1996), .ZN(n814) );
  NOR2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n927) );
  INV_X1 U911 ( .A(n816), .ZN(n832) );
  NOR2_X1 U912 ( .A1(n927), .A2(n832), .ZN(n825) );
  INV_X1 U913 ( .A(n825), .ZN(n817) );
  AND2_X1 U914 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n835) );
  NOR2_X1 U916 ( .A1(n821), .A2(n887), .ZN(n922) );
  INV_X1 U917 ( .A(n822), .ZN(n829) );
  NOR2_X1 U918 ( .A1(G1996), .A2(n902), .ZN(n937) );
  NOR2_X1 U919 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U920 ( .A1(G1991), .A2(n903), .ZN(n929) );
  NOR2_X1 U921 ( .A1(n823), .A2(n929), .ZN(n824) );
  NOR2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U923 ( .A1(n937), .A2(n826), .ZN(n827) );
  XOR2_X1 U924 ( .A(KEYINPUT39), .B(n827), .Z(n828) );
  NOR2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U926 ( .A1(n922), .A2(n830), .ZN(n831) );
  NOR2_X1 U927 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U928 ( .A(n833), .B(KEYINPUT107), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n836), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n837), .ZN(G217) );
  INV_X1 U932 ( .A(n837), .ZN(G223) );
  NAND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n838) );
  XOR2_X1 U934 ( .A(KEYINPUT110), .B(n838), .Z(n839) );
  NAND2_X1 U935 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U937 ( .A1(n841), .A2(n840), .ZN(G188) );
  NOR2_X1 U938 ( .A1(n843), .A2(n842), .ZN(G325) );
  XNOR2_X1 U939 ( .A(KEYINPUT111), .B(G325), .ZN(G261) );
  INV_X1 U941 ( .A(G96), .ZN(G221) );
  XOR2_X1 U942 ( .A(G2678), .B(G2084), .Z(n845) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2090), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n849) );
  XNOR2_X1 U946 ( .A(G2078), .B(G2072), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U948 ( .A(G2096), .B(KEYINPUT113), .Z(n851) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U951 ( .A(n853), .B(n852), .Z(G227) );
  XOR2_X1 U952 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n855) );
  XNOR2_X1 U953 ( .A(KEYINPUT115), .B(G2474), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U955 ( .A(n856), .B(KEYINPUT41), .Z(n858) );
  XNOR2_X1 U956 ( .A(G1991), .B(G1996), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n866) );
  XOR2_X1 U958 ( .A(G1986), .B(G1961), .Z(n860) );
  XNOR2_X1 U959 ( .A(G1976), .B(G1971), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U961 ( .A(KEYINPUT114), .B(G1956), .Z(n862) );
  XNOR2_X1 U962 ( .A(G1981), .B(G1966), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U964 ( .A(n864), .B(n863), .Z(n865) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G124), .A2(n890), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U968 ( .A1(n889), .A2(G112), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G100), .A2(n515), .ZN(n871) );
  NAND2_X1 U971 ( .A1(G136), .A2(n609), .ZN(n870) );
  NAND2_X1 U972 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U973 ( .A1(n873), .A2(n872), .ZN(G162) );
  XOR2_X1 U974 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n875) );
  XNOR2_X1 U975 ( .A(n925), .B(KEYINPUT46), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U977 ( .A(n876), .B(KEYINPUT121), .Z(n885) );
  NAND2_X1 U978 ( .A1(G103), .A2(n515), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G139), .A2(n609), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n883) );
  NAND2_X1 U981 ( .A1(G115), .A2(n889), .ZN(n880) );
  NAND2_X1 U982 ( .A1(G127), .A2(n890), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n932) );
  XNOR2_X1 U986 ( .A(n932), .B(KEYINPUT48), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U988 ( .A(n886), .B(G164), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n888), .B(n887), .ZN(n909) );
  NAND2_X1 U990 ( .A1(G118), .A2(n889), .ZN(n892) );
  NAND2_X1 U991 ( .A1(G130), .A2(n890), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U993 ( .A(KEYINPUT118), .B(n893), .ZN(n901) );
  XNOR2_X1 U994 ( .A(KEYINPUT45), .B(KEYINPUT120), .ZN(n899) );
  NAND2_X1 U995 ( .A1(n609), .A2(G142), .ZN(n897) );
  NAND2_X1 U996 ( .A1(n515), .A2(G106), .ZN(n895) );
  XOR2_X1 U997 ( .A(KEYINPUT119), .B(n895), .Z(n896) );
  NAND2_X1 U998 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U999 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U1000 ( .A1(n901), .A2(n900), .ZN(n907) );
  XOR2_X1 U1001 ( .A(G162), .B(G160), .Z(n905) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G395) );
  XOR2_X1 U1007 ( .A(n970), .B(n911), .Z(n913) );
  XOR2_X1 U1008 ( .A(G286), .B(G301), .Z(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n914), .B(n975), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n915), .ZN(G397) );
  XOR2_X1 U1012 ( .A(KEYINPUT112), .B(n916), .Z(G319) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n918), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n919) );
  AND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n921), .A2(G319), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n931) );
  XOR2_X1 U1022 ( .A(G2084), .B(G160), .Z(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n942) );
  XOR2_X1 U1027 ( .A(G2072), .B(n932), .Z(n934) );
  XOR2_X1 U1028 ( .A(G164), .B(G2078), .Z(n933) );
  NOR2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(KEYINPUT50), .B(n935), .ZN(n940) );
  XOR2_X1 U1031 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1033 ( .A(KEYINPUT51), .B(n938), .Z(n939) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(KEYINPUT52), .B(n943), .ZN(n944) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n964) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n964), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n945), .A2(G29), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(KEYINPUT124), .B(n946), .ZN(n1022) );
  XOR2_X1 U1041 ( .A(G29), .B(KEYINPUT126), .Z(n967) );
  XNOR2_X1 U1042 ( .A(KEYINPUT125), .B(G2072), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(n947), .B(G33), .ZN(n957) );
  XOR2_X1 U1044 ( .A(G32), .B(G1996), .Z(n948) );
  NAND2_X1 U1045 ( .A1(n948), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1046 ( .A(G27), .B(n949), .ZN(n953) );
  XNOR2_X1 U1047 ( .A(G1991), .B(G25), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(G26), .B(G2067), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(n958), .B(KEYINPUT53), .ZN(n961) );
  XOR2_X1 U1054 ( .A(G2084), .B(G34), .Z(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n959), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G35), .B(G2090), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n965) );
  XOR2_X1 U1059 ( .A(n965), .B(n964), .Z(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(G11), .A2(n968), .ZN(n1020) );
  XNOR2_X1 U1062 ( .A(KEYINPUT56), .B(KEYINPUT127), .ZN(n969) );
  XOR2_X1 U1063 ( .A(G16), .B(n969), .Z(n992) );
  XNOR2_X1 U1064 ( .A(G1348), .B(n970), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n983) );
  XOR2_X1 U1066 ( .A(G301), .B(G1961), .Z(n981) );
  XOR2_X1 U1067 ( .A(G1956), .B(G299), .Z(n974) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n979) );
  XOR2_X1 U1069 ( .A(G1341), .B(n975), .Z(n977) );
  NAND2_X1 U1070 ( .A1(G1971), .A2(G303), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n990) );
  XNOR2_X1 U1075 ( .A(G168), .B(G1966), .ZN(n985) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1077 ( .A(KEYINPUT57), .B(n986), .Z(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n1018) );
  INV_X1 U1081 ( .A(G16), .ZN(n1016) );
  XNOR2_X1 U1082 ( .A(G20), .B(n993), .ZN(n998) );
  XNOR2_X1 U1083 ( .A(G1981), .B(G6), .ZN(n996) );
  XOR2_X1 U1084 ( .A(n994), .B(G19), .Z(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n1001) );
  XOR2_X1 U1087 ( .A(KEYINPUT59), .B(G1348), .Z(n999) );
  XNOR2_X1 U1088 ( .A(G4), .B(n999), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(KEYINPUT60), .B(n1002), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(G1966), .B(G21), .ZN(n1004) );
  XNOR2_X1 U1092 ( .A(G5), .B(G1961), .ZN(n1003) );
  NOR2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1013) );
  XNOR2_X1 U1095 ( .A(G1976), .B(G23), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1010) );
  XOR2_X1 U1098 ( .A(G1986), .B(G24), .Z(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(KEYINPUT58), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1023), .ZN(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

