//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT0), .Z(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G50), .ZN(new_n209));
  INV_X1    g0009(.A(G226), .ZN(new_n210));
  INV_X1    g0010(.A(G116), .ZN(new_n211));
  INV_X1    g0011(.A(G270), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G58), .B2(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G68), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G244), .ZN(new_n217));
  XOR2_X1   g0017(.A(KEYINPUT65), .B(G77), .Z(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n204), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(new_n215), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n207), .B(new_n225), .C1(new_n228), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G264), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n212), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT66), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT67), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n246), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT13), .ZN(new_n252));
  INV_X1    g0052(.A(G274), .ZN(new_n253));
  XOR2_X1   g0053(.A(KEYINPUT69), .B(G45), .Z(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  AOI211_X1 g0055(.A(G1), .B(new_n253), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  OAI211_X1 g0057(.A(G1), .B(G13), .C1(new_n257), .C2(new_n255), .ZN(new_n258));
  INV_X1    g0058(.A(G232), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G1698), .ZN(new_n260));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  OAI221_X1 g0062(.A(new_n260), .B1(G226), .B2(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G97), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n258), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n258), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n269), .A2(new_n216), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n252), .B1(new_n266), .B2(new_n271), .ZN(new_n272));
  NOR4_X1   g0072(.A1(new_n256), .A2(new_n265), .A3(KEYINPUT13), .A4(new_n270), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G190), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n215), .A2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(G13), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n276), .A2(G1), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n278), .B(KEYINPUT12), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n226), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(new_n267), .B2(G20), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n279), .B1(G68), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G77), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n227), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT70), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(new_n227), .A3(new_n257), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n288));
  AND2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI221_X1 g0089(.A(new_n276), .B1(new_n284), .B2(new_n285), .C1(new_n289), .C2(new_n209), .ZN(new_n290));
  XOR2_X1   g0090(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n281), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n281), .ZN(new_n293));
  INV_X1    g0093(.A(new_n291), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n275), .A2(new_n283), .A3(new_n292), .A4(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G200), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n274), .A2(new_n297), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n266), .A2(new_n271), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT13), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n266), .A2(new_n252), .A3(new_n271), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT76), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT14), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n274), .A2(G179), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n304), .B(G169), .C1(new_n272), .C2(new_n273), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT14), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n295), .A2(new_n283), .A3(new_n292), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n299), .A2(new_n312), .A3(KEYINPUT77), .ZN(new_n313));
  OAI21_X1  g0113(.A(G20), .B1(new_n230), .B2(G50), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT8), .B(G58), .ZN(new_n315));
  INV_X1    g0115(.A(G150), .ZN(new_n316));
  OAI221_X1 g0116(.A(new_n314), .B1(new_n285), .B2(new_n315), .C1(new_n289), .C2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n267), .A2(G13), .A3(G20), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n317), .A2(new_n281), .B1(new_n209), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n282), .A2(G50), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n257), .ZN(new_n324));
  NAND2_X1  g0124(.A1(KEYINPUT3), .A2(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G1698), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G222), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G223), .A2(G1698), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n330), .B(new_n331), .C1(new_n218), .C2(new_n326), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n254), .A2(new_n255), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(new_n267), .A3(G274), .ZN(new_n334));
  INV_X1    g0134(.A(new_n269), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(G226), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n332), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G169), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n322), .B(new_n339), .C1(G179), .C2(new_n337), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT72), .B(G200), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT9), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n342), .B(new_n344), .C1(new_n322), .C2(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT9), .B1(new_n320), .B2(new_n321), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT10), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n346), .A2(KEYINPUT10), .A3(new_n347), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n340), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G238), .A2(G1698), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n326), .B(new_n353), .C1(new_n259), .C2(G1698), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n354), .B(new_n331), .C1(G107), .C2(new_n326), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n335), .A2(G244), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n334), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n343), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n282), .A2(G77), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  OR3_X1    g0160(.A1(new_n360), .A2(KEYINPUT71), .A3(new_n285), .ZN(new_n361));
  INV_X1    g0161(.A(new_n315), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n287), .A2(new_n288), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n218), .A2(G20), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT71), .B1(new_n360), .B2(new_n285), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n361), .A2(new_n364), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n281), .B1(new_n219), .B2(new_n319), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n358), .A2(new_n359), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT73), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n357), .A2(new_n341), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT73), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n358), .A2(new_n372), .A3(new_n368), .A4(new_n359), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n368), .A2(new_n359), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n357), .A2(new_n338), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n375), .B(new_n376), .C1(G179), .C2(new_n357), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT74), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n374), .A2(KEYINPUT74), .A3(new_n377), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n352), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n299), .A2(new_n312), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT77), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n261), .A2(new_n262), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT7), .B1(new_n386), .B2(new_n227), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n324), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n325), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n363), .A2(G159), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n227), .B1(new_n230), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n390), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n324), .A2(new_n227), .A3(new_n325), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n388), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n393), .B1(new_n401), .B2(G68), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(KEYINPUT16), .A3(new_n391), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n397), .A2(new_n281), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n210), .A2(G1698), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n405), .B1(G223), .B2(G1698), .C1(new_n261), .C2(new_n262), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G87), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n258), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n256), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n269), .A2(new_n259), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G200), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n256), .A2(new_n408), .A3(new_n410), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G190), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n267), .A2(G20), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n362), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT78), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n319), .A2(new_n281), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n418), .A2(new_n419), .B1(new_n319), .B2(new_n315), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n404), .A2(new_n413), .A3(new_n415), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n412), .A2(G169), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n414), .A2(G179), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n404), .A2(KEYINPUT79), .A3(new_n420), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT79), .B1(new_n404), .B2(new_n420), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT79), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT16), .B1(new_n402), .B2(new_n391), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n215), .B1(new_n400), .B2(new_n388), .ZN(new_n434));
  INV_X1    g0234(.A(new_n391), .ZN(new_n435));
  NOR4_X1   g0235(.A1(new_n434), .A2(new_n435), .A3(new_n396), .A4(new_n393), .ZN(new_n436));
  INV_X1    g0236(.A(new_n281), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n420), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n432), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n404), .A2(KEYINPUT79), .A3(new_n420), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n442), .A2(KEYINPUT18), .A3(new_n426), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n423), .B1(new_n431), .B2(new_n443), .ZN(new_n444));
  AND4_X1   g0244(.A1(new_n313), .A2(new_n382), .A3(new_n385), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G264), .A2(G1698), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n326), .B(new_n447), .C1(new_n222), .C2(G1698), .ZN(new_n448));
  INV_X1    g0248(.A(G303), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n258), .B1(new_n386), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(KEYINPUT5), .A2(G41), .ZN(new_n452));
  NOR2_X1   g0252(.A1(KEYINPUT5), .A2(G41), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n267), .A2(G45), .ZN(new_n455));
  OAI211_X1 g0255(.A(G270), .B(new_n258), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n267), .A2(G45), .A3(G274), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n454), .A2(KEYINPUT81), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT81), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT5), .B(G41), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n267), .A2(G45), .A3(G274), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n456), .B(KEYINPUT89), .C1(new_n458), .C2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT81), .B1(new_n454), .B2(new_n457), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n460), .A2(new_n459), .A3(new_n461), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT89), .B1(new_n467), .B2(new_n456), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n451), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G200), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n437), .B(new_n318), .C1(G1), .C2(new_n257), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G116), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n267), .A2(new_n211), .A3(G13), .A4(G20), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n474), .B(KEYINPUT90), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT91), .ZN(new_n477));
  AOI21_X1  g0277(.A(G20), .B1(G33), .B2(G283), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n257), .A2(G97), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n479), .A3(new_n477), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n280), .A2(new_n226), .B1(G20), .B2(new_n211), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT20), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n482), .ZN(new_n486));
  OAI211_X1 g0286(.A(KEYINPUT20), .B(new_n484), .C1(new_n486), .C2(new_n480), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n473), .B(new_n476), .C1(new_n485), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n470), .B(new_n490), .C1(new_n341), .C2(new_n469), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n456), .B1(new_n458), .B2(new_n462), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT89), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n494), .A2(new_n463), .B1(new_n448), .B2(new_n450), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(G179), .A3(new_n489), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT21), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n463), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n338), .B1(new_n498), .B2(new_n451), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n497), .B1(new_n499), .B2(new_n489), .ZN(new_n500));
  AND4_X1   g0300(.A1(new_n497), .A2(new_n469), .A3(G169), .A4(new_n489), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n491), .B(new_n496), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(G244), .B1(new_n261), .B2(new_n262), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n504), .A2(G1698), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n507), .B(G244), .C1(new_n262), .C2(new_n261), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(G250), .B1(new_n261), .B2(new_n262), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n327), .B1(new_n510), .B2(KEYINPUT4), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n331), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(G179), .ZN(new_n513));
  INV_X1    g0313(.A(new_n455), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n331), .B1(new_n460), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n515), .A2(G257), .B1(new_n465), .B2(new_n466), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(G257), .B(new_n258), .C1(new_n454), .C2(new_n455), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n467), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n503), .A2(new_n504), .B1(G33), .B2(G283), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n504), .B1(new_n326), .B2(G250), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n520), .B(new_n508), .C1(new_n327), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n519), .B1(new_n331), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n517), .B(KEYINPUT84), .C1(new_n523), .C2(G169), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT84), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n525), .A3(new_n513), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n471), .A2(new_n221), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n401), .A2(G107), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n363), .A2(G77), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT6), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT80), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT80), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT6), .ZN(new_n534));
  INV_X1    g0334(.A(G107), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n532), .A2(new_n534), .A3(G97), .A4(new_n535), .ZN(new_n536));
  XOR2_X1   g0336(.A(G97), .B(G107), .Z(new_n537));
  XNOR2_X1  g0337(.A(KEYINPUT80), .B(KEYINPUT6), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G20), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n529), .A2(new_n530), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n528), .B1(new_n541), .B2(new_n281), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n319), .A2(new_n221), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n542), .A2(KEYINPUT83), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT83), .B1(new_n542), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n527), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n227), .A2(G107), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n547), .B(KEYINPUT23), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n227), .A2(G33), .A3(G116), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT22), .ZN(new_n550));
  AOI21_X1  g0350(.A(G20), .B1(new_n324), .B2(new_n325), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(G87), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n227), .B(G87), .C1(new_n261), .C2(new_n262), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(KEYINPUT22), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n548), .B(new_n549), .C1(new_n552), .C2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n551), .A2(new_n550), .A3(G87), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n553), .A2(KEYINPUT22), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(KEYINPUT24), .A3(new_n548), .A4(new_n549), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n557), .A2(new_n281), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n472), .A2(G107), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n319), .B(new_n535), .C1(KEYINPUT92), .C2(KEYINPUT25), .ZN(new_n564));
  NAND2_X1  g0364(.A1(KEYINPUT92), .A2(KEYINPUT25), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n562), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G250), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n327), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n222), .A2(G1698), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n569), .B(new_n570), .C1(new_n261), .C2(new_n262), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G294), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n331), .ZN(new_n574));
  OAI211_X1 g0374(.A(G264), .B(new_n258), .C1(new_n454), .C2(new_n455), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n467), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G169), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT93), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n574), .A2(new_n575), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(G179), .A3(new_n467), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT93), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n576), .A2(new_n581), .A3(G169), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n578), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n567), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n576), .A2(new_n297), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(G190), .B2(new_n576), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n586), .A2(new_n562), .A3(new_n563), .A4(new_n566), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT82), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G200), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n523), .A2(new_n341), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n512), .A2(new_n516), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n588), .B2(new_n297), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n543), .A3(new_n542), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n546), .A2(new_n584), .A3(new_n587), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n216), .A2(new_n327), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n217), .A2(G1698), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n596), .B(new_n597), .C1(new_n261), .C2(new_n262), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G33), .A2(G116), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n258), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n258), .A2(G250), .A3(new_n455), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT85), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n457), .B(new_n603), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n600), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT87), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n605), .A2(new_n606), .A3(G190), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n606), .B1(new_n605), .B2(G190), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT88), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(G190), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT87), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT88), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n607), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n551), .A2(G68), .ZN(new_n615));
  OR3_X1    g0415(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n264), .A2(new_n227), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(KEYINPUT19), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n264), .A2(G20), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n615), .B(new_n618), .C1(KEYINPUT19), .C2(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n620), .A2(new_n281), .B1(new_n319), .B2(new_n360), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n472), .A2(G87), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n343), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n605), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n610), .A2(new_n614), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n605), .A2(G179), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n338), .B2(new_n605), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT86), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n621), .B1(new_n360), .B2(new_n471), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT86), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n628), .B(new_n632), .C1(new_n338), .C2(new_n605), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n627), .A2(new_n634), .ZN(new_n635));
  NOR4_X1   g0435(.A1(new_n446), .A2(new_n502), .A3(new_n595), .A4(new_n635), .ZN(G372));
  NOR2_X1   g0436(.A1(new_n296), .A2(new_n298), .ZN(new_n637));
  AOI211_X1 g0437(.A(new_n637), .B(new_n423), .C1(new_n312), .C2(new_n377), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n426), .B1(new_n438), .B2(new_n439), .ZN(new_n639));
  XNOR2_X1  g0439(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI22_X1  g0442(.A1(new_n638), .A2(new_n642), .B1(new_n350), .B2(new_n351), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n643), .A2(new_n340), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n629), .A2(new_n631), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n584), .B(new_n496), .C1(new_n500), .C2(new_n501), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n612), .A2(new_n607), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n626), .A2(new_n647), .B1(new_n631), .B2(new_n629), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n546), .A2(new_n587), .A3(new_n594), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n645), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT26), .B1(new_n635), .B2(new_n546), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n542), .A2(new_n543), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n648), .A2(new_n654), .A3(new_n655), .A4(new_n527), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n644), .B1(new_n446), .B2(new_n660), .ZN(G369));
  OAI21_X1  g0461(.A(new_n496), .B1(new_n500), .B2(new_n501), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n267), .A2(new_n227), .A3(G13), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n490), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n662), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n671), .B1(new_n502), .B2(new_n670), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n672), .A2(G330), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n584), .A2(new_n587), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n567), .A2(new_n668), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n674), .A2(new_n675), .B1(new_n584), .B2(new_n669), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  AND4_X1   g0477(.A1(new_n662), .A2(new_n584), .A3(new_n587), .A4(new_n669), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n584), .A2(new_n668), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(G399));
  NOR2_X1   g0481(.A1(new_n616), .A2(G116), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n205), .A2(new_n255), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(G1), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n231), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  AOI211_X1 g0486(.A(KEYINPUT29), .B(new_n668), .C1(new_n652), .C2(new_n658), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n546), .A2(new_n587), .A3(new_n594), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n689), .A2(new_n646), .A3(new_n648), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n648), .A2(new_n655), .A3(new_n527), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(KEYINPUT26), .ZN(new_n692));
  INV_X1    g0492(.A(new_n635), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT83), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n655), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n542), .A2(KEYINPUT83), .A3(new_n543), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n695), .A2(new_n696), .B1(new_n524), .B2(new_n526), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n693), .A2(new_n654), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n690), .A2(new_n645), .A3(new_n692), .A4(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n688), .B1(new_n699), .B2(new_n669), .ZN(new_n700));
  INV_X1    g0500(.A(G330), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n655), .B1(new_n592), .B2(new_n590), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n697), .A2(new_n674), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n502), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n693), .A3(new_n704), .A4(new_n669), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n495), .A2(new_n579), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n523), .A2(G179), .A3(new_n605), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n591), .A2(new_n628), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(KEYINPUT30), .A3(new_n495), .A4(new_n579), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n605), .B1(new_n579), .B2(new_n467), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n712), .A2(new_n469), .A3(new_n513), .A4(new_n591), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n668), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT31), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n717), .A3(new_n668), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n701), .B1(new_n705), .B2(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n687), .A2(new_n700), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n686), .B1(new_n721), .B2(G1), .ZN(G364));
  NAND2_X1  g0522(.A1(new_n250), .A2(G45), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n232), .A2(new_n254), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n386), .A2(new_n205), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT95), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(G355), .A2(new_n205), .A3(new_n326), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n727), .B(new_n728), .C1(G116), .C2(new_n205), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G13), .A2(G33), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT96), .Z(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n226), .B1(G20), .B2(new_n338), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n729), .A2(new_n735), .ZN(new_n736));
  AND3_X1   g0536(.A1(KEYINPUT97), .A2(G20), .A3(G179), .ZN(new_n737));
  AOI21_X1  g0537(.A(KEYINPUT97), .B1(G20), .B2(G179), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G190), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n227), .A2(G179), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(new_n741), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n743), .A2(G311), .B1(G329), .B2(new_n746), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n739), .A2(new_n341), .A3(new_n297), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G326), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n343), .A2(new_n744), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n341), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G303), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n747), .A2(new_n386), .A3(new_n749), .A4(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT98), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(new_n750), .B2(G190), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n343), .A2(KEYINPUT98), .A3(new_n341), .A4(new_n744), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n753), .B1(G283), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G294), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n341), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n513), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G20), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G322), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n740), .A2(new_n761), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n759), .B1(new_n760), .B2(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n739), .A2(G190), .A3(new_n297), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT33), .B(G317), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n746), .A2(G159), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT32), .ZN(new_n772));
  INV_X1    g0572(.A(new_n768), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n326), .B1(new_n773), .B2(new_n215), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(G97), .B2(new_n763), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n751), .A2(G87), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n743), .A2(new_n218), .B1(new_n748), .B2(G50), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n758), .A2(G107), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n766), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n772), .B(new_n779), .C1(G58), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n770), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT99), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n736), .B1(new_n783), .B2(new_n734), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n277), .A2(G20), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G45), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n683), .A2(G1), .A3(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n733), .B(KEYINPUT100), .Z(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI211_X1 g0590(.A(new_n784), .B(new_n788), .C1(new_n672), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n673), .A2(new_n788), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G330), .B2(new_n672), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  INV_X1    g0595(.A(new_n374), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n375), .A2(new_n668), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT102), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n377), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n377), .A2(new_n668), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n660), .B2(new_n668), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT102), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n797), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n374), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n800), .B1(new_n806), .B2(new_n377), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n669), .B(new_n807), .C1(new_n651), .C2(new_n657), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(new_n720), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n787), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n758), .A2(G87), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n812), .B1(new_n211), .B2(new_n742), .C1(new_n760), .C2(new_n766), .ZN(new_n813));
  INV_X1    g0613(.A(new_n751), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n814), .A2(new_n535), .B1(new_n764), .B2(new_n221), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n386), .B1(new_n773), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n813), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n748), .ZN(new_n819));
  INV_X1    g0619(.A(G311), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n818), .B1(new_n449), .B2(new_n819), .C1(new_n820), .C2(new_n745), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G143), .A2(new_n780), .B1(new_n743), .B2(G159), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n748), .A2(G137), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n768), .A2(G150), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT101), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(KEYINPUT101), .B1(new_n823), .B2(new_n824), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n822), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT34), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n745), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n757), .A2(new_n215), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(G50), .C2(new_n751), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n829), .A2(new_n326), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n764), .A2(new_n229), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n821), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n734), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n802), .A2(new_n731), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n734), .A2(new_n730), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n284), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n837), .A2(new_n838), .A3(new_n788), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n811), .A2(new_n841), .ZN(G384));
  AOI21_X1  g0642(.A(new_n211), .B1(new_n539), .B2(KEYINPUT35), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n843), .B(new_n228), .C1(KEYINPUT35), .C2(new_n539), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT36), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n232), .A2(new_n218), .A3(new_n392), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(G50), .B2(new_n215), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(G1), .A3(new_n277), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT103), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT40), .ZN(new_n851));
  XNOR2_X1  g0651(.A(new_n421), .B(KEYINPUT17), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT18), .B1(new_n442), .B2(new_n426), .ZN(new_n853));
  INV_X1    g0653(.A(new_n426), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n430), .B(new_n854), .C1(new_n440), .C2(new_n441), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n852), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n666), .B1(new_n404), .B2(new_n420), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n666), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n427), .B2(new_n428), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n421), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n429), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n639), .A2(new_n421), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n864), .B2(new_n857), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT38), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n857), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT38), .B(new_n866), .C1(new_n444), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NOR4_X1   g0671(.A1(new_n595), .A2(new_n502), .A3(new_n635), .A4(new_n668), .ZN(new_n872));
  INV_X1    g0672(.A(new_n718), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n717), .B1(new_n714), .B2(new_n668), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT107), .B1(new_n872), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n310), .A2(new_n311), .A3(new_n668), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n311), .A2(new_n668), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n299), .A2(new_n312), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n802), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT107), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n705), .A2(new_n881), .A3(new_n719), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n876), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n851), .B1(new_n871), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n876), .A2(new_n882), .ZN(new_n885));
  XNOR2_X1  g0685(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n860), .A2(new_n421), .A3(new_n639), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n442), .B1(new_n426), .B2(new_n859), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n887), .A2(KEYINPUT37), .B1(new_n888), .B2(new_n862), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n860), .B1(new_n641), .B2(new_n852), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n851), .B1(new_n891), .B2(new_n869), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n892), .A2(new_n880), .A3(new_n876), .A4(new_n882), .ZN(new_n893));
  AND4_X1   g0693(.A1(new_n445), .A2(new_n884), .A3(new_n885), .A4(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n884), .A2(G330), .A3(new_n893), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n445), .A2(G330), .A3(new_n876), .A4(new_n882), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n866), .B1(new_n444), .B2(new_n868), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n869), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n879), .A2(new_n877), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT105), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n800), .B(KEYINPUT104), .Z(new_n904));
  AND3_X1   g0704(.A1(new_n808), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n903), .B1(new_n808), .B2(new_n904), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n901), .B(new_n902), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n642), .A2(new_n666), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n891), .A2(new_n869), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n900), .A2(KEYINPUT39), .A3(new_n869), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n312), .A2(new_n668), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AND3_X1   g0714(.A1(new_n907), .A2(new_n908), .A3(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n897), .B(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n445), .B1(new_n687), .B2(new_n700), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n644), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n785), .A2(new_n267), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n850), .B1(new_n919), .B2(new_n920), .ZN(G367));
  NAND2_X1  g0721(.A1(new_n655), .A2(new_n668), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n922), .B1(new_n524), .B2(new_n526), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT108), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n546), .A2(new_n594), .A3(new_n922), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n926), .A2(new_n924), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n925), .B1(new_n927), .B2(new_n923), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n678), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT42), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(new_n567), .A3(new_n583), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n668), .B1(new_n931), .B2(new_n546), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT43), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n623), .A2(new_n668), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n648), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g0736(.A1(new_n645), .A2(new_n935), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n933), .A2(new_n934), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n934), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n941), .B(new_n942), .C1(new_n930), .C2(new_n932), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n928), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n944), .B1(new_n677), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n721), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n928), .A2(KEYINPUT44), .A3(new_n680), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT44), .B1(new_n928), .B2(new_n680), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n928), .A2(KEYINPUT45), .A3(new_n680), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT45), .B1(new_n928), .B2(new_n680), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n948), .B(new_n949), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n677), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n676), .B1(new_n662), .B2(new_n669), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n955), .A2(new_n678), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n673), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n947), .B1(new_n953), .B2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n683), .B(KEYINPUT41), .Z(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OAI211_X1 g0761(.A(G1), .B(new_n786), .C1(new_n959), .C2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n677), .A2(new_n945), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n940), .A2(new_n963), .A3(new_n943), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n946), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT110), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n780), .A2(G150), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n763), .A2(G68), .ZN(new_n969));
  INV_X1    g0769(.A(G137), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n970), .B2(new_n745), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n386), .B1(new_n748), .B2(G143), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n229), .B2(new_n814), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n971), .B(new_n973), .C1(new_n218), .C2(new_n758), .ZN(new_n974));
  INV_X1    g0774(.A(G159), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(new_n773), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n968), .B(new_n976), .C1(G50), .C2(new_n743), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n757), .A2(new_n221), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(G283), .B2(new_n743), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n979), .B(new_n386), .C1(new_n760), .C2(new_n773), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n819), .A2(new_n820), .B1(new_n766), .B2(new_n449), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT109), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n982), .A2(KEYINPUT109), .ZN(new_n985));
  INV_X1    g0785(.A(G317), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n984), .A2(new_n985), .B1(new_n986), .B2(new_n745), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n980), .B(new_n987), .C1(G107), .C2(new_n763), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n751), .A2(G116), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT46), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n977), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT47), .Z(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n734), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n939), .A2(new_n789), .ZN(new_n994));
  INV_X1    g0794(.A(new_n726), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n735), .B1(new_n205), .B2(new_n360), .C1(new_n236), .C2(new_n995), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n993), .A2(new_n788), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  AND3_X1   g0797(.A1(new_n965), .A2(new_n966), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n966), .B1(new_n965), .B2(new_n997), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(new_n999), .ZN(G387));
  NAND2_X1  g0800(.A1(new_n786), .A2(G1), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n958), .A2(new_n1001), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT111), .Z(new_n1003));
  NOR2_X1   g0803(.A1(new_n764), .A2(new_n360), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n751), .A2(new_n218), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1005), .B(new_n326), .C1(new_n215), .C2(new_n742), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(G150), .C2(new_n746), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT112), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(new_n748), .B2(G159), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1009), .B(new_n978), .C1(new_n362), .C2(new_n768), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n748), .A2(new_n1008), .A3(G159), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n780), .A2(G50), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n780), .A2(G317), .B1(new_n768), .B2(G311), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n449), .B2(new_n742), .C1(new_n765), .C2(new_n819), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT48), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n816), .B2(new_n764), .C1(new_n760), .C2(new_n814), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT49), .Z(new_n1018));
  AOI21_X1  g0818(.A(new_n326), .B1(new_n746), .B2(G326), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n757), .B2(new_n211), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1013), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n734), .ZN(new_n1022));
  OR3_X1    g0822(.A1(new_n315), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1023));
  OAI21_X1  g0823(.A(KEYINPUT50), .B1(new_n315), .B2(G50), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n682), .A3(new_n1024), .ZN(new_n1025));
  AOI211_X1 g0825(.A(G45), .B(new_n1025), .C1(G68), .C2(G77), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n726), .B1(new_n241), .B2(new_n254), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n326), .B(new_n205), .C1(new_n616), .C2(G116), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n205), .A2(G107), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n735), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n676), .A2(new_n790), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1022), .A2(new_n788), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n721), .A2(new_n958), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n721), .A2(new_n958), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n683), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1003), .B(new_n1033), .C1(new_n1034), .C2(new_n1037), .ZN(G393));
  OR2_X1    g0838(.A1(new_n953), .A2(new_n954), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n953), .A2(new_n954), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n1035), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n953), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1036), .C1(new_n1035), .C2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1039), .A2(new_n1001), .A3(new_n1040), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n787), .B1(new_n945), .B2(new_n733), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n726), .A2(new_n245), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n735), .B(new_n1047), .C1(new_n221), .C2(new_n205), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n743), .A2(G294), .B1(G283), .B2(new_n751), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n778), .B(new_n1049), .C1(new_n765), .C2(new_n745), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n819), .A2(new_n986), .B1(new_n766), .B2(new_n820), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT52), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n386), .B1(new_n211), .B2(new_n764), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1050), .B(new_n1057), .C1(G303), .C2(new_n768), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n764), .A2(new_n284), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n386), .B1(new_n768), .B2(G50), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n743), .A2(new_n362), .B1(G143), .B2(new_n746), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n812), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n819), .A2(new_n316), .B1(new_n766), .B2(new_n975), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT51), .Z(new_n1065));
  AOI211_X1 g0865(.A(new_n1063), .B(new_n1065), .C1(G68), .C2(new_n751), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1058), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT113), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n734), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1046), .B(new_n1048), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n1045), .A2(KEYINPUT114), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(KEYINPUT114), .B1(new_n1045), .B2(new_n1070), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1044), .B1(new_n1071), .B2(new_n1072), .ZN(G390));
  NAND4_X1  g0873(.A1(new_n876), .A2(new_n880), .A3(G330), .A4(new_n882), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n913), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1076), .A2(new_n1077), .B1(new_n911), .B2(new_n912), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n698), .A2(new_n692), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n668), .B1(new_n1079), .B2(new_n652), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n800), .B1(new_n1080), .B2(new_n799), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT115), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n902), .B(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n909), .B(new_n1077), .C1(new_n1081), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1075), .B1(new_n1078), .B2(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n720), .A2(new_n807), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n902), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n808), .A2(new_n904), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(KEYINPUT105), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n808), .A2(new_n903), .A3(new_n904), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n913), .B1(new_n1092), .B2(new_n902), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n911), .A2(new_n912), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1084), .B(new_n1088), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1086), .A2(new_n1095), .A3(new_n1001), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1094), .A2(new_n732), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n839), .A2(new_n315), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n768), .A2(G107), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n1100), .B(new_n832), .C1(G97), .C2(new_n743), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n386), .B1(new_n760), .B2(new_n745), .C1(new_n819), .C2(new_n816), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G87), .B2(new_n751), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n780), .A2(G116), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1101), .A2(new_n1060), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT54), .B(G143), .Z(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n773), .A2(new_n970), .B1(new_n742), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT116), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1108), .A2(new_n1109), .B1(new_n975), .B2(new_n764), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n1109), .B2(new_n1108), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n751), .A2(G150), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT53), .Z(new_n1113));
  INV_X1    g0913(.A(G128), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n819), .A2(new_n1114), .B1(new_n766), .B2(new_n830), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT118), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n326), .B1(new_n757), .B2(new_n209), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1117), .A2(KEYINPUT117), .B1(G125), .B2(new_n746), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1111), .A2(new_n1113), .A3(new_n1116), .A4(new_n1118), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1117), .A2(KEYINPUT117), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1105), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n734), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1097), .A2(new_n788), .A3(new_n1098), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1096), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n917), .A2(new_n896), .A3(new_n644), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1074), .B1(new_n1087), .B2(new_n902), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1092), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n876), .A2(G330), .A3(new_n807), .A4(new_n882), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1083), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n1088), .A3(new_n1081), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1125), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1086), .A2(new_n1095), .A3(new_n1131), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1132), .A2(new_n1036), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1086), .A2(new_n1095), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1125), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1124), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(G378));
  XOR2_X1   g0940(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1141));
  XNOR2_X1  g0941(.A(new_n352), .B(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n322), .A2(new_n859), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1142), .B(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n895), .A2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n884), .A2(G330), .A3(new_n893), .A4(new_n1144), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1146), .A2(new_n915), .A3(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n915), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n1001), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1144), .A2(new_n731), .B1(new_n209), .B2(new_n839), .ZN(new_n1152));
  INV_X1    g0952(.A(G124), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n257), .B1(new_n745), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n764), .A2(new_n316), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n814), .A2(new_n1107), .B1(new_n970), .B2(new_n742), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(G125), .C2(new_n748), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n1114), .B2(new_n766), .C1(new_n830), .C2(new_n773), .ZN(new_n1158));
  AOI211_X1 g0958(.A(G41), .B(new_n1154), .C1(new_n1158), .C2(KEYINPUT59), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(KEYINPUT59), .B2(new_n1158), .C1(new_n975), .C2(new_n757), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n209), .B1(new_n261), .B2(G41), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n742), .A2(new_n360), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n768), .A2(G97), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1162), .A2(new_n969), .A3(new_n1005), .A4(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(G41), .B1(new_n748), .B2(G116), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n326), .B1(new_n746), .B2(G283), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(new_n535), .C2(new_n766), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n757), .A2(new_n229), .ZN(new_n1168));
  NOR3_X1   g0968(.A1(new_n1164), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  XOR2_X1   g0969(.A(new_n1169), .B(KEYINPUT58), .Z(new_n1170));
  NAND3_X1  g0970(.A1(new_n1160), .A2(new_n1161), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n734), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1152), .A2(new_n788), .A3(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT119), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1151), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1150), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n683), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1150), .A2(new_n1176), .A3(KEYINPUT57), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1175), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(G375));
  NAND2_X1  g0982(.A1(new_n1135), .A2(new_n1001), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1083), .A2(new_n730), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n814), .A2(new_n975), .B1(new_n764), .B2(new_n209), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G128), .B2(new_n746), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1168), .A2(new_n386), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n1186), .B(new_n1187), .C1(new_n316), .C2(new_n742), .ZN(new_n1188));
  XNOR2_X1  g0988(.A(new_n1188), .B(KEYINPUT120), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G132), .B2(new_n748), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1190), .B1(new_n970), .B2(new_n766), .C1(new_n773), .C2(new_n1107), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n386), .B1(new_n819), .B2(new_n760), .C1(new_n757), .C2(new_n284), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n745), .A2(new_n449), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n535), .A2(new_n742), .B1(new_n766), .B2(new_n816), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1192), .A2(new_n1004), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n221), .B2(new_n814), .C1(new_n211), .C2(new_n773), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1069), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n839), .A2(new_n215), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1184), .A2(new_n1198), .A3(new_n788), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1183), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT121), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1183), .A2(KEYINPUT121), .A3(new_n1200), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1125), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1137), .A2(new_n960), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1205), .A2(new_n1207), .ZN(G381));
  NAND2_X1  g1008(.A1(new_n1181), .A2(new_n1139), .ZN(new_n1209));
  OR3_X1    g1009(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(G387), .A2(G384), .A3(G381), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(G407));
  OAI211_X1 g1013(.A(G407), .B(G213), .C1(G343), .C2(new_n1209), .ZN(G409));
  INV_X1    g1014(.A(new_n1173), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1150), .A2(new_n1176), .A3(new_n960), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(KEYINPUT122), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT122), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1150), .A2(new_n1176), .A3(new_n1218), .A4(new_n960), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1217), .A2(new_n1139), .A3(new_n1151), .A4(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(G213), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1221), .A2(G343), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1220), .B(new_n1223), .C1(new_n1181), .C2(new_n1139), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT60), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1206), .A2(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(KEYINPUT123), .A3(new_n1137), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1125), .A2(new_n1127), .A3(new_n1130), .A4(KEYINPUT60), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT124), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1128), .A2(new_n1083), .B1(new_n1087), .B2(new_n902), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1232), .A2(new_n1081), .B1(new_n1126), .B2(new_n1092), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1233), .A2(KEYINPUT124), .A3(KEYINPUT60), .A4(new_n1125), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1231), .A2(new_n1234), .A3(new_n1036), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT123), .B1(new_n1226), .B2(new_n1137), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1228), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1238));
  INV_X1    g1038(.A(G384), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT123), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT60), .B1(new_n1233), .B2(new_n1125), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1242), .B1(new_n1243), .B2(new_n1131), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1244), .A3(new_n1036), .A4(new_n1227), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G384), .B1(new_n1245), .B2(new_n1205), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1240), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(KEYINPUT62), .B1(new_n1224), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1222), .A2(G2897), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1240), .B2(new_n1246), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1239), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1245), .A2(G384), .A3(new_n1205), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1250), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1251), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT61), .B1(new_n1224), .B2(new_n1256), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1220), .A2(new_n1223), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT62), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1260), .A2(new_n1036), .A3(new_n1180), .ZN(new_n1261));
  OAI21_X1  g1061(.A(G378), .B1(new_n1261), .B2(new_n1175), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1258), .A2(new_n1259), .A3(new_n1247), .A4(new_n1262), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1249), .A2(new_n1257), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT126), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(G390), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1044), .B(KEYINPUT126), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1266), .B(new_n1267), .C1(new_n998), .C2(new_n999), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(new_n794), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n965), .A2(new_n997), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(G390), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1268), .A2(new_n1270), .A3(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1271), .A2(G390), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1271), .A2(G390), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1269), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1224), .A2(new_n1248), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1240), .A2(new_n1246), .A3(new_n1250), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1254), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1280));
  OAI21_X1  g1080(.A(KEYINPUT125), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT125), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1251), .A2(new_n1255), .A3(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1281), .A2(new_n1224), .A3(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1278), .B1(new_n1284), .B2(KEYINPUT63), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1258), .A2(KEYINPUT63), .A3(new_n1247), .A4(new_n1262), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT61), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1286), .A2(new_n1287), .A3(new_n1277), .ZN(new_n1288));
  OAI22_X1  g1088(.A1(new_n1264), .A2(new_n1277), .B1(new_n1285), .B2(new_n1288), .ZN(G405));
  NAND2_X1  g1089(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1175), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1290), .A2(new_n1139), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1139), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1248), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1262), .A2(new_n1209), .A3(new_n1247), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT127), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1294), .A2(new_n1296), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1277), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1294), .A2(new_n1295), .A3(new_n1296), .A4(KEYINPUT127), .ZN(new_n1302));
  AND3_X1   g1102(.A1(new_n1299), .A2(new_n1301), .A3(new_n1302), .ZN(G402));
endmodule


