//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1285,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n206), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n225), .A2(G50), .A3(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI211_X1 g0028(.A(new_n209), .B(new_n217), .C1(new_n224), .C2(new_n228), .ZN(G361));
  XOR2_X1   g0029(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n230));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G226), .B(G232), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  INV_X1    g0040(.A(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT67), .B(G107), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n202), .A2(G68), .ZN(new_n245));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n244), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(KEYINPUT7), .A3(new_n218), .ZN(new_n257));
  AOI21_X1  g0057(.A(KEYINPUT7), .B1(new_n222), .B2(new_n256), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(KEYINPUT77), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT7), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT64), .B(G20), .ZN(new_n261));
  XNOR2_X1  g0061(.A(KEYINPUT3), .B(G33), .ZN(new_n262));
  OAI211_X1 g0062(.A(KEYINPUT77), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(G68), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G58), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n246), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n267), .A2(new_n201), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n268), .A2(G20), .B1(G159), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n265), .A2(KEYINPUT16), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n256), .A2(new_n260), .A3(new_n218), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n219), .A2(new_n221), .B1(new_n253), .B2(new_n255), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n272), .B1(new_n273), .B2(new_n260), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n270), .B1(new_n274), .B2(new_n246), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT16), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT70), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND4_X1  g0080(.A1(KEYINPUT70), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(new_n223), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n271), .A2(new_n277), .A3(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G13), .A3(G20), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n285), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n218), .A2(G1), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n289), .B1(new_n292), .B2(new_n285), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G41), .ZN(new_n295));
  INV_X1    g0095(.A(G45), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g0097(.A1(G1), .A2(G13), .ZN(new_n298));
  NAND2_X1  g0098(.A1(G33), .A2(G41), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n286), .A2(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G232), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n286), .B(G274), .C1(G41), .C2(G45), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT68), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT68), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n297), .A2(new_n304), .A3(new_n286), .A4(G274), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n253), .A2(new_n255), .A3(G226), .A4(G1698), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT78), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n262), .A2(KEYINPUT78), .A3(G226), .A4(G1698), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G87), .ZN(new_n312));
  INV_X1    g0112(.A(G1698), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n262), .A2(G223), .A3(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n310), .A2(new_n311), .A3(new_n312), .A4(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n298), .A2(new_n299), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT69), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT69), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n298), .A2(new_n318), .A3(new_n299), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n307), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(G200), .B2(new_n321), .ZN(new_n324));
  NAND2_X1  g0124(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n325));
  AND4_X1   g0125(.A1(new_n283), .A2(new_n294), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n283), .A2(new_n294), .A3(new_n324), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT80), .B(KEYINPUT17), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n315), .A2(new_n320), .ZN(new_n330));
  OAI21_X1  g0130(.A(G169), .B1(new_n330), .B2(new_n307), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n321), .A2(G179), .ZN(new_n332));
  AOI221_X4 g0132(.A(KEYINPUT18), .B1(new_n331), .B2(new_n332), .C1(new_n283), .C2(new_n294), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT18), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n283), .A2(new_n294), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n332), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT79), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n282), .ZN(new_n339));
  INV_X1    g0139(.A(new_n270), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT77), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n273), .B2(KEYINPUT7), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(new_n263), .A3(new_n257), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n340), .B1(new_n343), .B2(G68), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n339), .B1(new_n344), .B2(KEYINPUT16), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n293), .B1(new_n345), .B2(new_n277), .ZN(new_n346));
  INV_X1    g0146(.A(new_n336), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT18), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT79), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n335), .A2(new_n334), .A3(new_n336), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n329), .B1(new_n338), .B2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT71), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n261), .B2(new_n252), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n222), .A2(KEYINPUT71), .A3(G33), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G150), .ZN(new_n357));
  INV_X1    g0157(.A(new_n269), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n356), .A2(new_n284), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT72), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n359), .A2(new_n360), .B1(G20), .B2(new_n203), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n339), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n288), .A2(G50), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n364), .B1(new_n292), .B2(G50), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n365), .A2(KEYINPUT73), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(KEYINPUT73), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT9), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT9), .B1(new_n363), .B2(new_n368), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n262), .A2(G222), .A3(new_n313), .ZN(new_n374));
  INV_X1    g0174(.A(G77), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n262), .A2(G1698), .ZN(new_n376));
  INV_X1    g0176(.A(G223), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n374), .B1(new_n375), .B2(new_n262), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n320), .ZN(new_n379));
  INV_X1    g0179(.A(new_n306), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(G226), .B2(new_n300), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(new_n322), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n383), .A2(KEYINPUT75), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(KEYINPUT75), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n384), .A2(new_n385), .B1(G200), .B2(new_n382), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n373), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT10), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT10), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n373), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G169), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n382), .A2(new_n392), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n393), .B1(G179), .B2(new_n382), .C1(new_n363), .C2(new_n368), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n262), .A2(G232), .A3(new_n313), .ZN(new_n395));
  INV_X1    g0195(.A(G107), .ZN(new_n396));
  INV_X1    g0196(.A(G238), .ZN(new_n397));
  OAI221_X1 g0197(.A(new_n395), .B1(new_n396), .B2(new_n262), .C1(new_n376), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n320), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n380), .B1(G244), .B2(new_n300), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n401), .A2(G179), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(new_n392), .B2(new_n401), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT15), .B(G87), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n356), .A2(new_n404), .B1(new_n358), .B2(new_n284), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n405), .A2(new_n282), .B1(new_n375), .B2(new_n288), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n339), .A2(new_n222), .ZN(new_n407));
  OAI21_X1  g0207(.A(G77), .B1(new_n407), .B2(new_n291), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n401), .A2(G200), .ZN(new_n411));
  AND3_X1   g0211(.A1(new_n406), .A2(KEYINPUT74), .A3(new_n408), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT74), .B1(new_n406), .B2(new_n408), .ZN(new_n413));
  OAI221_X1 g0213(.A(new_n411), .B1(new_n322), .B2(new_n401), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n354), .A2(new_n355), .A3(G77), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n269), .A2(G50), .B1(G20), .B2(new_n246), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(KEYINPUT11), .B1(new_n417), .B2(new_n282), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT11), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n419), .B(new_n339), .C1(new_n415), .C2(new_n416), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n288), .A2(new_n246), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT12), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n292), .B2(new_n246), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n418), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n253), .A2(new_n255), .A3(G232), .A4(G1698), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n253), .A2(new_n255), .A3(G226), .A4(new_n313), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G97), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n320), .ZN(new_n430));
  AOI22_X1  g0230(.A1(G238), .A2(new_n300), .B1(new_n303), .B2(new_n305), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT13), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT13), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n430), .A2(new_n434), .A3(new_n431), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(G179), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n392), .B1(new_n433), .B2(new_n435), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT14), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n430), .A2(new_n434), .A3(new_n431), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n434), .B1(new_n430), .B2(new_n431), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n438), .B(G169), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n425), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT76), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n440), .A2(new_n441), .ZN(new_n446));
  INV_X1    g0246(.A(G200), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(G190), .ZN(new_n449));
  OAI211_X1 g0249(.A(KEYINPUT76), .B(G200), .C1(new_n440), .C2(new_n441), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n448), .A2(new_n424), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  AND4_X1   g0251(.A1(new_n410), .A2(new_n414), .A3(new_n444), .A4(new_n451), .ZN(new_n452));
  AND4_X1   g0252(.A1(new_n352), .A2(new_n391), .A3(new_n394), .A4(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(KEYINPUT23), .A2(G107), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n261), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(KEYINPUT23), .A2(G107), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n455), .B(new_n456), .C1(G20), .C2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n222), .A2(new_n262), .A3(G87), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n461), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n463), .A2(G87), .A3(new_n222), .A4(new_n262), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n459), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT24), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n339), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n458), .B1(new_n464), .B2(new_n462), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT24), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n287), .B1(G1), .B2(new_n252), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n282), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G107), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n287), .A2(G107), .ZN(new_n474));
  XNOR2_X1  g0274(.A(new_n474), .B(KEYINPUT25), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT86), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n473), .A2(new_n475), .A3(KEYINPUT86), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n468), .A2(new_n470), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n286), .B(G45), .C1(new_n295), .C2(KEYINPUT5), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT5), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G41), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n316), .B(G264), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n253), .A2(new_n255), .A3(G250), .A4(new_n313), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT87), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n262), .A2(KEYINPUT87), .A3(G250), .A4(new_n313), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G294), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n262), .A2(G257), .A3(G1698), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n488), .A2(new_n489), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n485), .B1(new_n492), .B2(new_n320), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT88), .ZN(new_n494));
  INV_X1    g0294(.A(new_n483), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n286), .A2(G45), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n482), .A2(G41), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n495), .A2(new_n497), .A3(G274), .A4(new_n498), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n493), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n494), .B1(new_n493), .B2(new_n499), .ZN(new_n501));
  OAI21_X1  g0301(.A(G169), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n493), .A2(new_n499), .ZN(new_n503));
  INV_X1    g0303(.A(G179), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n480), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n478), .A2(new_n479), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n282), .B1(new_n469), .B2(KEYINPUT24), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n466), .A2(new_n467), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n503), .A2(KEYINPUT88), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n493), .A2(new_n494), .A3(new_n499), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n512), .A2(new_n322), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n503), .A2(new_n447), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n507), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT21), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n253), .A2(new_n255), .A3(G264), .A4(G1698), .ZN(new_n519));
  INV_X1    g0319(.A(G303), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(new_n262), .ZN(new_n521));
  INV_X1    g0321(.A(G257), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n256), .A2(new_n522), .A3(G1698), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n320), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n316), .B(G270), .C1(new_n481), .C2(new_n483), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n525), .A2(new_n499), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G169), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n290), .A2(G13), .B1(new_n286), .B2(G33), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n298), .B1(new_n279), .B2(new_n278), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n529), .A2(new_n530), .A3(G116), .A4(new_n281), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(G116), .B2(new_n287), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT20), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G283), .ZN(new_n534));
  INV_X1    g0334(.A(G97), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n534), .B1(new_n535), .B2(G33), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n261), .A2(new_n536), .B1(new_n218), .B2(G116), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n533), .B1(new_n339), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n536), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n539), .A2(new_n222), .B1(G20), .B2(new_n241), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n540), .A2(KEYINPUT20), .A3(new_n282), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n532), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n518), .B1(new_n528), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT84), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n524), .A2(new_n526), .A3(G179), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n542), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n287), .A2(G116), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n547), .B1(new_n472), .B2(G116), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n339), .A2(new_n537), .A3(new_n533), .ZN(new_n549));
  AOI21_X1  g0349(.A(KEYINPUT20), .B1(new_n540), .B2(new_n282), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n551), .A2(KEYINPUT21), .A3(G169), .A4(new_n527), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n524), .A2(new_n526), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n551), .A2(new_n553), .A3(KEYINPUT84), .A4(G179), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n543), .A2(new_n546), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n553), .A2(new_n447), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n527), .A2(new_n322), .ZN(new_n557));
  NOR3_X1   g0357(.A1(new_n556), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n497), .A2(G274), .ZN(new_n560));
  INV_X1    g0360(.A(new_n316), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n496), .A2(G250), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n262), .A2(G244), .A3(G1698), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G33), .A2(G116), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n253), .A2(new_n255), .A3(G238), .A4(new_n313), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n567), .B2(new_n320), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(new_n447), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(G190), .B2(new_n568), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n404), .A2(new_n288), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n472), .A2(G87), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G97), .A2(G107), .ZN(new_n573));
  INV_X1    g0373(.A(G87), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT19), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n428), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n575), .B1(new_n261), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n222), .A2(new_n262), .A3(G68), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n354), .A2(new_n355), .A3(G97), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n580), .B1(new_n581), .B2(new_n576), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n571), .B(new_n572), .C1(new_n582), .C2(new_n339), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n568), .A2(G169), .ZN(new_n585));
  AOI211_X1 g0385(.A(G179), .B(new_n563), .C1(new_n567), .C2(new_n320), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n404), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n472), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n589), .B(new_n571), .C1(new_n582), .C2(new_n339), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n570), .A2(new_n584), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT81), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n358), .A2(new_n375), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n396), .A2(KEYINPUT6), .A3(G97), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT6), .ZN(new_n597));
  XNOR2_X1  g0397(.A(G97), .B(G107), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n592), .B(new_n594), .C1(new_n599), .C2(new_n222), .ZN(new_n600));
  AND2_X1   g0400(.A1(G97), .A2(G107), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n597), .B1(new_n601), .B2(new_n573), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n222), .B1(new_n602), .B2(new_n595), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT81), .B1(new_n603), .B2(new_n593), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n272), .B(G107), .C1(new_n273), .C2(new_n260), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n600), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n282), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n287), .A2(new_n535), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n472), .B2(new_n535), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT82), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT82), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(new_n608), .C1(new_n472), .C2(new_n535), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n316), .B1(new_n481), .B2(new_n483), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n499), .B1(new_n615), .B2(new_n522), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n253), .A2(new_n255), .A3(G244), .A4(new_n313), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT4), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .A4(new_n313), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n262), .A2(G250), .A3(G1698), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n534), .A4(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n616), .B1(new_n622), .B2(new_n320), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(G169), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n616), .A2(KEYINPUT83), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT83), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n499), .B(new_n626), .C1(new_n615), .C2(new_n522), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n622), .A2(new_n320), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n628), .A2(new_n504), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n614), .A2(new_n624), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(G200), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n623), .A2(G190), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n633), .A2(new_n613), .A3(new_n607), .A4(new_n634), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n591), .A2(new_n631), .A3(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n453), .A2(new_n517), .A3(new_n559), .A4(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n516), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n636), .B(new_n638), .C1(new_n507), .C2(new_n555), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n585), .A2(new_n586), .ZN(new_n641));
  INV_X1    g0441(.A(new_n590), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n568), .A2(G190), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n447), .B2(new_n568), .ZN(new_n644));
  OAI22_X1  g0444(.A1(new_n641), .A2(new_n642), .B1(new_n583), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n640), .B1(new_n645), .B2(new_n631), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n614), .A2(new_n624), .A3(new_n630), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n591), .A2(new_n647), .A3(KEYINPUT26), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n646), .A2(new_n648), .B1(new_n590), .B2(new_n587), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n639), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n453), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n394), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n333), .A2(new_n337), .ZN(new_n653));
  INV_X1    g0453(.A(new_n410), .ZN(new_n654));
  OAI21_X1  g0454(.A(G169), .B1(new_n440), .B2(new_n441), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT14), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n442), .A3(new_n436), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n654), .A2(new_n451), .B1(new_n425), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n653), .B1(new_n658), .B2(new_n329), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n652), .B1(new_n391), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n651), .A2(new_n660), .ZN(G369));
  OR2_X1    g0461(.A1(new_n559), .A2(KEYINPUT90), .ZN(new_n662));
  INV_X1    g0462(.A(G213), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n222), .A2(new_n286), .A3(G13), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(KEYINPUT27), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT27), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n222), .A2(new_n666), .A3(new_n286), .A4(G13), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT89), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT89), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n665), .A2(new_n670), .A3(new_n667), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n669), .A2(G343), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(new_n542), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n559), .A2(KEYINPUT90), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n662), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n555), .A2(new_n673), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(KEYINPUT91), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n517), .B1(new_n480), .B2(new_n672), .ZN(new_n681));
  INV_X1    g0481(.A(new_n672), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n507), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n555), .A2(new_n672), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n686), .A2(new_n507), .A3(new_n516), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n507), .B2(new_n672), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n685), .A2(new_n688), .ZN(G399));
  INV_X1    g0489(.A(new_n207), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n575), .A2(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n227), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n682), .B1(new_n639), .B2(new_n649), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT93), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n635), .A2(new_n631), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n701), .B1(new_n635), .B2(new_n631), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n591), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n638), .B1(new_n507), .B2(new_n555), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n649), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n700), .B1(new_n706), .B2(new_n672), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n699), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n517), .A2(new_n559), .A3(new_n636), .A4(new_n672), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n567), .A2(new_n320), .ZN(new_n710));
  INV_X1    g0510(.A(new_n563), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n545), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n713), .A2(KEYINPUT30), .A3(new_n493), .A4(new_n623), .ZN(new_n714));
  AOI21_X1  g0514(.A(G179), .B1(new_n524), .B2(new_n526), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n632), .A2(new_n503), .A3(new_n712), .A4(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT30), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n493), .A2(new_n623), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n568), .A2(G179), .A3(new_n524), .A4(new_n526), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n714), .A2(new_n716), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n682), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g0524(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n725));
  OAI211_X1 g0525(.A(new_n709), .B(new_n724), .C1(new_n722), .C2(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n708), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n696), .B1(new_n728), .B2(G1), .ZN(G364));
  NOR2_X1   g0529(.A1(new_n679), .A2(G330), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n222), .A2(G13), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n286), .B1(new_n731), .B2(G45), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n730), .B(new_n680), .C1(new_n692), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n732), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n691), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n690), .A2(new_n256), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G355), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(G116), .B2(new_n207), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n256), .A2(new_n207), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT94), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n296), .B2(new_n228), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n250), .A2(new_n296), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n738), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n223), .B1(G20), .B2(new_n392), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n735), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  NOR4_X1   g0551(.A1(new_n218), .A2(new_n322), .A3(new_n447), .A4(G179), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n256), .B1(new_n752), .B2(G87), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n322), .A2(G179), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n222), .A2(new_n754), .ZN(new_n755));
  NOR4_X1   g0555(.A1(new_n222), .A2(G179), .A3(G190), .A4(new_n447), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n753), .B1(new_n535), .B2(new_n755), .C1(new_n757), .C2(new_n396), .ZN(new_n758));
  NOR3_X1   g0558(.A1(G179), .A2(G190), .A3(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n261), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G159), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT32), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n261), .A2(G179), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT96), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n758), .B(new_n763), .C1(new_n767), .C2(G77), .ZN(new_n768));
  INV_X1    g0568(.A(new_n764), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(KEYINPUT97), .A3(G200), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT97), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(new_n764), .B2(new_n447), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n770), .A2(G190), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n770), .A2(new_n322), .A3(new_n772), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G50), .A2(new_n774), .B1(new_n776), .B2(G68), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n769), .A2(G190), .A3(new_n447), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT95), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT95), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n768), .B(new_n777), .C1(new_n266), .C2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT98), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n761), .A2(G329), .ZN(new_n786));
  INV_X1    g0586(.A(G283), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n757), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G294), .ZN(new_n789));
  INV_X1    g0589(.A(new_n752), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n256), .B1(new_n755), .B2(new_n789), .C1(new_n790), .C2(new_n520), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G311), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n793), .B2(new_n766), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G322), .B2(new_n781), .ZN(new_n795));
  INV_X1    g0595(.A(G326), .ZN(new_n796));
  XOR2_X1   g0596(.A(KEYINPUT33), .B(G317), .Z(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(new_n796), .B2(new_n773), .C1(new_n775), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n783), .A2(new_n784), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n785), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n751), .B1(new_n800), .B2(new_n748), .ZN(new_n801));
  INV_X1    g0601(.A(new_n747), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n678), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT99), .Z(new_n804));
  NOR2_X1   g0604(.A1(new_n733), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  NOR2_X1   g0606(.A1(new_n748), .A2(new_n745), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n775), .B(KEYINPUT100), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n787), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n256), .B1(new_n790), .B2(new_n396), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n756), .A2(G87), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n793), .B2(new_n760), .ZN(new_n813));
  INV_X1    g0613(.A(new_n755), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n811), .B(new_n813), .C1(G97), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n767), .A2(G116), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(new_n789), .C2(new_n782), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n810), .B(new_n817), .C1(G303), .C2(new_n774), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n767), .A2(G159), .B1(new_n781), .B2(G143), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n819), .B1(new_n820), .B2(new_n773), .C1(new_n357), .C2(new_n775), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT34), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n756), .A2(G68), .B1(G50), .B2(new_n752), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n266), .B2(new_n755), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n761), .A2(G132), .ZN(new_n825));
  AOI21_X1  g0625(.A(KEYINPUT101), .B1(new_n825), .B2(new_n262), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n825), .A2(KEYINPUT101), .A3(new_n262), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n818), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n748), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n735), .B1(G77), .B2(new_n808), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT102), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n682), .A2(new_n409), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n414), .A2(new_n410), .A3(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT103), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n403), .A2(new_n837), .A3(new_n409), .A4(new_n682), .ZN(new_n838));
  INV_X1    g0638(.A(new_n402), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n401), .A2(new_n392), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n839), .A2(new_n682), .A3(new_n409), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT103), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n836), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n833), .B(new_n834), .C1(new_n745), .C2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n698), .A2(new_n845), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n502), .A2(new_n506), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n555), .B1(new_n848), .B2(new_n511), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n591), .A2(new_n631), .A3(new_n635), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n849), .A2(new_n516), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n587), .A2(new_n590), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n645), .A2(new_n640), .A3(new_n631), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT26), .B1(new_n591), .B2(new_n647), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n672), .B(new_n844), .C1(new_n851), .C2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n847), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n727), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n735), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n727), .A2(new_n847), .A3(new_n856), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n846), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G384));
  INV_X1    g0663(.A(new_n599), .ZN(new_n864));
  OAI211_X1 g0664(.A(G116), .B(new_n224), .C1(new_n864), .C2(KEYINPUT35), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n865), .B1(KEYINPUT35), .B2(new_n864), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT36), .ZN(new_n867));
  OR3_X1    g0667(.A1(new_n227), .A2(new_n375), .A3(new_n267), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n286), .B(G13), .C1(new_n868), .C2(new_n245), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT108), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT108), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n721), .A2(new_n873), .A3(KEYINPUT31), .A4(new_n682), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n722), .A2(new_n725), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n709), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n453), .A2(G330), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n424), .A2(new_n672), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n444), .A2(new_n451), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT105), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT104), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n657), .A2(new_n884), .A3(new_n880), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n884), .B1(new_n657), .B2(new_n880), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n882), .B(new_n883), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n657), .A2(new_n880), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT104), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n885), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n883), .B1(new_n892), .B2(new_n882), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n877), .B(new_n844), .C1(new_n889), .C2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT37), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n669), .A2(new_n671), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n331), .A2(new_n332), .A3(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n327), .B(new_n896), .C1(new_n346), .C2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT106), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n331), .A2(new_n332), .A3(new_n897), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n335), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n903), .A2(KEYINPUT106), .A3(new_n896), .A4(new_n327), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n345), .B1(KEYINPUT16), .B2(new_n344), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n898), .B1(new_n906), .B2(new_n294), .ZN(new_n907));
  INV_X1    g0707(.A(new_n327), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT37), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n906), .A2(new_n294), .ZN(new_n911));
  INV_X1    g0711(.A(new_n897), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n910), .B(KEYINPUT38), .C1(new_n352), .C2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT38), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n896), .B1(new_n903), .B2(new_n327), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n901), .B2(new_n904), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n335), .A2(new_n912), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n327), .A2(new_n328), .ZN(new_n919));
  INV_X1    g0719(.A(new_n325), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n919), .B1(new_n327), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n918), .B1(new_n653), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n915), .B1(new_n917), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n914), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n879), .B1(new_n895), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n882), .B1(new_n886), .B2(new_n887), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT105), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n888), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n928), .A2(new_n879), .A3(new_n844), .A4(new_n877), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n338), .A2(new_n351), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n913), .B1(new_n930), .B2(new_n921), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n911), .A2(new_n902), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n896), .B1(new_n932), .B2(new_n327), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n901), .B2(new_n904), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n915), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n929), .B1(new_n914), .B2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n925), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(G330), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n878), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT109), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n935), .A2(new_n914), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n894), .B1(new_n914), .B2(new_n923), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n942), .A2(new_n929), .B1(new_n943), .B2(new_n879), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n944), .A2(new_n453), .A3(new_n877), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n444), .A2(new_n682), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT39), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n935), .B2(new_n914), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n914), .A2(new_n948), .A3(new_n923), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n653), .A2(new_n912), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n410), .A2(new_n682), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n697), .B2(new_n844), .ZN(new_n954));
  INV_X1    g0754(.A(new_n928), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n952), .B1(new_n941), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n951), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT107), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT107), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n951), .A2(new_n960), .A3(new_n957), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n946), .B(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n708), .A2(new_n453), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n964), .A2(new_n660), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n286), .B2(new_n731), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n963), .A2(new_n965), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n870), .B1(new_n967), .B2(new_n968), .ZN(G367));
  NOR2_X1   g0769(.A1(new_n631), .A2(new_n672), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT110), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n682), .A2(new_n614), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n702), .B2(new_n703), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n687), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT42), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n507), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n682), .B1(new_n977), .B2(new_n631), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n682), .A2(new_n583), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n591), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n980), .A2(new_n852), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n979), .B1(KEYINPUT43), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n685), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n974), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n986), .B(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n691), .B(KEYINPUT41), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n684), .B1(new_n555), .B2(new_n672), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n680), .B(KEYINPUT112), .C1(new_n687), .C2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n680), .A2(KEYINPUT112), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n992), .A2(new_n687), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n680), .A2(KEYINPUT112), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n688), .A2(new_n974), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT45), .Z(new_n1000));
  NOR2_X1   g0800(.A1(new_n688), .A2(new_n974), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT44), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT111), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n685), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n987), .A2(KEYINPUT111), .A3(new_n1003), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n998), .A2(new_n728), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n991), .B1(new_n1007), .B2(new_n728), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n989), .B1(new_n1008), .B2(new_n734), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n256), .B1(new_n755), .B2(new_n396), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n752), .A2(G116), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT46), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n756), .A2(G97), .B1(new_n761), .B2(G317), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1010), .B(new_n1014), .C1(G303), .C2(new_n781), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n767), .A2(G283), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(new_n793), .C2(new_n773), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n809), .A2(new_n789), .ZN(new_n1018));
  INV_X1    g0818(.A(G159), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n809), .A2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n767), .A2(G50), .B1(new_n781), .B2(G150), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n774), .A2(G143), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n761), .A2(G137), .B1(G58), .B2(new_n752), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(KEYINPUT113), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n814), .A2(G68), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1025), .B(new_n262), .C1(new_n757), .C2(new_n375), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1023), .A2(KEYINPUT113), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .A4(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1017), .A2(new_n1018), .B1(new_n1020), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT47), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n830), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n1031), .B2(new_n1030), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n735), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n238), .A2(new_n740), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n750), .B1(new_n690), .B2(new_n588), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1033), .B(new_n1037), .C1(new_n802), .C2(new_n983), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1009), .A2(new_n1038), .ZN(G387));
  NAND2_X1  g0839(.A1(new_n998), .A2(new_n728), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n993), .B1(new_n708), .B2(new_n727), .C1(new_n996), .C2(new_n997), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n1041), .A3(new_n691), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n741), .B1(new_n234), .B2(G45), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n693), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n736), .ZN(new_n1045));
  AOI21_X1  g0845(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n285), .A2(new_n202), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n693), .B(new_n1046), .C1(new_n1047), .C2(KEYINPUT50), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(KEYINPUT50), .B2(new_n1047), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1045), .A2(new_n1049), .B1(G107), .B2(new_n207), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1034), .B1(new_n1050), .B2(new_n749), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n684), .B2(new_n802), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n767), .A2(G303), .B1(new_n781), .B2(G317), .ZN(new_n1053));
  INV_X1    g0853(.A(G322), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1053), .B1(new_n1054), .B2(new_n773), .C1(new_n809), .C2(new_n793), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT48), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n787), .B2(new_n755), .C1(new_n789), .C2(new_n790), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT49), .Z(new_n1058));
  OAI221_X1 g0858(.A(new_n256), .B1(new_n796), .B2(new_n760), .C1(new_n757), .C2(new_n241), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n776), .A2(new_n285), .B1(G68), .B2(new_n765), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1061), .A2(KEYINPUT114), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(KEYINPUT114), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n752), .A2(G77), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n262), .B(new_n1064), .C1(new_n757), .C2(new_n535), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n814), .A2(new_n588), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n357), .B2(new_n760), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1065), .B(new_n1067), .C1(new_n781), .C2(G50), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n774), .A2(G159), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1063), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n1058), .A2(new_n1059), .B1(new_n1062), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1052), .B1(new_n1071), .B2(new_n748), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n998), .B2(new_n734), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1042), .A2(new_n1073), .ZN(G393));
  AOI22_X1  g0874(.A1(new_n781), .A2(G311), .B1(G317), .B2(new_n774), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n755), .A2(new_n241), .B1(new_n760), .B2(new_n1054), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n256), .B1(new_n790), .B2(new_n787), .C1(new_n757), .C2(new_n396), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G294), .C2(new_n765), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1077), .B(new_n1080), .C1(new_n520), .C2(new_n809), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n781), .A2(G159), .B1(G150), .B2(new_n774), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT115), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n814), .A2(G77), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n256), .B1(new_n752), .B2(G68), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n761), .A2(G143), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n812), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n767), .B2(new_n285), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1084), .B(new_n1089), .C1(new_n202), .C2(new_n809), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1081), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n748), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n244), .A2(new_n740), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n750), .B1(G97), .B2(new_n690), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1034), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1093), .B(new_n1096), .C1(new_n974), .C2(new_n802), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n685), .B(new_n1003), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1007), .A2(new_n691), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n728), .B2(new_n998), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n1097), .B1(new_n732), .B2(new_n1099), .C1(new_n1100), .C2(new_n1101), .ZN(G390));
  NAND3_X1  g0902(.A1(new_n964), .A2(new_n660), .A3(new_n878), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n727), .A2(new_n844), .A3(new_n928), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n706), .A2(new_n672), .A3(new_n844), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n953), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n877), .A2(G330), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n955), .B1(new_n1110), .B2(new_n845), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1105), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n928), .A2(new_n844), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1113), .A2(new_n1110), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n727), .A2(new_n844), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n1115), .B2(new_n955), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1112), .B1(new_n1116), .B2(new_n954), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1104), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT117), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n856), .A2(new_n1107), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n947), .B1(new_n1120), .B2(new_n928), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n949), .A2(new_n950), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1108), .A2(new_n928), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n947), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n924), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1114), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n333), .A2(new_n337), .A3(KEYINPUT79), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n349), .B1(new_n348), .B2(new_n350), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n921), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n913), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(KEYINPUT38), .B1(new_n1131), .B2(new_n910), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n914), .ZN(new_n1133));
  OAI21_X1  g0933(.A(KEYINPUT39), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n914), .A2(new_n948), .A3(new_n923), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1124), .B1(new_n954), .B2(new_n955), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1123), .A2(new_n1124), .A3(new_n924), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n1138), .A3(new_n1105), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1119), .B1(new_n1126), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1141));
  AOI21_X1  g0941(.A(KEYINPUT117), .B1(new_n1141), .B2(new_n1114), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1118), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1105), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1122), .A2(new_n1125), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1114), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1147));
  OAI21_X1  g0947(.A(KEYINPUT117), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1126), .A2(new_n1119), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1115), .A2(new_n955), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n954), .B1(new_n1150), .B2(new_n1146), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1112), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1153), .A2(new_n1103), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1148), .A2(new_n1149), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1143), .A2(new_n1155), .A3(new_n691), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n735), .B1(new_n285), .B2(new_n808), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n949), .A2(new_n950), .A3(new_n746), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT54), .B(G143), .Z(new_n1159));
  AOI22_X1  g0959(.A1(new_n767), .A2(new_n1159), .B1(G159), .B2(new_n814), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n809), .B2(new_n820), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT118), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n1163));
  OR3_X1    g0963(.A1(new_n790), .A2(new_n357), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n790), .B2(new_n357), .ZN(new_n1165));
  INV_X1    g0965(.A(G125), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1164), .B(new_n1165), .C1(new_n1166), .C2(new_n760), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n256), .B(new_n1167), .C1(G50), .C2(new_n756), .ZN(new_n1168));
  INV_X1    g0968(.A(G128), .ZN(new_n1169));
  INV_X1    g0969(.A(G132), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1168), .B1(new_n1169), .B2(new_n773), .C1(new_n1170), .C2(new_n782), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n809), .A2(new_n396), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n256), .B1(new_n790), .B2(new_n574), .C1(new_n757), .C2(new_n246), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1085), .B1(new_n789), .B2(new_n760), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n767), .C2(G97), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n241), .B2(new_n782), .C1(new_n787), .C2(new_n773), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n1162), .A2(new_n1171), .B1(new_n1172), .B2(new_n1176), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1157), .B(new_n1158), .C1(new_n748), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1126), .A2(new_n1139), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1142), .B1(KEYINPUT117), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1178), .B1(new_n1180), .B2(new_n734), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1156), .A2(new_n1181), .ZN(G378));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n912), .B1(new_n363), .B2(new_n368), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n391), .B2(new_n394), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n373), .A2(new_n386), .A3(new_n389), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n389), .B1(new_n373), .B2(new_n386), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n394), .B(new_n1185), .C1(new_n1187), .C2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1184), .B1(new_n1186), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n394), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1185), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1194), .A2(new_n1189), .A3(new_n1183), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1191), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(new_n944), .B2(G330), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1196), .B(G330), .C1(new_n925), .C2(new_n936), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n959), .B(new_n961), .C1(new_n1197), .C2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1196), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n937), .B2(new_n938), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n951), .A2(new_n960), .A3(new_n957), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n960), .B1(new_n951), .B2(new_n957), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1202), .B(new_n1198), .C1(new_n1203), .C2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT121), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1200), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1202), .A2(new_n1198), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1208), .A2(KEYINPUT121), .A3(new_n961), .A4(new_n959), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1207), .A2(new_n734), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1201), .A2(new_n745), .ZN(new_n1211));
  AOI21_X1  g1011(.A(G50), .B1(new_n252), .B2(new_n295), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n262), .B2(G41), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT120), .Z(new_n1214));
  NOR2_X1   g1014(.A1(new_n782), .A2(new_n396), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n766), .A2(new_n404), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1025), .A2(new_n295), .A3(new_n256), .A4(new_n1064), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n756), .A2(G58), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n787), .B2(new_n760), .ZN(new_n1219));
  NOR4_X1   g1019(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n535), .B2(new_n775), .C1(new_n241), .C2(new_n773), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT58), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1214), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n814), .A2(G150), .B1(new_n752), .B2(new_n1159), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n766), .B2(new_n820), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n781), .B2(G128), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n1166), .B2(new_n773), .C1(new_n1170), .C2(new_n775), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n756), .A2(G159), .ZN(new_n1230));
  AOI211_X1 g1030(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1223), .B1(new_n1222), .B2(new_n1221), .C1(new_n1228), .C2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n748), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n807), .A2(new_n202), .ZN(new_n1235));
  AND4_X1   g1035(.A1(new_n735), .A2(new_n1211), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1210), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1155), .A2(new_n1104), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT57), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1200), .B2(new_n1205), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1241), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n691), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1239), .B1(new_n1242), .B2(new_n1246), .ZN(G375));
  INV_X1    g1047(.A(KEYINPUT122), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1153), .B2(new_n1103), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1153), .A2(new_n1248), .A3(new_n1103), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1252), .A2(new_n990), .A3(new_n1118), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n782), .A2(new_n820), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1218), .B(new_n262), .C1(new_n1019), .C2(new_n790), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n766), .A2(new_n357), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n755), .A2(new_n202), .B1(new_n760), .B2(new_n1169), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1159), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1258), .B1(new_n1170), .B2(new_n773), .C1(new_n809), .C2(new_n1259), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n809), .A2(new_n241), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n256), .B1(new_n790), .B2(new_n535), .C1(new_n757), .C2(new_n375), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1066), .B1(new_n520), .B2(new_n760), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1262), .B(new_n1263), .C1(new_n767), .C2(G107), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1264), .B1(new_n787), .B2(new_n782), .C1(new_n789), .C2(new_n773), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1260), .B1(new_n1261), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n830), .B1(new_n1266), .B2(KEYINPUT123), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(KEYINPUT123), .B2(new_n1266), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1034), .B1(new_n246), .B2(new_n807), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(new_n928), .C2(new_n746), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1270), .B1(new_n1153), .B2(new_n732), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1253), .A2(new_n1272), .ZN(G381));
  NAND3_X1  g1073(.A1(new_n1042), .A2(new_n805), .A3(new_n1073), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(G384), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(KEYINPUT124), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(G387), .A2(G390), .A3(G381), .ZN(new_n1277));
  INV_X1    g1077(.A(G378), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1103), .B1(new_n1180), .B2(new_n1117), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1243), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n692), .B1(new_n1241), .B2(new_n1244), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1238), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1276), .A2(new_n1277), .A3(new_n1278), .A4(new_n1283), .ZN(G407));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1278), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G407), .B(G213), .C1(G343), .C2(new_n1285), .ZN(G409));
  NOR2_X1   g1086(.A1(new_n663), .A2(G343), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1200), .A2(new_n1205), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1236), .B1(new_n1288), .B2(new_n734), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1289), .A2(new_n1156), .A3(new_n1181), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1240), .A2(new_n990), .A3(new_n1241), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1287), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n1278), .B2(new_n1283), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1153), .A2(new_n1103), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT60), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n691), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1118), .A2(KEYINPUT60), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1252), .B2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n862), .B1(new_n1298), .B2(new_n1271), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1251), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1297), .B1(new_n1300), .B2(new_n1249), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1296), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(G384), .A3(new_n1272), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1299), .A2(new_n1304), .A3(G2897), .A4(new_n1287), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1287), .A2(G2897), .ZN(new_n1306));
  AOI21_X1  g1106(.A(G384), .B1(new_n1303), .B2(new_n1272), .ZN(new_n1307));
  AOI211_X1 g1107(.A(new_n862), .B(new_n1271), .C1(new_n1301), .C2(new_n1302), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1306), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1305), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT61), .B1(new_n1293), .B2(new_n1310), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1312));
  OAI211_X1 g1112(.A(new_n1292), .B(new_n1312), .C1(new_n1278), .C2(new_n1283), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(KEYINPUT62), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G375), .A2(G378), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT62), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1315), .A2(new_n1316), .A3(new_n1312), .A4(new_n1292), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1311), .A2(new_n1314), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1274), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n805), .B1(new_n1042), .B2(new_n1073), .ZN(new_n1320));
  OAI21_X1  g1120(.A(KEYINPUT126), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1320), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT126), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1322), .A2(new_n1323), .A3(new_n1274), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1321), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(G390), .A2(new_n1038), .A3(new_n1009), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(G390), .B1(new_n1009), .B2(new_n1038), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1325), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(G390), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(G387), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1331), .A2(new_n1321), .A3(new_n1324), .A4(new_n1326), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1329), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1318), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1313), .A2(KEYINPUT63), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT63), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1315), .A2(new_n1337), .A3(new_n1312), .A4(new_n1292), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(KEYINPUT61), .B1(new_n1329), .B2(new_n1332), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1278), .B1(new_n1341), .B2(new_n1239), .ZN(new_n1342));
  NOR3_X1   g1142(.A1(new_n1279), .A2(new_n1280), .A3(new_n991), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1289), .A2(new_n1156), .A3(new_n1181), .ZN(new_n1344));
  OAI22_X1  g1144(.A1(new_n1343), .A2(new_n1344), .B1(new_n663), .B2(G343), .ZN(new_n1345));
  OAI21_X1  g1145(.A(KEYINPUT125), .B1(new_n1342), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT125), .ZN(new_n1347));
  OAI211_X1 g1147(.A(new_n1292), .B(new_n1347), .C1(new_n1278), .C2(new_n1283), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1346), .A2(new_n1310), .A3(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1339), .A2(new_n1340), .A3(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1335), .A2(new_n1350), .ZN(G405));
  INV_X1    g1151(.A(new_n1285), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1312), .B1(new_n1352), .B2(new_n1342), .ZN(new_n1353));
  OAI211_X1 g1153(.A(new_n1315), .B(new_n1285), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1334), .A2(new_n1353), .A3(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1353), .A2(new_n1354), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1333), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1355), .A2(new_n1357), .ZN(G402));
endmodule


