//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT75), .ZN(new_n203));
  OR2_X1    g002(.A1(G197gat), .A2(G204gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  NAND2_X1  g005(.A1(G211gat), .A2(G218gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n203), .A2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n202), .A2(KEYINPUT75), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n202), .A2(KEYINPUT75), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n208), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  INV_X1    g015(.A(G162gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT78), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G141gat), .B(G148gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n220), .B1(G155gat), .B2(G162gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n218), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g021(.A(G155gat), .B(G162gat), .Z(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n222), .B(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n215), .B1(new_n226), .B2(KEYINPUT29), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT29), .B1(new_n210), .B2(new_n213), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n225), .B1(new_n228), .B2(KEYINPUT3), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT83), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G228gat), .ZN(new_n233));
  INV_X1    g032(.A(G233gat), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G22gat), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n230), .B(new_n231), .C1(new_n233), .C2(new_n234), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT84), .ZN(new_n240));
  XNOR2_X1  g039(.A(G78gat), .B(G106gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT31), .B(G50gat), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n241), .B(new_n242), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n236), .A2(new_n238), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(G22gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n239), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g047(.A1(new_n240), .A2(new_n246), .A3(new_n239), .A4(new_n243), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G1gat), .B(G29gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(KEYINPUT0), .ZN(new_n252));
  XNOR2_X1  g051(.A(G57gat), .B(G85gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n222), .A2(new_n223), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n222), .A2(new_n223), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n261));
  XNOR2_X1  g060(.A(G113gat), .B(G120gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(KEYINPUT1), .ZN(new_n263));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(new_n261), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT81), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n225), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n264), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n263), .B(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT4), .B1(new_n258), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n268), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n269), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n258), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n225), .A2(new_n265), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n276), .B(KEYINPUT81), .C1(new_n277), .C2(KEYINPUT4), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n267), .B1(new_n274), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G225gat), .A2(G233gat), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n279), .A2(KEYINPUT39), .A3(new_n280), .ZN(new_n281));
  OR2_X1    g080(.A1(new_n279), .A2(new_n280), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT39), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n258), .A2(new_n272), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n225), .A2(new_n265), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n283), .B1(new_n287), .B2(new_n280), .ZN(new_n288));
  AOI211_X1 g087(.A(new_n255), .B(new_n281), .C1(new_n282), .C2(new_n288), .ZN(new_n289));
  OR2_X1    g088(.A1(KEYINPUT85), .A2(KEYINPUT40), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT5), .B1(new_n287), .B2(new_n280), .ZN(new_n292));
  INV_X1    g091(.A(new_n280), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n293), .B1(new_n284), .B2(new_n269), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n258), .A2(KEYINPUT4), .A3(new_n272), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(new_n266), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT80), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n294), .A2(new_n266), .A3(KEYINPUT80), .A4(new_n295), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n292), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n280), .A2(new_n301), .ZN(new_n302));
  AOI211_X1 g101(.A(new_n302), .B(new_n267), .C1(new_n274), .C2(new_n278), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n255), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n305), .B1(new_n289), .B2(new_n290), .ZN(new_n306));
  NAND2_X1  g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(KEYINPUT24), .ZN(new_n309));
  INV_X1    g108(.A(G183gat), .ZN(new_n310));
  INV_X1    g109(.A(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OR3_X1    g113(.A1(new_n309), .A2(new_n314), .A3(KEYINPUT64), .ZN(new_n315));
  INV_X1    g114(.A(G169gat), .ZN(new_n316));
  INV_X1    g115(.A(G176gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(KEYINPUT65), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT65), .ZN(new_n321));
  NOR2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n321), .B1(new_n322), .B2(KEYINPUT23), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n316), .A2(new_n317), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(KEYINPUT23), .B2(new_n322), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT64), .B1(new_n309), .B2(new_n314), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n315), .A2(new_n324), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT25), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT66), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT24), .B1(new_n307), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n330), .B2(new_n307), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(new_n312), .A3(new_n313), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n324), .A2(KEYINPUT25), .A3(new_n326), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n328), .A2(new_n329), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT70), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT27), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT67), .B1(new_n339), .B2(G183gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT67), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n310), .A3(KEYINPUT27), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n342), .A3(new_n311), .ZN(new_n343));
  OAI21_X1  g142(.A(G183gat), .B1(KEYINPUT68), .B2(KEYINPUT27), .ZN(new_n344));
  AND2_X1   g143(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n338), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT27), .B(G183gat), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(KEYINPUT28), .A3(new_n311), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n337), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n337), .A3(new_n349), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n318), .A2(KEYINPUT26), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n318), .B1(new_n325), .B2(KEYINPUT26), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n355), .B2(KEYINPUT71), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT71), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n357), .B(new_n318), .C1(new_n325), .C2(KEYINPUT26), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n308), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT72), .B1(new_n353), .B2(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n347), .A2(new_n337), .A3(new_n349), .ZN(new_n361));
  OAI211_X1 g160(.A(KEYINPUT72), .B(new_n359), .C1(new_n361), .C2(new_n350), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n336), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n359), .B1(new_n361), .B2(new_n350), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT72), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n362), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(KEYINPUT76), .A3(new_n336), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n366), .A2(KEYINPUT77), .A3(new_n368), .A4(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT76), .B1(new_n372), .B2(new_n336), .ZN(new_n375));
  AOI211_X1 g174(.A(new_n365), .B(new_n335), .C1(new_n371), .C2(new_n362), .ZN(new_n376));
  NOR3_X1   g175(.A1(new_n375), .A2(new_n376), .A3(new_n367), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT77), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT29), .B1(new_n336), .B2(new_n369), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n378), .B1(new_n379), .B2(new_n368), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n214), .B(new_n374), .C1(new_n377), .C2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G8gat), .B(G36gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(G64gat), .B(G92gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OR2_X1    g184(.A1(new_n368), .A2(KEYINPUT29), .ZN(new_n386));
  NOR3_X1   g185(.A1(new_n375), .A2(new_n376), .A3(new_n386), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n336), .A2(new_n368), .A3(new_n369), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n215), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n381), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n385), .B1(new_n381), .B2(new_n389), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(KEYINPUT30), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT30), .ZN(new_n393));
  AOI211_X1 g192(.A(new_n393), .B(new_n385), .C1(new_n381), .C2(new_n389), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n291), .B(new_n306), .C1(new_n392), .C2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n300), .A2(new_n303), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n254), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n304), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n305), .A2(KEYINPUT6), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(new_n391), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n381), .A2(new_n389), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n385), .A2(KEYINPUT37), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n403), .A2(KEYINPUT37), .B1(new_n390), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT38), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n402), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT38), .B1(new_n390), .B2(new_n404), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n215), .B(new_n374), .C1(new_n377), .C2(new_n380), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n214), .B1(new_n387), .B2(new_n388), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(KEYINPUT86), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n366), .A2(new_n368), .A3(new_n373), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n412), .B(new_n378), .C1(new_n368), .C2(new_n379), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT86), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n413), .A2(new_n414), .A3(new_n215), .A4(new_n374), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(new_n415), .A3(KEYINPUT37), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n408), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n250), .B(new_n395), .C1(new_n407), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n248), .A2(new_n249), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n381), .A2(new_n389), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n384), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n393), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n304), .A2(KEYINPUT82), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT82), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n424), .B(new_n255), .C1(new_n300), .C2(new_n303), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n423), .A2(new_n397), .A3(new_n398), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n400), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n391), .A2(KEYINPUT30), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n422), .A2(new_n427), .A3(new_n390), .A4(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT74), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n364), .A2(new_n265), .ZN(new_n431));
  NAND2_X1  g230(.A1(G227gat), .A2(G233gat), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n372), .A2(new_n272), .A3(new_n336), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT34), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n434), .A2(KEYINPUT73), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n431), .A2(new_n432), .A3(new_n433), .A4(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n272), .B1(new_n372), .B2(new_n336), .ZN(new_n438));
  AOI211_X1 g237(.A(new_n265), .B(new_n335), .C1(new_n371), .C2(new_n362), .ZN(new_n439));
  INV_X1    g238(.A(new_n432), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n437), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n440), .B1(new_n438), .B2(new_n439), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT32), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  XOR2_X1   g246(.A(G15gat), .B(G43gat), .Z(new_n448));
  XNOR2_X1  g247(.A(G71gat), .B(G99gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n445), .A2(new_n447), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n450), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n444), .B(KEYINPUT32), .C1(new_n446), .C2(new_n452), .ZN(new_n453));
  AOI211_X1 g252(.A(new_n430), .B(new_n443), .C1(new_n451), .C2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n453), .A3(new_n443), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n443), .A2(new_n430), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT36), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n451), .A2(new_n453), .ZN(new_n459));
  INV_X1    g258(.A(new_n443), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT36), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n455), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n419), .A2(new_n429), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n250), .B1(new_n454), .B2(new_n457), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT35), .B1(new_n429), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n392), .A2(new_n394), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n419), .B1(new_n461), .B2(new_n455), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT35), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n467), .A2(new_n468), .A3(new_n469), .A4(new_n401), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n418), .A2(new_n464), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(G8gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(G15gat), .B(G22gat), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n473), .A2(G1gat), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT92), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT16), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n473), .B1(new_n477), .B2(G1gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n476), .B(new_n479), .Z(new_n480));
  XNOR2_X1  g279(.A(G43gat), .B(G50gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT15), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g283(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n485));
  OR2_X1    g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT87), .B(G36gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(G29gat), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n482), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n485), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n483), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT90), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n481), .A2(KEYINPUT88), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT15), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT91), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n488), .B(new_n497), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n489), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT17), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI211_X1 g301(.A(KEYINPUT17), .B(new_n489), .C1(new_n494), .C2(new_n499), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n480), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G229gat), .A2(G233gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n500), .ZN(new_n506));
  INV_X1    g305(.A(new_n480), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT18), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n504), .A2(new_n508), .A3(KEYINPUT18), .A4(new_n505), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(new_n500), .B2(new_n480), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n506), .A2(new_n513), .A3(new_n507), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n505), .B(KEYINPUT13), .Z(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n511), .A2(new_n512), .A3(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G113gat), .B(G141gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(G197gat), .ZN(new_n521));
  XOR2_X1   g320(.A(KEYINPUT11), .B(G169gat), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n523), .B(KEYINPUT12), .Z(new_n524));
  NAND2_X1  g323(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n524), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n511), .A2(new_n518), .A3(new_n526), .A4(new_n512), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(KEYINPUT94), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT94), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n519), .A2(new_n529), .A3(new_n524), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT21), .ZN(new_n532));
  XOR2_X1   g331(.A(G57gat), .B(G64gat), .Z(new_n533));
  NAND2_X1  g332(.A1(G71gat), .A2(G78gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(G71gat), .A2(G78gat), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT95), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n534), .A2(new_n539), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n534), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n543), .A2(new_n538), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n533), .B(new_n536), .C1(new_n544), .C2(new_n540), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n480), .B1(new_n532), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT97), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n546), .A2(KEYINPUT21), .ZN(new_n550));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G127gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n549), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT96), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(G155gat), .ZN(new_n558));
  XOR2_X1   g357(.A(G183gat), .B(G211gat), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT98), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n558), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n555), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G134gat), .B(G162gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n564), .B(new_n565), .Z(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G99gat), .ZN(new_n572));
  INV_X1    g371(.A(G106gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n571), .A2(new_n567), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n567), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n566), .A2(new_n576), .A3(new_n570), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(KEYINPUT100), .A3(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n577), .A2(KEYINPUT100), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT41), .ZN(new_n582));
  AND2_X1   g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  OAI22_X1  g383(.A1(new_n500), .A2(new_n581), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n492), .B(KEYINPUT90), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n496), .A2(new_n498), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT17), .B1(new_n588), .B2(new_n489), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n500), .A2(new_n501), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n580), .A2(KEYINPUT101), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT101), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n593), .A3(new_n579), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n585), .B1(new_n591), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G190gat), .B(G218gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT102), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n563), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n598), .A2(new_n599), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n584), .A2(new_n582), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n600), .ZN(new_n605));
  INV_X1    g404(.A(new_n563), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n595), .B1(new_n589), .B2(new_n590), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n585), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n601), .A2(new_n604), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n604), .B1(new_n601), .B2(new_n608), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n562), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n546), .B1(new_n578), .B2(new_n579), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n547), .B1(new_n577), .B2(new_n575), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n580), .A2(KEYINPUT10), .A3(new_n546), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(KEYINPUT103), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  OR3_X1    g421(.A1(new_n614), .A2(new_n621), .A3(new_n615), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G120gat), .B(G148gat), .Z(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT104), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n626), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n624), .A2(new_n625), .A3(new_n630), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n612), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT106), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n471), .A2(new_n531), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n427), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G1gat), .ZN(G1324gat));
  INV_X1    g441(.A(new_n467), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT16), .B(G8gat), .Z(new_n645));
  AND3_X1   g444(.A1(new_n644), .A2(KEYINPUT42), .A3(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n646), .A2(KEYINPUT107), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(KEYINPUT107), .ZN(new_n648));
  OAI21_X1  g447(.A(KEYINPUT42), .B1(new_n644), .B2(new_n472), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n644), .A2(new_n645), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n647), .B1(new_n648), .B2(new_n651), .ZN(G1325gat));
  INV_X1    g451(.A(G15gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n461), .A2(new_n455), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n639), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n458), .A2(new_n463), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n639), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n655), .B1(new_n658), .B2(new_n653), .ZN(G1326gat));
  NAND2_X1  g458(.A1(new_n639), .A2(new_n419), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT43), .B(G22gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  INV_X1    g461(.A(new_n611), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n471), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n562), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n531), .A2(new_n665), .A3(new_n634), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n667), .A2(G29gat), .A3(new_n427), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(KEYINPUT45), .Z(new_n669));
  NAND2_X1  g468(.A1(new_n418), .A2(new_n464), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n466), .A2(new_n470), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT44), .B1(new_n672), .B2(new_n611), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT44), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n471), .A2(new_n674), .A3(new_n663), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n666), .ZN(new_n677));
  OAI21_X1  g476(.A(G29gat), .B1(new_n677), .B2(new_n427), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n669), .A2(new_n678), .ZN(G1328gat));
  OAI21_X1  g478(.A(new_n487), .B1(new_n677), .B2(new_n467), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n667), .A2(new_n467), .A3(new_n487), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT46), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n681), .B1(KEYINPUT108), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n680), .B(new_n683), .C1(new_n681), .C2(new_n684), .ZN(G1329gat));
  NAND2_X1  g484(.A1(new_n657), .A2(G43gat), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n667), .B1(new_n455), .B2(new_n461), .ZN(new_n687));
  OAI22_X1  g486(.A1(new_n677), .A2(new_n686), .B1(new_n687), .B2(G43gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g488(.A1(new_n667), .A2(G50gat), .A3(new_n250), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n676), .A2(new_n419), .A3(new_n666), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n691), .B2(G50gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g492(.A1(new_n612), .A2(new_n531), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n672), .A2(new_n634), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n640), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT109), .B(G57gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1332gat));
  AOI21_X1  g497(.A(new_n467), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1333gat));
  INV_X1    g501(.A(G71gat), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n695), .A2(new_n703), .A3(new_n654), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n695), .A2(new_n657), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n704), .B1(new_n705), .B2(new_n703), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g506(.A1(new_n695), .A2(new_n419), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G78gat), .ZN(G1335gat));
  INV_X1    g508(.A(new_n676), .ZN(new_n710));
  INV_X1    g509(.A(new_n531), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n665), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n635), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n710), .A2(new_n427), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT51), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n672), .A2(new_n611), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(new_n713), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n664), .A2(KEYINPUT51), .A3(new_n712), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n640), .A2(new_n568), .A3(new_n634), .ZN(new_n723));
  OAI22_X1  g522(.A1(new_n716), .A2(new_n568), .B1(new_n722), .B2(new_n723), .ZN(G1336gat));
  NAND3_X1  g523(.A1(new_n676), .A2(new_n643), .A3(new_n714), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(G92gat), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n721), .A2(new_n569), .A3(new_n643), .A4(new_n634), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(new_n730), .A3(KEYINPUT52), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT52), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n726), .B(new_n727), .C1(new_n729), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(G1337gat));
  NOR3_X1   g533(.A1(new_n710), .A2(new_n656), .A3(new_n715), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n654), .A2(new_n572), .A3(new_n634), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT111), .Z(new_n737));
  OAI22_X1  g536(.A1(new_n735), .A2(new_n572), .B1(new_n722), .B2(new_n737), .ZN(G1338gat));
  NAND3_X1  g537(.A1(new_n672), .A2(KEYINPUT44), .A3(new_n611), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n674), .B1(new_n471), .B2(new_n663), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n739), .A2(new_n740), .A3(new_n419), .A4(new_n714), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G106gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n419), .A2(new_n573), .A3(new_n634), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n722), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT53), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n573), .B1(new_n741), .B2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n676), .A2(KEYINPUT112), .A3(new_n419), .A4(new_n714), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT113), .ZN(new_n750));
  INV_X1    g549(.A(new_n743), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT53), .B1(new_n721), .B2(new_n751), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n750), .B1(new_n749), .B2(new_n752), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n745), .B1(new_n753), .B2(new_n754), .ZN(G1339gat));
  NAND3_X1  g554(.A1(new_n616), .A2(new_n620), .A3(new_n617), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n622), .A2(KEYINPUT54), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n620), .B1(new_n616), .B2(new_n617), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n631), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n622), .A2(new_n623), .A3(new_n631), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n757), .A2(KEYINPUT55), .A3(new_n760), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n517), .B1(new_n515), .B2(new_n516), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n505), .B1(new_n504), .B2(new_n508), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n523), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n527), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n611), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT114), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n611), .A2(new_n766), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n528), .A2(new_n766), .A3(new_n530), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n770), .A2(new_n634), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n611), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n562), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n694), .A2(new_n635), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n640), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n782), .A2(new_n643), .A3(new_n465), .ZN(new_n783));
  AOI21_X1  g582(.A(G113gat), .B1(new_n783), .B2(new_n711), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n781), .A2(new_n468), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n467), .A2(new_n640), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n711), .A2(G113gat), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n784), .B1(new_n788), .B2(new_n789), .ZN(G1340gat));
  AOI21_X1  g589(.A(G120gat), .B1(new_n783), .B2(new_n634), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n634), .A2(G120gat), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n791), .B1(new_n788), .B2(new_n792), .ZN(G1341gat));
  INV_X1    g592(.A(new_n788), .ZN(new_n794));
  OAI21_X1  g593(.A(G127gat), .B1(new_n794), .B2(new_n562), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n783), .A2(new_n553), .A3(new_n665), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1342gat));
  OAI21_X1  g596(.A(G134gat), .B1(new_n794), .B2(new_n663), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799));
  INV_X1    g598(.A(G134gat), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n799), .A3(new_n800), .A4(new_n611), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n783), .A2(new_n800), .A3(new_n611), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT56), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n798), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT115), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n798), .A2(new_n803), .A3(new_n806), .A4(new_n801), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1343gat));
  NOR2_X1   g607(.A1(new_n657), .A2(new_n786), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n250), .B1(new_n779), .B2(new_n780), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(KEYINPUT57), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812));
  AOI211_X1 g611(.A(new_n812), .B(new_n250), .C1(new_n779), .C2(new_n780), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n711), .B(new_n809), .C1(new_n811), .C2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n814), .A2(G141gat), .B1(new_n815), .B2(KEYINPUT58), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n782), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n781), .A2(KEYINPUT117), .A3(new_n640), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n657), .A2(new_n250), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n467), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n531), .A2(G141gat), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n818), .A2(new_n819), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n816), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(KEYINPUT118), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n821), .B1(new_n782), .B2(new_n817), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n819), .A4(new_n823), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n814), .A2(new_n815), .A3(G141gat), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n830), .A2(new_n831), .A3(new_n816), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n825), .B1(new_n832), .B2(new_n833), .ZN(G1344gat));
  AND2_X1   g633(.A1(new_n827), .A2(new_n819), .ZN(new_n835));
  INV_X1    g634(.A(G148gat), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n835), .A2(new_n836), .A3(new_n634), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n811), .A2(new_n813), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(new_n657), .A3(new_n786), .ZN(new_n839));
  AOI211_X1 g638(.A(KEYINPUT59), .B(new_n836), .C1(new_n839), .C2(new_n634), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n638), .A2(new_n711), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n843));
  OR3_X1    g642(.A1(new_n663), .A2(KEYINPUT121), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT121), .B1(new_n663), .B2(new_n843), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n770), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n778), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n665), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n419), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n812), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n810), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT120), .B1(new_n810), .B2(KEYINPUT57), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n634), .B1(new_n809), .B2(KEYINPUT119), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(KEYINPUT119), .B2(new_n809), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n841), .B1(new_n856), .B2(G148gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n837), .B1(new_n840), .B2(new_n857), .ZN(G1345gat));
  NAND3_X1  g657(.A1(new_n835), .A2(new_n216), .A3(new_n665), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n839), .A2(new_n665), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n859), .B1(new_n861), .B2(new_n216), .ZN(G1346gat));
  AOI21_X1  g661(.A(G162gat), .B1(new_n835), .B2(new_n611), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n663), .A2(new_n217), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n839), .B2(new_n864), .ZN(G1347gat));
  AOI21_X1  g664(.A(new_n640), .B1(new_n779), .B2(new_n780), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n465), .A2(new_n467), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(G169gat), .B1(new_n868), .B2(new_n711), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n643), .A2(new_n427), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT122), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n785), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n531), .A2(new_n316), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(G1348gat));
  INV_X1    g673(.A(new_n872), .ZN(new_n875));
  OAI21_X1  g674(.A(G176gat), .B1(new_n875), .B2(new_n635), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n868), .A2(new_n317), .A3(new_n634), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1349gat));
  NAND3_X1  g677(.A1(new_n785), .A2(new_n665), .A3(new_n871), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n665), .A2(new_n348), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n879), .A2(G183gat), .B1(new_n868), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT123), .B1(new_n881), .B2(KEYINPUT124), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT60), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n881), .B2(KEYINPUT123), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n883), .B1(new_n882), .B2(new_n885), .ZN(G1350gat));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n311), .A3(new_n611), .ZN(new_n887));
  OAI21_X1  g686(.A(G190gat), .B1(new_n875), .B2(new_n663), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(KEYINPUT61), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(KEYINPUT61), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(G1351gat));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n871), .A2(new_n656), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n711), .A2(G197gat), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n853), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n820), .A2(new_n643), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n897), .A2(KEYINPUT125), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(KEYINPUT125), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n898), .A2(new_n866), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(new_n531), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(G197gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n892), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n853), .A2(new_n893), .ZN(new_n904));
  OAI221_X1 g703(.A(KEYINPUT126), .B1(G197gat), .B2(new_n901), .C1(new_n904), .C2(new_n894), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1352gat));
  XNOR2_X1  g705(.A(KEYINPUT127), .B(G204gat), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n900), .A2(new_n635), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT62), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n904), .B2(new_n635), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1353gat));
  OR3_X1    g710(.A1(new_n900), .A2(G211gat), .A3(new_n562), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n853), .A2(new_n665), .A3(new_n893), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n913), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT63), .B1(new_n913), .B2(G211gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(G1354gat));
  OAI21_X1  g715(.A(G218gat), .B1(new_n904), .B2(new_n663), .ZN(new_n917));
  OR2_X1    g716(.A1(new_n663), .A2(G218gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n900), .B2(new_n918), .ZN(G1355gat));
endmodule


