//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977;
  XNOR2_X1  g000(.A(KEYINPUT2), .B(G113), .ZN(new_n187));
  AND2_X1   g001(.A1(KEYINPUT67), .A2(G119), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT67), .A2(G119), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NOR3_X1   g004(.A1(new_n188), .A2(new_n189), .A3(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G116), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n187), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n187), .ZN(new_n195));
  OR2_X1    g009(.A1(KEYINPUT67), .A2(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT67), .A2(G119), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(G116), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n193), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT66), .A2(G134), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT66), .A2(G134), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n203), .B1(new_n206), .B2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G134), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(new_n206), .B2(G137), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n202), .B(new_n207), .C1(new_n211), .C2(new_n203), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(G146), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(KEYINPUT65), .A3(G143), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT1), .B1(new_n214), .B2(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G128), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G143), .B(G146), .ZN(new_n223));
  INV_X1    g037(.A(G128), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n206), .A2(G137), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n208), .A2(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(G131), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n212), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(KEYINPUT0), .A2(G128), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT0), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n224), .A3(KEYINPUT64), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(KEYINPUT0), .B2(G128), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n233), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n219), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n223), .A2(new_n233), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  OR2_X1    g055(.A1(KEYINPUT66), .A2(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(KEYINPUT66), .A2(G134), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(G137), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n203), .B1(new_n244), .B2(new_n209), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT66), .B(G134), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT11), .B1(new_n246), .B2(new_n208), .ZN(new_n247));
  OAI21_X1  g061(.A(G131), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n241), .B1(new_n248), .B2(new_n212), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n232), .A2(new_n249), .A3(KEYINPUT30), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT30), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n238), .A2(new_n219), .B1(new_n233), .B2(new_n223), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n204), .A2(new_n205), .A3(new_n208), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT11), .B1(new_n253), .B2(new_n210), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n202), .B1(new_n254), .B2(new_n207), .ZN(new_n255));
  NOR3_X1   g069(.A1(new_n245), .A2(new_n247), .A3(G131), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n252), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n251), .B1(new_n257), .B2(new_n231), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n201), .B1(new_n250), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n201), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n260), .A3(new_n231), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G237), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT68), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G237), .ZN(new_n266));
  AOI21_X1  g080(.A(G953), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G210), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT26), .B(G101), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n275));
  NOR3_X1   g089(.A1(new_n232), .A2(new_n249), .A3(new_n201), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n260), .B1(new_n257), .B2(new_n231), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT28), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(KEYINPUT70), .B1(new_n276), .B2(KEYINPUT28), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT28), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n261), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n274), .B(new_n275), .C1(new_n273), .C2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  OR2_X1    g099(.A1(new_n283), .A2(new_n273), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n284), .B(new_n285), .C1(new_n275), .C2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G472), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n283), .A2(new_n273), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n259), .A2(new_n272), .A3(new_n261), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT31), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n259), .A2(new_n292), .A3(new_n272), .A4(new_n261), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n289), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G472), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n295), .A3(new_n285), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n296), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT32), .B1(new_n296), .B2(KEYINPUT71), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n288), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(G113), .B(G122), .ZN(new_n300));
  INV_X1    g114(.A(G104), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n300), .B(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n264), .A2(new_n266), .ZN(new_n303));
  INV_X1    g117(.A(G953), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n214), .A2(KEYINPUT83), .ZN(new_n305));
  AND4_X1   g119(.A1(G214), .A2(new_n303), .A3(new_n304), .A4(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT83), .B(G143), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n307), .B1(new_n267), .B2(G214), .ZN(new_n308));
  OAI21_X1  g122(.A(G131), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n265), .A2(G237), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n263), .A2(KEYINPUT68), .ZN(new_n311));
  OAI211_X1 g125(.A(G214), .B(new_n304), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n307), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n267), .A2(G214), .A3(new_n305), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n202), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G125), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n321), .A3(KEYINPUT16), .ZN(new_n322));
  OR3_X1    g136(.A1(new_n320), .A2(KEYINPUT16), .A3(G140), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(G146), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(new_n321), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT19), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n317), .B(new_n326), .C1(G146), .C2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n327), .B(new_n217), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n306), .A2(new_n308), .ZN(new_n331));
  NAND2_X1  g145(.A1(KEYINPUT18), .A2(G131), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT84), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n314), .A2(new_n315), .ZN(new_n335));
  INV_X1    g149(.A(new_n332), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n334), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI211_X1 g151(.A(KEYINPUT84), .B(new_n332), .C1(new_n314), .C2(new_n315), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n333), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n302), .B1(new_n329), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT85), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n336), .B1(new_n306), .B2(new_n308), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(KEYINPUT84), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n335), .A2(new_n334), .A3(new_n336), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT17), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n309), .A2(new_n347), .A3(new_n316), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n322), .A2(new_n323), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n217), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n324), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n202), .B1(new_n314), .B2(new_n315), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(KEYINPUT17), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n346), .A2(new_n333), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n342), .B1(new_n354), .B2(new_n302), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n348), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n339), .A2(new_n356), .A3(new_n342), .A4(new_n302), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n341), .B1(new_n355), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(G475), .A2(G902), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n339), .A2(new_n356), .A3(new_n302), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT85), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n340), .B1(new_n364), .B2(new_n357), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT86), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n361), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT20), .ZN(new_n368));
  INV_X1    g182(.A(new_n362), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(KEYINPUT20), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n359), .A2(KEYINPUT87), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT87), .ZN(new_n372));
  INV_X1    g186(.A(new_n370), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n372), .B1(new_n365), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n368), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n354), .ZN(new_n378));
  INV_X1    g192(.A(new_n302), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n364), .A2(new_n357), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(G475), .B1(new_n380), .B2(G902), .ZN(new_n381));
  XOR2_X1   g195(.A(G128), .B(G143), .Z(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(new_n246), .ZN(new_n383));
  XNOR2_X1  g197(.A(G116), .B(G122), .ZN(new_n384));
  INV_X1    g198(.A(G107), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n190), .A2(KEYINPUT14), .A3(G122), .ZN(new_n387));
  INV_X1    g201(.A(new_n384), .ZN(new_n388));
  OAI211_X1 g202(.A(G107), .B(new_n387), .C1(new_n388), .C2(KEYINPUT14), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n383), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n384), .B(new_n385), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT13), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n214), .A3(G128), .ZN(new_n393));
  OAI211_X1 g207(.A(G134), .B(new_n393), .C1(new_n382), .C2(new_n392), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n391), .B(new_n394), .C1(new_n246), .C2(new_n382), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT9), .B(G234), .ZN(new_n396));
  INV_X1    g210(.A(G217), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n396), .A2(new_n397), .A3(G953), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n390), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n390), .B2(new_n395), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT15), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G478), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n285), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n285), .B1(new_n399), .B2(new_n400), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n402), .A3(G478), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(G234), .A2(G237), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(G952), .A3(new_n304), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT88), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(G902), .A3(G953), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT21), .B(G898), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n407), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n377), .A2(new_n381), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n397), .B1(G234), .B2(new_n285), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT24), .B(G110), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n188), .A2(new_n189), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(G128), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT72), .B1(new_n192), .B2(G128), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT72), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n424), .A2(new_n224), .A3(G119), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n422), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT23), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n421), .B2(G128), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n224), .A2(KEYINPUT23), .A3(G119), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n428), .A2(new_n422), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(G110), .ZN(new_n431));
  OAI221_X1 g245(.A(new_n351), .B1(new_n420), .B2(new_n426), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n327), .A2(G146), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n428), .A2(new_n431), .A3(new_n422), .A4(new_n429), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n188), .A2(new_n189), .A3(new_n224), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n423), .A2(new_n425), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n420), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n433), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n438), .A2(new_n326), .A3(KEYINPUT74), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT74), .B1(new_n438), .B2(new_n326), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n432), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT75), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT75), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n443), .B(new_n432), .C1(new_n439), .C2(new_n440), .ZN(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT22), .B(G137), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n304), .A2(G221), .A3(G234), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n445), .B(new_n446), .Z(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n442), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n441), .A2(KEYINPUT75), .A3(new_n447), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT25), .B1(new_n451), .B2(new_n285), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT25), .ZN(new_n453));
  AOI211_X1 g267(.A(new_n453), .B(G902), .C1(new_n449), .C2(new_n450), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n419), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n419), .A2(G902), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT3), .B1(new_n301), .B2(G107), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT3), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(new_n385), .A3(G104), .ZN(new_n462));
  INV_X1    g276(.A(G101), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n301), .A2(G107), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n460), .A2(new_n462), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n301), .A2(G107), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n385), .A2(G104), .ZN(new_n467));
  OAI21_X1  g281(.A(G101), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n217), .A2(G143), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n220), .A2(G128), .B1(new_n470), .B2(new_n216), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT78), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n226), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n224), .B1(new_n470), .B2(KEYINPUT1), .ZN(new_n474));
  NOR3_X1   g288(.A1(new_n474), .A2(new_n223), .A3(KEYINPUT78), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n469), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT10), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n255), .A2(new_n256), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n460), .A2(new_n462), .A3(new_n464), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G101), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(KEYINPUT4), .A3(new_n465), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT4), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(new_n483), .A3(G101), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n252), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n227), .A2(new_n469), .A3(KEYINPUT10), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n478), .A2(new_n479), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n465), .A2(new_n468), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n222), .A3(new_n226), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n476), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n248), .A2(new_n212), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(KEYINPUT12), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT12), .B1(new_n490), .B2(new_n491), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G110), .B(G140), .ZN(new_n496));
  INV_X1    g310(.A(G227), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n497), .A2(G953), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n496), .B(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n499), .B(KEYINPUT77), .Z(new_n500));
  INV_X1    g314(.A(new_n499), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n487), .A2(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n225), .A2(new_n470), .A3(new_n216), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT1), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(G143), .B2(new_n217), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n214), .A2(G146), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n217), .A2(G143), .ZN(new_n507));
  OAI22_X1  g321(.A1(new_n505), .A2(new_n224), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n503), .B1(new_n508), .B2(KEYINPUT78), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n471), .A2(new_n472), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n488), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n485), .B(new_n486), .C1(new_n511), .C2(KEYINPUT10), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n491), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n495), .A2(new_n500), .B1(new_n502), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(G469), .B1(new_n514), .B2(G902), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT79), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(KEYINPUT79), .B(G469), .C1(new_n514), .C2(G902), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n487), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n499), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n487), .B(new_n501), .C1(new_n493), .C2(new_n494), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(G469), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n523), .A3(new_n285), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n517), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(G214), .B1(G237), .B2(G902), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n201), .A2(new_n482), .A3(new_n484), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n198), .A2(KEYINPUT5), .A3(new_n199), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT5), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n196), .A2(new_n531), .A3(G116), .A4(new_n197), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G113), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n469), .B(new_n200), .C1(new_n530), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(G110), .B(G122), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n528), .A2(new_n534), .A3(new_n536), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(KEYINPUT6), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT6), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n535), .A2(new_n541), .A3(new_n537), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n222), .A2(new_n320), .A3(new_n226), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n543), .B1(new_n252), .B2(new_n320), .ZN(new_n544));
  INV_X1    g358(.A(G224), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G953), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n544), .B(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n540), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT7), .B1(new_n545), .B2(G953), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n543), .B(new_n550), .C1(new_n320), .C2(new_n252), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n539), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n200), .B(new_n488), .C1(new_n530), .C2(new_n533), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n536), .B(KEYINPUT8), .ZN(new_n554));
  INV_X1    g368(.A(new_n200), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT80), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n533), .B1(new_n556), .B2(new_n529), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n198), .A2(KEYINPUT80), .A3(KEYINPUT5), .A4(new_n199), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n555), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n553), .B(new_n554), .C1(new_n559), .C2(new_n488), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT81), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n222), .A2(new_n561), .A3(new_n320), .A4(new_n226), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n562), .A2(new_n549), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n543), .B(KEYINPUT81), .C1(new_n320), .C2(new_n252), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT82), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT82), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n563), .A2(new_n564), .A3(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n552), .A2(new_n560), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n548), .A2(new_n569), .A3(new_n285), .ZN(new_n570));
  OAI21_X1  g384(.A(G210), .B1(G237), .B2(G902), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n548), .A2(new_n569), .A3(new_n285), .A4(new_n571), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n527), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G221), .ZN(new_n576));
  INV_X1    g390(.A(new_n396), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n577), .B2(new_n285), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n578), .B(KEYINPUT76), .Z(new_n579));
  NAND3_X1  g393(.A1(new_n525), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n299), .A2(new_n418), .A3(new_n459), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  INV_X1    g397(.A(new_n415), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n455), .A2(new_n457), .A3(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(new_n580), .ZN(new_n586));
  INV_X1    g400(.A(new_n381), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n368), .B2(new_n376), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n401), .B(KEYINPUT33), .Z(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G478), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n405), .A2(G478), .ZN(new_n591));
  NAND2_X1  g405(.A1(G478), .A2(G902), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n294), .A2(new_n285), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G472), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(KEYINPUT89), .A3(new_n296), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT89), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n595), .A2(new_n598), .A3(G472), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n586), .A2(new_n594), .A3(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT34), .B(G104), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT90), .B(KEYINPUT91), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  INV_X1    g419(.A(KEYINPUT20), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n361), .A2(new_n366), .A3(new_n606), .A4(new_n362), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n368), .A2(KEYINPUT92), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT92), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n367), .A2(new_n609), .A3(KEYINPUT20), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n381), .A2(KEYINPUT93), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT93), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n612), .B(G475), .C1(new_n380), .C2(G902), .ZN(new_n613));
  AND3_X1   g427(.A1(new_n611), .A2(new_n407), .A3(new_n613), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n608), .A2(new_n610), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n586), .A3(new_n600), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT35), .B(G107), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  NOR2_X1   g432(.A1(new_n448), .A2(KEYINPUT36), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n441), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n456), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n455), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n418), .A2(new_n600), .A3(new_n581), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT37), .B(G110), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT94), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n623), .B(new_n625), .ZN(G12));
  INV_X1    g440(.A(new_n410), .ZN(new_n627));
  INV_X1    g441(.A(G900), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n627), .B1(new_n628), .B2(new_n412), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT95), .Z(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n615), .A2(KEYINPUT96), .A3(new_n575), .A4(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n608), .A2(new_n610), .A3(new_n614), .A4(new_n631), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n566), .A2(new_n560), .A3(new_n568), .ZN(new_n635));
  AOI21_X1  g449(.A(G902), .B1(new_n635), .B2(new_n552), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n571), .B1(new_n636), .B2(new_n548), .ZN(new_n637));
  INV_X1    g451(.A(new_n574), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n526), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n633), .B1(new_n634), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n622), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n296), .A2(KEYINPUT71), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT32), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n296), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n641), .B1(new_n646), .B2(new_n288), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n525), .A2(new_n579), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n632), .A2(new_n640), .A3(new_n647), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G128), .ZN(G30));
  NAND2_X1  g465(.A1(new_n377), .A2(new_n381), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n630), .B(KEYINPUT39), .Z(new_n653));
  NAND2_X1  g467(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT40), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n637), .A2(new_n638), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n658), .A2(new_n622), .A3(new_n527), .ZN(new_n659));
  AND4_X1   g473(.A1(new_n652), .A2(new_n655), .A3(new_n407), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n262), .A2(new_n272), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n276), .A2(new_n277), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n285), .B1(new_n663), .B2(new_n272), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n646), .A2(new_n665), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n660), .B(new_n666), .C1(KEYINPUT40), .C2(new_n654), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT98), .B(G143), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G45));
  INV_X1    g483(.A(new_n593), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n375), .B1(KEYINPUT20), .B2(new_n367), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n670), .B(new_n631), .C1(new_n671), .C2(new_n587), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n580), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n647), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G146), .ZN(G48));
  INV_X1    g489(.A(new_n299), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n676), .A2(new_n458), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n523), .B1(new_n522), .B2(new_n285), .ZN(new_n678));
  AOI211_X1 g492(.A(G469), .B(G902), .C1(new_n520), .C2(new_n521), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n578), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n680), .A2(new_n575), .A3(new_n681), .A4(new_n584), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n588), .A2(new_n682), .A3(new_n593), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  INV_X1    g500(.A(new_n494), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(new_n492), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n688), .A2(new_n502), .B1(new_n519), .B2(new_n499), .ZN(new_n689));
  OAI21_X1  g503(.A(G469), .B1(new_n689), .B2(G902), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n681), .A3(new_n524), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n639), .A2(new_n691), .A3(new_n415), .ZN(new_n692));
  AND4_X1   g506(.A1(new_n610), .A2(new_n608), .A3(new_n692), .A4(new_n614), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n677), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  INV_X1    g509(.A(KEYINPUT99), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n639), .B2(new_n691), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n680), .A2(new_n575), .A3(KEYINPUT99), .A4(new_n681), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n417), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n647), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  INV_X1    g516(.A(new_n407), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n588), .A2(new_n682), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n595), .A2(KEYINPUT100), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G472), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n595), .A2(KEYINPUT100), .A3(new_n295), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(KEYINPUT101), .B1(new_n708), .B2(new_n459), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n295), .B1(new_n595), .B2(KEYINPUT100), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT100), .ZN(new_n711));
  AOI211_X1 g525(.A(new_n711), .B(G472), .C1(new_n294), .C2(new_n285), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT101), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n713), .A2(new_n714), .A3(new_n458), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n704), .B1(new_n709), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT102), .B(G122), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G24));
  NOR2_X1   g532(.A1(new_n672), .A2(new_n699), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n706), .A2(new_n707), .B1(new_n455), .B2(new_n621), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  INV_X1    g536(.A(new_n672), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n578), .B1(new_n515), .B2(new_n524), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n637), .A2(new_n638), .A3(new_n527), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n723), .A2(new_n299), .A3(new_n459), .A4(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n728), .A2(KEYINPUT103), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT42), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n730), .B1(new_n728), .B2(KEYINPUT103), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n296), .A2(new_n643), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n288), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n296), .A2(new_n643), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n459), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n723), .A2(KEYINPUT42), .A3(new_n727), .ZN(new_n736));
  OAI22_X1  g550(.A1(new_n729), .A2(new_n731), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G131), .ZN(G33));
  INV_X1    g552(.A(new_n634), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n739), .A2(new_n299), .A3(new_n459), .A4(new_n727), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT104), .B(G134), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G36));
  NOR3_X1   g556(.A1(new_n652), .A2(KEYINPUT43), .A3(new_n593), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n593), .B1(new_n652), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n744), .B2(new_n652), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n743), .B1(new_n746), .B2(KEYINPUT43), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n600), .A2(new_n641), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT44), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n725), .ZN(new_n750));
  OAI21_X1  g564(.A(G469), .B1(new_n514), .B2(KEYINPUT45), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT105), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n752), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n514), .A2(KEYINPUT45), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(G469), .A2(G902), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT46), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n679), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n757), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n681), .A3(new_n653), .ZN(new_n762));
  NOR3_X1   g576(.A1(new_n749), .A2(new_n750), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n747), .A2(KEYINPUT44), .A3(new_n748), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT107), .B(G137), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G39));
  NAND3_X1  g581(.A1(new_n723), .A2(new_n458), .A3(new_n725), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(new_n299), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n578), .B1(new_n759), .B2(new_n760), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n770), .A2(KEYINPUT47), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(KEYINPUT47), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g587(.A(KEYINPUT108), .B(G140), .Z(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G42));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n647), .A2(new_n673), .B1(new_n719), .B2(new_n720), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n588), .A2(new_n639), .A3(new_n703), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n630), .B(KEYINPUT113), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n724), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n666), .A2(new_n641), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n650), .A2(new_n777), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n650), .A2(new_n777), .A3(KEYINPUT52), .A4(new_n781), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n608), .A2(new_n610), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n404), .A2(KEYINPUT111), .A3(new_n406), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT111), .B1(new_n404), .B2(new_n406), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n788), .A2(new_n789), .A3(new_n630), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n725), .A2(new_n611), .A3(new_n613), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n648), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n299), .A2(new_n787), .A3(new_n622), .A4(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n723), .A2(new_n720), .A3(new_n727), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n740), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT112), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n740), .A2(new_n793), .A3(KEYINPUT112), .A4(new_n794), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n299), .B(new_n459), .C1(new_n693), .C2(new_n683), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n716), .A2(new_n701), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n788), .A2(new_n789), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n671), .A2(new_n587), .A3(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n586), .B(new_n600), .C1(new_n594), .C2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n582), .A3(new_n623), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n799), .A2(new_n806), .A3(new_n737), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n776), .B1(new_n786), .B2(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n804), .A2(new_n582), .A3(new_n623), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n714), .B1(new_n713), .B2(new_n458), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n708), .A2(new_n459), .A3(KEYINPUT101), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n812), .A2(new_n704), .B1(new_n647), .B2(new_n700), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n809), .A2(new_n813), .A3(new_n800), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n797), .B2(new_n798), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n784), .A2(new_n785), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n815), .A2(new_n816), .A3(KEYINPUT53), .A4(new_n737), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n808), .A2(KEYINPUT115), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n807), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n820), .A3(KEYINPUT53), .A4(new_n816), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n823), .B1(new_n808), .B2(new_n817), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(KEYINPUT114), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n829), .A2(KEYINPUT51), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n410), .B1(new_n810), .B2(new_n811), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n747), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n658), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n834), .A2(new_n526), .A3(new_n691), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XOR2_X1   g650(.A(new_n836), .B(KEYINPUT50), .Z(new_n837));
  NOR3_X1   g651(.A1(new_n750), .A2(new_n410), .A3(new_n691), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n747), .A2(new_n720), .A3(new_n838), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n646), .A2(new_n459), .A3(new_n665), .A4(new_n838), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n588), .A3(new_n593), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n680), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n771), .B(new_n772), .C1(new_n579), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n832), .A2(new_n750), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n830), .B1(new_n837), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n837), .A2(new_n830), .A3(new_n846), .ZN(new_n848));
  INV_X1    g662(.A(G952), .ZN(new_n849));
  OAI21_X1  g663(.A(KEYINPUT117), .B1(new_n849), .B2(G953), .ZN(new_n850));
  OAI221_X1 g664(.A(new_n850), .B1(new_n829), .B2(KEYINPUT51), .C1(KEYINPUT117), .C2(G953), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n840), .B2(new_n594), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(new_n832), .B2(new_n699), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n747), .A2(new_n838), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(new_n735), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n855), .A2(KEYINPUT48), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(KEYINPUT48), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n848), .A2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n828), .A2(new_n847), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(G952), .A2(G953), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n459), .A2(new_n526), .A3(new_n579), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT109), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n746), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(KEYINPUT110), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(KEYINPUT110), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n680), .B(KEYINPUT49), .Z(new_n867));
  NOR3_X1   g681(.A1(new_n666), .A2(new_n834), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n860), .A2(new_n861), .B1(new_n865), .B2(new_n869), .ZN(G75));
  INV_X1    g684(.A(new_n822), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(G210), .A3(G902), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT56), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n540), .A2(new_n542), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT118), .Z(new_n875));
  XOR2_X1   g689(.A(new_n547), .B(KEYINPUT55), .Z(new_n876));
  XNOR2_X1  g690(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n872), .A2(new_n873), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n877), .B1(new_n872), .B2(new_n873), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n304), .A2(G952), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G51));
  XOR2_X1   g695(.A(new_n757), .B(KEYINPUT57), .Z(new_n882));
  INV_X1    g696(.A(new_n824), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n822), .A2(new_n823), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n522), .ZN(new_n886));
  OR3_X1    g700(.A1(new_n822), .A2(new_n285), .A3(new_n756), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n880), .B1(new_n886), .B2(new_n887), .ZN(G54));
  NAND4_X1  g702(.A1(new_n871), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n361), .A2(new_n366), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n889), .A2(KEYINPUT119), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n880), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n889), .B2(new_n890), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT119), .B1(new_n889), .B2(new_n890), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n891), .A2(new_n893), .A3(new_n894), .ZN(G60));
  INV_X1    g709(.A(new_n589), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n592), .B(KEYINPUT59), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n896), .B(new_n897), .C1(new_n883), .C2(new_n884), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n892), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n896), .B1(new_n828), .B2(new_n897), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(G63));
  NAND2_X1  g715(.A1(G217), .A2(G902), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT60), .Z(new_n903));
  NAND3_X1  g717(.A1(new_n818), .A2(new_n821), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n451), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n818), .A2(new_n620), .A3(new_n821), .A4(new_n903), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n906), .A2(KEYINPUT61), .A3(new_n892), .A4(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n880), .B1(new_n904), .B2(new_n905), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(KEYINPUT121), .A3(KEYINPUT61), .A4(new_n907), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AOI211_X1 g727(.A(KEYINPUT120), .B(KEYINPUT61), .C1(new_n911), .C2(new_n907), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n911), .A2(new_n907), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT61), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n913), .B1(new_n914), .B2(new_n918), .ZN(G66));
  OAI21_X1  g733(.A(G953), .B1(new_n413), .B2(new_n545), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n806), .B2(G953), .ZN(new_n921));
  INV_X1    g735(.A(new_n875), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(G898), .B2(new_n304), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT122), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n921), .B(new_n924), .ZN(G69));
  OAI21_X1  g739(.A(G953), .B1(new_n497), .B2(new_n628), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n250), .A2(new_n258), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(new_n328), .Z(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n773), .B1(new_n763), .B2(new_n764), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n594), .A2(new_n803), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n933), .A2(new_n654), .A3(new_n750), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n932), .B1(new_n677), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n650), .A2(new_n777), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT123), .Z(new_n937));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n937), .B(new_n667), .C1(KEYINPUT124), .C2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n667), .ZN(new_n940));
  XOR2_X1   g754(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n935), .A2(new_n939), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n930), .B1(new_n943), .B2(new_n304), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n778), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n946), .A2(new_n735), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n770), .A2(new_n947), .A3(new_n653), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n737), .A2(new_n740), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n931), .A2(new_n937), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n304), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n304), .A2(G900), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT125), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n929), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n927), .B1(new_n945), .B2(new_n956), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n944), .A2(new_n955), .A3(new_n926), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n957), .A2(new_n958), .ZN(G72));
  NAND4_X1  g773(.A1(new_n935), .A2(new_n806), .A3(new_n939), .A4(new_n942), .ZN(new_n960));
  NAND2_X1  g774(.A1(G472), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT63), .Z(new_n962));
  NAND2_X1  g776(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n662), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n808), .A2(new_n817), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n274), .A2(new_n290), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n962), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT126), .Z(new_n968));
  NAND2_X1  g782(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n962), .B1(new_n951), .B2(new_n814), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n262), .A2(new_n272), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n880), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n964), .A2(KEYINPUT127), .A3(new_n969), .A4(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT127), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n661), .B1(new_n960), .B2(new_n962), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n972), .A2(new_n969), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n973), .A2(new_n977), .ZN(G57));
endmodule


