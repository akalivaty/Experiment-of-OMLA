

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U554 ( .A1(n984), .A2(G138), .ZN(n522) );
  NOR2_X1 U555 ( .A1(n530), .A2(n529), .ZN(G164) );
  NOR2_X1 U556 ( .A1(n538), .A2(n537), .ZN(G160) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n699) );
  INV_X1 U558 ( .A(KEYINPUT93), .ZN(n717) );
  XNOR2_X1 U559 ( .A(n718), .B(n717), .ZN(n724) );
  NOR2_X1 U560 ( .A1(G164), .A2(G1384), .ZN(n766) );
  NOR2_X1 U561 ( .A1(n764), .A2(n763), .ZN(n765) );
  INV_X1 U562 ( .A(KEYINPUT17), .ZN(n520) );
  NOR2_X1 U563 ( .A1(G543), .A2(G651), .ZN(n645) );
  NOR2_X2 U564 ( .A1(G2105), .A2(n526), .ZN(n983) );
  NOR2_X1 U565 ( .A1(n633), .A2(G651), .ZN(n639) );
  INV_X1 U566 ( .A(KEYINPUT83), .ZN(n523) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  XNOR2_X2 U568 ( .A(n521), .B(n520), .ZN(n984) );
  XNOR2_X1 U569 ( .A(n523), .B(n522), .ZN(n525) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n979) );
  NAND2_X1 U571 ( .A1(n979), .A2(G114), .ZN(n524) );
  NAND2_X1 U572 ( .A1(n525), .A2(n524), .ZN(n530) );
  INV_X1 U573 ( .A(G2104), .ZN(n526) );
  NAND2_X1 U574 ( .A1(G102), .A2(n983), .ZN(n528) );
  AND2_X1 U575 ( .A1(n526), .A2(G2105), .ZN(n980) );
  NAND2_X1 U576 ( .A1(G126), .A2(n980), .ZN(n527) );
  NAND2_X1 U577 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U578 ( .A1(G101), .A2(n983), .ZN(n531) );
  XOR2_X1 U579 ( .A(KEYINPUT23), .B(n531), .Z(n534) );
  NAND2_X1 U580 ( .A1(G113), .A2(n979), .ZN(n532) );
  XOR2_X1 U581 ( .A(KEYINPUT65), .B(n532), .Z(n533) );
  NAND2_X1 U582 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U583 ( .A1(G137), .A2(n984), .ZN(n536) );
  NAND2_X1 U584 ( .A1(G125), .A2(n980), .ZN(n535) );
  NAND2_X1 U585 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  NAND2_X1 U587 ( .A1(G52), .A2(n639), .ZN(n541) );
  XOR2_X1 U588 ( .A(G651), .B(KEYINPUT66), .Z(n543) );
  NOR2_X1 U589 ( .A1(G543), .A2(n543), .ZN(n539) );
  XOR2_X2 U590 ( .A(KEYINPUT1), .B(n539), .Z(n641) );
  NAND2_X1 U591 ( .A1(G64), .A2(n641), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U593 ( .A(KEYINPUT70), .B(n542), .ZN(n549) );
  NAND2_X1 U594 ( .A1(G90), .A2(n645), .ZN(n546) );
  OR2_X1 U595 ( .A1(n633), .A2(n543), .ZN(n544) );
  XNOR2_X1 U596 ( .A(KEYINPUT67), .B(n544), .ZN(n646) );
  NAND2_X1 U597 ( .A1(G77), .A2(n646), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U599 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U600 ( .A1(n549), .A2(n548), .ZN(G171) );
  AND2_X1 U601 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U602 ( .A(G132), .ZN(G219) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  INV_X1 U604 ( .A(G57), .ZN(G237) );
  NAND2_X1 U605 ( .A1(n639), .A2(G50), .ZN(n556) );
  NAND2_X1 U606 ( .A1(G62), .A2(n641), .ZN(n551) );
  NAND2_X1 U607 ( .A1(G75), .A2(n646), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n551), .A2(n550), .ZN(n554) );
  NAND2_X1 U609 ( .A1(G88), .A2(n645), .ZN(n552) );
  XNOR2_X1 U610 ( .A(KEYINPUT79), .B(n552), .ZN(n553) );
  NOR2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U613 ( .A(KEYINPUT80), .B(n557), .Z(G166) );
  INV_X1 U614 ( .A(G166), .ZN(G303) );
  NAND2_X1 U615 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U616 ( .A(n558), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U617 ( .A(G223), .ZN(n819) );
  NAND2_X1 U618 ( .A1(n819), .A2(G567), .ZN(n559) );
  XOR2_X1 U619 ( .A(KEYINPUT11), .B(n559), .Z(G234) );
  NAND2_X1 U620 ( .A1(G56), .A2(n641), .ZN(n560) );
  XOR2_X1 U621 ( .A(KEYINPUT14), .B(n560), .Z(n566) );
  NAND2_X1 U622 ( .A1(n645), .A2(G81), .ZN(n561) );
  XNOR2_X1 U623 ( .A(n561), .B(KEYINPUT12), .ZN(n563) );
  NAND2_X1 U624 ( .A1(G68), .A2(n646), .ZN(n562) );
  NAND2_X1 U625 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT13), .B(n564), .Z(n565) );
  NOR2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U628 ( .A1(n639), .A2(G43), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n681) );
  INV_X1 U630 ( .A(G860), .ZN(n599) );
  OR2_X1 U631 ( .A1(n681), .A2(n599), .ZN(G153) );
  INV_X1 U632 ( .A(G171), .ZN(G301) );
  NAND2_X1 U633 ( .A1(G868), .A2(G301), .ZN(n577) );
  NAND2_X1 U634 ( .A1(G54), .A2(n639), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G79), .A2(n646), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U637 ( .A1(G92), .A2(n645), .ZN(n572) );
  NAND2_X1 U638 ( .A1(G66), .A2(n641), .ZN(n571) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT15), .ZN(n904) );
  INV_X1 U642 ( .A(G868), .ZN(n659) );
  NAND2_X1 U643 ( .A1(n904), .A2(n659), .ZN(n576) );
  NAND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(G284) );
  NAND2_X1 U645 ( .A1(n645), .A2(G89), .ZN(n578) );
  XNOR2_X1 U646 ( .A(n578), .B(KEYINPUT4), .ZN(n580) );
  NAND2_X1 U647 ( .A1(G76), .A2(n646), .ZN(n579) );
  NAND2_X1 U648 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U649 ( .A(KEYINPUT5), .B(n581), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n641), .A2(G63), .ZN(n582) );
  XOR2_X1 U651 ( .A(KEYINPUT73), .B(n582), .Z(n584) );
  NAND2_X1 U652 ( .A1(n639), .A2(G51), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U654 ( .A(KEYINPUT6), .B(n585), .Z(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U656 ( .A(KEYINPUT7), .B(n588), .ZN(G168) );
  XOR2_X1 U657 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U658 ( .A1(n639), .A2(G53), .ZN(n589) );
  XOR2_X1 U659 ( .A(KEYINPUT71), .B(n589), .Z(n591) );
  NAND2_X1 U660 ( .A1(n641), .A2(G65), .ZN(n590) );
  NAND2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U662 ( .A(KEYINPUT72), .B(n592), .Z(n596) );
  NAND2_X1 U663 ( .A1(G91), .A2(n645), .ZN(n594) );
  NAND2_X1 U664 ( .A1(G78), .A2(n646), .ZN(n593) );
  AND2_X1 U665 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n596), .A2(n595), .ZN(G299) );
  NOR2_X1 U667 ( .A1(G286), .A2(n659), .ZN(n598) );
  NOR2_X1 U668 ( .A1(G868), .A2(G299), .ZN(n597) );
  NOR2_X1 U669 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n599), .A2(G559), .ZN(n600) );
  INV_X1 U671 ( .A(n904), .ZN(n1008) );
  NAND2_X1 U672 ( .A1(n600), .A2(n1008), .ZN(n601) );
  XNOR2_X1 U673 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U674 ( .A1(n904), .A2(n659), .ZN(n602) );
  XOR2_X1 U675 ( .A(KEYINPUT74), .B(n602), .Z(n603) );
  NOR2_X1 U676 ( .A1(G559), .A2(n603), .ZN(n605) );
  NOR2_X1 U677 ( .A1(G868), .A2(n681), .ZN(n604) );
  NOR2_X1 U678 ( .A1(n605), .A2(n604), .ZN(G282) );
  NAND2_X1 U679 ( .A1(G111), .A2(n979), .ZN(n607) );
  NAND2_X1 U680 ( .A1(G135), .A2(n984), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n980), .A2(G123), .ZN(n608) );
  XOR2_X1 U683 ( .A(KEYINPUT18), .B(n608), .Z(n609) );
  NOR2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n983), .A2(G99), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n996) );
  XOR2_X1 U687 ( .A(n996), .B(G2096), .Z(n614) );
  XNOR2_X1 U688 ( .A(G2100), .B(KEYINPUT75), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(G156) );
  XNOR2_X1 U690 ( .A(n681), .B(KEYINPUT76), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n1008), .A2(G559), .ZN(n615) );
  XNOR2_X1 U692 ( .A(n616), .B(n615), .ZN(n657) );
  NOR2_X1 U693 ( .A1(G860), .A2(n657), .ZN(n624) );
  NAND2_X1 U694 ( .A1(G93), .A2(n645), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G80), .A2(n646), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n623) );
  NAND2_X1 U697 ( .A1(G55), .A2(n639), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G67), .A2(n641), .ZN(n619) );
  NAND2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U700 ( .A(KEYINPUT77), .B(n621), .Z(n622) );
  OR2_X1 U701 ( .A1(n623), .A2(n622), .ZN(n660) );
  XOR2_X1 U702 ( .A(n624), .B(n660), .Z(G145) );
  NAND2_X1 U703 ( .A1(n645), .A2(G86), .ZN(n631) );
  NAND2_X1 U704 ( .A1(G48), .A2(n639), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G61), .A2(n641), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G73), .A2(n646), .ZN(n627) );
  XOR2_X1 U708 ( .A(KEYINPUT2), .B(n627), .Z(n628) );
  NOR2_X1 U709 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U711 ( .A(n632), .B(KEYINPUT78), .ZN(G305) );
  NAND2_X1 U712 ( .A1(G74), .A2(G651), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G87), .A2(n633), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U715 ( .A1(n641), .A2(n636), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(G49), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(G288) );
  NAND2_X1 U718 ( .A1(n639), .A2(G47), .ZN(n640) );
  XNOR2_X1 U719 ( .A(n640), .B(KEYINPUT68), .ZN(n643) );
  NAND2_X1 U720 ( .A1(G60), .A2(n641), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U722 ( .A(KEYINPUT69), .B(n644), .ZN(n650) );
  NAND2_X1 U723 ( .A1(G85), .A2(n645), .ZN(n648) );
  NAND2_X1 U724 ( .A1(G72), .A2(n646), .ZN(n647) );
  AND2_X1 U725 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(G290) );
  INV_X1 U727 ( .A(G299), .ZN(n891) );
  XNOR2_X1 U728 ( .A(G305), .B(n891), .ZN(n656) );
  XNOR2_X1 U729 ( .A(KEYINPUT19), .B(G166), .ZN(n651) );
  XNOR2_X1 U730 ( .A(n651), .B(G288), .ZN(n652) );
  XNOR2_X1 U731 ( .A(KEYINPUT81), .B(n652), .ZN(n654) );
  XOR2_X1 U732 ( .A(G290), .B(n660), .Z(n653) );
  XNOR2_X1 U733 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n656), .B(n655), .ZN(n1007) );
  XOR2_X1 U735 ( .A(n1007), .B(n657), .Z(n658) );
  NOR2_X1 U736 ( .A1(n659), .A2(n658), .ZN(n662) );
  NOR2_X1 U737 ( .A1(G868), .A2(n660), .ZN(n661) );
  NOR2_X1 U738 ( .A1(n662), .A2(n661), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2078), .A2(G2084), .ZN(n663) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n663), .Z(n664) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n665), .ZN(n666) );
  NAND2_X1 U743 ( .A1(n666), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U745 ( .A1(G108), .A2(G120), .ZN(n667) );
  NOR2_X1 U746 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U747 ( .A1(G69), .A2(n668), .ZN(n954) );
  NAND2_X1 U748 ( .A1(G567), .A2(n954), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n669), .B(KEYINPUT82), .ZN(n674) );
  NOR2_X1 U750 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U751 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U752 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U753 ( .A1(G96), .A2(n672), .ZN(n955) );
  NAND2_X1 U754 ( .A1(G2106), .A2(n955), .ZN(n673) );
  NAND2_X1 U755 ( .A1(n674), .A2(n673), .ZN(n956) );
  NAND2_X1 U756 ( .A1(G661), .A2(G483), .ZN(n675) );
  NOR2_X1 U757 ( .A1(n956), .A2(n675), .ZN(n823) );
  NAND2_X1 U758 ( .A1(n823), .A2(G36), .ZN(G176) );
  NAND2_X1 U759 ( .A1(G160), .A2(G40), .ZN(n767) );
  INV_X1 U760 ( .A(n767), .ZN(n677) );
  AND2_X1 U761 ( .A1(n677), .A2(n766), .ZN(n701) );
  NAND2_X1 U762 ( .A1(n701), .A2(G1996), .ZN(n676) );
  XNOR2_X1 U763 ( .A(n676), .B(KEYINPUT26), .ZN(n679) );
  NAND2_X1 U764 ( .A1(n677), .A2(n766), .ZN(n719) );
  NAND2_X1 U765 ( .A1(n719), .A2(G1341), .ZN(n678) );
  NAND2_X1 U766 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U767 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U768 ( .A(n682), .B(KEYINPUT64), .Z(n687) );
  OR2_X1 U769 ( .A1(n687), .A2(n904), .ZN(n686) );
  NOR2_X1 U770 ( .A1(G2067), .A2(n719), .ZN(n684) );
  NOR2_X1 U771 ( .A1(n701), .A2(G1348), .ZN(n683) );
  NOR2_X1 U772 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U773 ( .A1(n686), .A2(n685), .ZN(n689) );
  NAND2_X1 U774 ( .A1(n687), .A2(n904), .ZN(n688) );
  NAND2_X1 U775 ( .A1(n689), .A2(n688), .ZN(n694) );
  NAND2_X1 U776 ( .A1(n701), .A2(G2072), .ZN(n690) );
  XNOR2_X1 U777 ( .A(n690), .B(KEYINPUT27), .ZN(n692) );
  AND2_X1 U778 ( .A1(G1956), .A2(n719), .ZN(n691) );
  NOR2_X1 U779 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U780 ( .A1(n891), .A2(n695), .ZN(n693) );
  NAND2_X1 U781 ( .A1(n694), .A2(n693), .ZN(n698) );
  NOR2_X1 U782 ( .A1(n891), .A2(n695), .ZN(n696) );
  XOR2_X1 U783 ( .A(n696), .B(KEYINPUT28), .Z(n697) );
  NAND2_X1 U784 ( .A1(n698), .A2(n697), .ZN(n700) );
  XNOR2_X1 U785 ( .A(n700), .B(n699), .ZN(n706) );
  XOR2_X1 U786 ( .A(G2078), .B(KEYINPUT25), .Z(n837) );
  NOR2_X1 U787 ( .A1(n837), .A2(n719), .ZN(n703) );
  NOR2_X1 U788 ( .A1(n701), .A2(G1961), .ZN(n702) );
  NOR2_X1 U789 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U790 ( .A(KEYINPUT91), .B(n704), .ZN(n711) );
  NAND2_X1 U791 ( .A1(G171), .A2(n711), .ZN(n705) );
  NAND2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n716) );
  NAND2_X1 U793 ( .A1(G8), .A2(n719), .ZN(n762) );
  NOR2_X1 U794 ( .A1(G1966), .A2(n762), .ZN(n730) );
  NOR2_X1 U795 ( .A1(G2084), .A2(n719), .ZN(n727) );
  NOR2_X1 U796 ( .A1(n730), .A2(n727), .ZN(n707) );
  NAND2_X1 U797 ( .A1(G8), .A2(n707), .ZN(n708) );
  XNOR2_X1 U798 ( .A(KEYINPUT30), .B(n708), .ZN(n709) );
  NOR2_X1 U799 ( .A1(G168), .A2(n709), .ZN(n710) );
  XOR2_X1 U800 ( .A(KEYINPUT92), .B(n710), .Z(n713) );
  OR2_X1 U801 ( .A1(n711), .A2(G171), .ZN(n712) );
  NAND2_X1 U802 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U803 ( .A(n714), .B(KEYINPUT31), .ZN(n715) );
  NAND2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n728) );
  NAND2_X1 U805 ( .A1(G286), .A2(n728), .ZN(n718) );
  NOR2_X1 U806 ( .A1(G1971), .A2(n762), .ZN(n721) );
  NOR2_X1 U807 ( .A1(G2090), .A2(n719), .ZN(n720) );
  NOR2_X1 U808 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U809 ( .A1(n722), .A2(G303), .ZN(n723) );
  NAND2_X1 U810 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U811 ( .A1(n725), .A2(G8), .ZN(n726) );
  XNOR2_X1 U812 ( .A(n726), .B(KEYINPUT32), .ZN(n747) );
  NAND2_X1 U813 ( .A1(G8), .A2(n727), .ZN(n732) );
  INV_X1 U814 ( .A(n728), .ZN(n729) );
  NOR2_X1 U815 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U816 ( .A1(n732), .A2(n731), .ZN(n745) );
  AND2_X1 U817 ( .A1(n745), .A2(n762), .ZN(n733) );
  NAND2_X1 U818 ( .A1(n747), .A2(n733), .ZN(n737) );
  INV_X1 U819 ( .A(n762), .ZN(n738) );
  NOR2_X1 U820 ( .A1(G303), .A2(G2090), .ZN(n734) );
  NAND2_X1 U821 ( .A1(G8), .A2(n734), .ZN(n735) );
  OR2_X1 U822 ( .A1(n738), .A2(n735), .ZN(n736) );
  AND2_X1 U823 ( .A1(n737), .A2(n736), .ZN(n757) );
  NAND2_X1 U824 ( .A1(G1976), .A2(G288), .ZN(n896) );
  AND2_X1 U825 ( .A1(n738), .A2(n896), .ZN(n739) );
  OR2_X1 U826 ( .A1(KEYINPUT33), .A2(n739), .ZN(n742) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n750) );
  NAND2_X1 U828 ( .A1(n750), .A2(KEYINPUT33), .ZN(n740) );
  OR2_X1 U829 ( .A1(n762), .A2(n740), .ZN(n741) );
  NAND2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n744) );
  XOR2_X1 U831 ( .A(G1981), .B(G305), .Z(n911) );
  INV_X1 U832 ( .A(n911), .ZN(n743) );
  NOR2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n748) );
  AND2_X1 U834 ( .A1(n745), .A2(n748), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n755) );
  INV_X1 U836 ( .A(n748), .ZN(n753) );
  NOR2_X1 U837 ( .A1(G303), .A2(G1971), .ZN(n749) );
  NOR2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n897) );
  INV_X1 U839 ( .A(KEYINPUT33), .ZN(n751) );
  AND2_X1 U840 ( .A1(n897), .A2(n751), .ZN(n752) );
  OR2_X1 U841 ( .A1(n753), .A2(n752), .ZN(n754) );
  AND2_X1 U842 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U843 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U844 ( .A(n758), .B(KEYINPUT94), .ZN(n764) );
  NOR2_X1 U845 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XOR2_X1 U846 ( .A(n759), .B(KEYINPUT90), .Z(n760) );
  XNOR2_X1 U847 ( .A(KEYINPUT24), .B(n760), .ZN(n761) );
  NOR2_X1 U848 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U849 ( .A(n765), .B(KEYINPUT95), .ZN(n803) );
  XNOR2_X1 U850 ( .A(G1986), .B(G290), .ZN(n893) );
  NOR2_X1 U851 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U852 ( .A(n768), .B(KEYINPUT84), .ZN(n814) );
  NAND2_X1 U853 ( .A1(n893), .A2(n814), .ZN(n801) );
  INV_X1 U854 ( .A(n814), .ZN(n788) );
  NAND2_X1 U855 ( .A1(n984), .A2(G131), .ZN(n769) );
  XOR2_X1 U856 ( .A(KEYINPUT85), .B(n769), .Z(n771) );
  NAND2_X1 U857 ( .A1(n983), .A2(G95), .ZN(n770) );
  NAND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U859 ( .A(KEYINPUT86), .B(n772), .ZN(n776) );
  NAND2_X1 U860 ( .A1(G107), .A2(n979), .ZN(n774) );
  NAND2_X1 U861 ( .A1(G119), .A2(n980), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  OR2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n992) );
  AND2_X1 U864 ( .A1(n992), .A2(G1991), .ZN(n787) );
  NAND2_X1 U865 ( .A1(n983), .A2(G105), .ZN(n778) );
  XNOR2_X1 U866 ( .A(KEYINPUT38), .B(KEYINPUT88), .ZN(n777) );
  XNOR2_X1 U867 ( .A(n778), .B(n777), .ZN(n785) );
  NAND2_X1 U868 ( .A1(G141), .A2(n984), .ZN(n780) );
  NAND2_X1 U869 ( .A1(G129), .A2(n980), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G117), .A2(n979), .ZN(n781) );
  XNOR2_X1 U872 ( .A(KEYINPUT87), .B(n781), .ZN(n782) );
  NOR2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n997) );
  AND2_X1 U875 ( .A1(G1996), .A2(n997), .ZN(n786) );
  NOR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n877) );
  NOR2_X1 U877 ( .A1(n788), .A2(n877), .ZN(n806) );
  XOR2_X1 U878 ( .A(KEYINPUT89), .B(n806), .Z(n799) );
  NAND2_X1 U879 ( .A1(G104), .A2(n983), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G140), .A2(n984), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U882 ( .A(KEYINPUT34), .B(n791), .ZN(n796) );
  NAND2_X1 U883 ( .A1(G116), .A2(n979), .ZN(n793) );
  NAND2_X1 U884 ( .A1(G128), .A2(n980), .ZN(n792) );
  NAND2_X1 U885 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U886 ( .A(KEYINPUT35), .B(n794), .Z(n795) );
  NOR2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U888 ( .A(KEYINPUT36), .B(n797), .ZN(n1004) );
  XNOR2_X1 U889 ( .A(G2067), .B(KEYINPUT37), .ZN(n811) );
  NOR2_X1 U890 ( .A1(n1004), .A2(n811), .ZN(n869) );
  NAND2_X1 U891 ( .A1(n869), .A2(n814), .ZN(n809) );
  INV_X1 U892 ( .A(n809), .ZN(n798) );
  NOR2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n800) );
  AND2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n817) );
  NOR2_X1 U896 ( .A1(G1996), .A2(n997), .ZN(n872) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U898 ( .A1(G1991), .A2(n992), .ZN(n879) );
  NOR2_X1 U899 ( .A1(n804), .A2(n879), .ZN(n805) );
  NOR2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U901 ( .A1(n872), .A2(n807), .ZN(n808) );
  XNOR2_X1 U902 ( .A(n808), .B(KEYINPUT39), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U904 ( .A1(n1004), .A2(n811), .ZN(n866) );
  NAND2_X1 U905 ( .A1(n812), .A2(n866), .ZN(n813) );
  XNOR2_X1 U906 ( .A(KEYINPUT96), .B(n813), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U909 ( .A(n818), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n819), .ZN(G217) );
  NAND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n820) );
  XOR2_X1 U912 ( .A(KEYINPUT98), .B(n820), .Z(n821) );
  NAND2_X1 U913 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(G188) );
  XNOR2_X1 U916 ( .A(G120), .B(KEYINPUT99), .ZN(G236) );
  NAND2_X1 U918 ( .A1(G124), .A2(n980), .ZN(n824) );
  XNOR2_X1 U919 ( .A(n824), .B(KEYINPUT44), .ZN(n827) );
  NAND2_X1 U920 ( .A1(G100), .A2(n983), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n825), .B(KEYINPUT106), .ZN(n826) );
  NAND2_X1 U922 ( .A1(n827), .A2(n826), .ZN(n831) );
  NAND2_X1 U923 ( .A1(G112), .A2(n979), .ZN(n829) );
  NAND2_X1 U924 ( .A1(G136), .A2(n984), .ZN(n828) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U926 ( .A1(n831), .A2(n830), .ZN(G162) );
  NOR2_X1 U927 ( .A1(KEYINPUT55), .A2(G29), .ZN(n850) );
  XNOR2_X1 U928 ( .A(G2090), .B(G35), .ZN(n845) );
  XOR2_X1 U929 ( .A(G25), .B(G1991), .Z(n836) );
  XOR2_X1 U930 ( .A(G2072), .B(G33), .Z(n832) );
  NAND2_X1 U931 ( .A1(n832), .A2(G28), .ZN(n834) );
  XNOR2_X1 U932 ( .A(G26), .B(G2067), .ZN(n833) );
  NOR2_X1 U933 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U934 ( .A1(n836), .A2(n835), .ZN(n842) );
  XNOR2_X1 U935 ( .A(n837), .B(G27), .ZN(n839) );
  XNOR2_X1 U936 ( .A(G32), .B(G1996), .ZN(n838) );
  NOR2_X1 U937 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n840), .B(KEYINPUT113), .ZN(n841) );
  NOR2_X1 U939 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U940 ( .A(KEYINPUT53), .B(n843), .ZN(n844) );
  NOR2_X1 U941 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U942 ( .A(n846), .B(KEYINPUT114), .ZN(n849) );
  XOR2_X1 U943 ( .A(G2084), .B(G34), .Z(n847) );
  XNOR2_X1 U944 ( .A(KEYINPUT54), .B(n847), .ZN(n848) );
  NAND2_X1 U945 ( .A1(n849), .A2(n848), .ZN(n852) );
  NAND2_X1 U946 ( .A1(n850), .A2(n852), .ZN(n851) );
  NAND2_X1 U947 ( .A1(G11), .A2(n851), .ZN(n890) );
  INV_X1 U948 ( .A(KEYINPUT55), .ZN(n884) );
  OR2_X1 U949 ( .A1(n884), .A2(n852), .ZN(n888) );
  NAND2_X1 U950 ( .A1(G115), .A2(n979), .ZN(n854) );
  NAND2_X1 U951 ( .A1(G127), .A2(n980), .ZN(n853) );
  NAND2_X1 U952 ( .A1(n854), .A2(n853), .ZN(n856) );
  XOR2_X1 U953 ( .A(KEYINPUT108), .B(KEYINPUT47), .Z(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n861) );
  NAND2_X1 U955 ( .A1(G103), .A2(n983), .ZN(n858) );
  NAND2_X1 U956 ( .A1(G139), .A2(n984), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U958 ( .A(KEYINPUT107), .B(n859), .Z(n860) );
  NOR2_X1 U959 ( .A1(n861), .A2(n860), .ZN(n991) );
  XOR2_X1 U960 ( .A(G2072), .B(n991), .Z(n863) );
  XOR2_X1 U961 ( .A(G164), .B(G2078), .Z(n862) );
  NOR2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U963 ( .A(KEYINPUT112), .B(n864), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n865), .B(KEYINPUT50), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n867), .A2(n866), .ZN(n882) );
  XOR2_X1 U966 ( .A(G2084), .B(G160), .Z(n868) );
  NOR2_X1 U967 ( .A1(n869), .A2(n868), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n870), .A2(n996), .ZN(n875) );
  XOR2_X1 U969 ( .A(G2090), .B(G162), .Z(n871) );
  NOR2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n873), .B(KEYINPUT51), .ZN(n874) );
  NOR2_X1 U972 ( .A1(n875), .A2(n874), .ZN(n876) );
  NAND2_X1 U973 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U974 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U975 ( .A(n880), .B(KEYINPUT111), .ZN(n881) );
  NOR2_X1 U976 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U977 ( .A(n883), .B(KEYINPUT52), .ZN(n885) );
  NAND2_X1 U978 ( .A1(n885), .A2(n884), .ZN(n886) );
  NAND2_X1 U979 ( .A1(G29), .A2(n886), .ZN(n887) );
  NAND2_X1 U980 ( .A1(n888), .A2(n887), .ZN(n889) );
  NOR2_X1 U981 ( .A1(n890), .A2(n889), .ZN(n952) );
  XNOR2_X1 U982 ( .A(G16), .B(KEYINPUT56), .ZN(n919) );
  XNOR2_X1 U983 ( .A(n891), .B(G1956), .ZN(n895) );
  XNOR2_X1 U984 ( .A(G1341), .B(n681), .ZN(n892) );
  NOR2_X1 U985 ( .A1(n893), .A2(n892), .ZN(n894) );
  NAND2_X1 U986 ( .A1(n895), .A2(n894), .ZN(n903) );
  NAND2_X1 U987 ( .A1(n897), .A2(n896), .ZN(n900) );
  INV_X1 U988 ( .A(G1971), .ZN(n898) );
  NOR2_X1 U989 ( .A1(G166), .A2(n898), .ZN(n899) );
  NOR2_X1 U990 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U991 ( .A(n901), .B(KEYINPUT119), .ZN(n902) );
  NOR2_X1 U992 ( .A1(n903), .A2(n902), .ZN(n917) );
  XNOR2_X1 U993 ( .A(G171), .B(G1961), .ZN(n907) );
  XNOR2_X1 U994 ( .A(G1348), .B(KEYINPUT117), .ZN(n905) );
  XNOR2_X1 U995 ( .A(n905), .B(n904), .ZN(n906) );
  NAND2_X1 U996 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U997 ( .A(n908), .B(KEYINPUT118), .ZN(n915) );
  XNOR2_X1 U998 ( .A(KEYINPUT57), .B(KEYINPUT116), .ZN(n913) );
  XOR2_X1 U999 ( .A(G1966), .B(G168), .Z(n909) );
  XNOR2_X1 U1000 ( .A(KEYINPUT115), .B(n909), .ZN(n910) );
  NAND2_X1 U1001 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1002 ( .A(n913), .B(n912), .Z(n914) );
  NOR2_X1 U1003 ( .A1(n915), .A2(n914), .ZN(n916) );
  NAND2_X1 U1004 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1005 ( .A1(n919), .A2(n918), .ZN(n949) );
  INV_X1 U1006 ( .A(G16), .ZN(n947) );
  XNOR2_X1 U1007 ( .A(G1971), .B(G22), .ZN(n921) );
  XNOR2_X1 U1008 ( .A(G1986), .B(G24), .ZN(n920) );
  NOR2_X1 U1009 ( .A1(n921), .A2(n920), .ZN(n924) );
  XNOR2_X1 U1010 ( .A(G1976), .B(KEYINPUT123), .ZN(n922) );
  XNOR2_X1 U1011 ( .A(n922), .B(G23), .ZN(n923) );
  NAND2_X1 U1012 ( .A1(n924), .A2(n923), .ZN(n927) );
  XNOR2_X1 U1013 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n925) );
  XNOR2_X1 U1014 ( .A(n925), .B(KEYINPUT58), .ZN(n926) );
  XNOR2_X1 U1015 ( .A(n927), .B(n926), .ZN(n942) );
  XNOR2_X1 U1016 ( .A(G1966), .B(KEYINPUT122), .ZN(n928) );
  XNOR2_X1 U1017 ( .A(n928), .B(G21), .ZN(n940) );
  XNOR2_X1 U1018 ( .A(KEYINPUT59), .B(G1348), .ZN(n929) );
  XNOR2_X1 U1019 ( .A(n929), .B(G4), .ZN(n937) );
  XNOR2_X1 U1020 ( .A(G1956), .B(G20), .ZN(n935) );
  XNOR2_X1 U1021 ( .A(G1981), .B(G6), .ZN(n930) );
  XNOR2_X1 U1022 ( .A(n930), .B(KEYINPUT120), .ZN(n932) );
  XNOR2_X1 U1023 ( .A(G19), .B(G1341), .ZN(n931) );
  NOR2_X1 U1024 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1025 ( .A(KEYINPUT121), .B(n933), .ZN(n934) );
  NOR2_X1 U1026 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1027 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1028 ( .A(KEYINPUT60), .B(n938), .ZN(n939) );
  NOR2_X1 U1029 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1030 ( .A1(n942), .A2(n941), .ZN(n944) );
  XNOR2_X1 U1031 ( .A(G5), .B(G1961), .ZN(n943) );
  NOR2_X1 U1032 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1033 ( .A(KEYINPUT61), .B(n945), .ZN(n946) );
  NAND2_X1 U1034 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1035 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1036 ( .A(KEYINPUT126), .B(n950), .Z(n951) );
  NAND2_X1 U1037 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1038 ( .A(KEYINPUT62), .B(n953), .Z(G311) );
  XNOR2_X1 U1039 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1040 ( .A(G108), .ZN(G238) );
  INV_X1 U1041 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1042 ( .A1(n955), .A2(n954), .ZN(G325) );
  INV_X1 U1043 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1044 ( .A(KEYINPUT100), .B(n956), .Z(G319) );
  XOR2_X1 U1045 ( .A(KEYINPUT41), .B(G2474), .Z(n958) );
  XNOR2_X1 U1046 ( .A(G1981), .B(G1976), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(n958), .B(n957), .ZN(n959) );
  XOR2_X1 U1048 ( .A(n959), .B(KEYINPUT104), .Z(n961) );
  XNOR2_X1 U1049 ( .A(G1996), .B(KEYINPUT105), .ZN(n960) );
  XNOR2_X1 U1050 ( .A(n961), .B(n960), .ZN(n965) );
  XOR2_X1 U1051 ( .A(G1986), .B(G1971), .Z(n963) );
  XNOR2_X1 U1052 ( .A(G1966), .B(G1961), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(n963), .B(n962), .ZN(n964) );
  XOR2_X1 U1054 ( .A(n965), .B(n964), .Z(n967) );
  XNOR2_X1 U1055 ( .A(G1956), .B(G1991), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(n967), .B(n966), .ZN(G229) );
  XNOR2_X1 U1057 ( .A(G2078), .B(G2072), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(n968), .B(G2100), .ZN(n978) );
  XOR2_X1 U1059 ( .A(KEYINPUT103), .B(KEYINPUT101), .Z(n970) );
  XNOR2_X1 U1060 ( .A(KEYINPUT102), .B(KEYINPUT43), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(n970), .B(n969), .ZN(n974) );
  XOR2_X1 U1062 ( .A(G2678), .B(G2096), .Z(n972) );
  XNOR2_X1 U1063 ( .A(G2090), .B(KEYINPUT42), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(n972), .B(n971), .ZN(n973) );
  XOR2_X1 U1065 ( .A(n974), .B(n973), .Z(n976) );
  XNOR2_X1 U1066 ( .A(G2067), .B(G2084), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(n976), .B(n975), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(n978), .B(n977), .ZN(G227) );
  NAND2_X1 U1069 ( .A1(G118), .A2(n979), .ZN(n982) );
  NAND2_X1 U1070 ( .A1(G130), .A2(n980), .ZN(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n989) );
  NAND2_X1 U1072 ( .A1(G106), .A2(n983), .ZN(n986) );
  NAND2_X1 U1073 ( .A1(G142), .A2(n984), .ZN(n985) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1075 ( .A(KEYINPUT45), .B(n987), .Z(n988) );
  NOR2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(n991), .B(n990), .ZN(n1003) );
  XOR2_X1 U1078 ( .A(G164), .B(n992), .Z(n1001) );
  XOR2_X1 U1079 ( .A(KEYINPUT109), .B(KEYINPUT48), .Z(n994) );
  XNOR2_X1 U1080 ( .A(G162), .B(KEYINPUT46), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(n994), .B(n993), .ZN(n995) );
  XNOR2_X1 U1082 ( .A(n996), .B(n995), .ZN(n999) );
  XOR2_X1 U1083 ( .A(G160), .B(n997), .Z(n998) );
  XNOR2_X1 U1084 ( .A(n999), .B(n998), .ZN(n1000) );
  XNOR2_X1 U1085 ( .A(n1001), .B(n1000), .ZN(n1002) );
  XNOR2_X1 U1086 ( .A(n1003), .B(n1002), .ZN(n1005) );
  XOR2_X1 U1087 ( .A(n1005), .B(n1004), .Z(n1006) );
  NOR2_X1 U1088 ( .A1(G37), .A2(n1006), .ZN(G395) );
  XOR2_X1 U1089 ( .A(KEYINPUT110), .B(n1007), .Z(n1010) );
  XNOR2_X1 U1090 ( .A(n1008), .B(G286), .ZN(n1009) );
  XNOR2_X1 U1091 ( .A(n1010), .B(n1009), .ZN(n1012) );
  XOR2_X1 U1092 ( .A(n681), .B(G171), .Z(n1011) );
  XNOR2_X1 U1093 ( .A(n1012), .B(n1011), .ZN(n1013) );
  NOR2_X1 U1094 ( .A1(G37), .A2(n1013), .ZN(G397) );
  XOR2_X1 U1095 ( .A(G2443), .B(G2454), .Z(n1015) );
  XNOR2_X1 U1096 ( .A(G1348), .B(G2435), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(n1015), .B(n1014), .ZN(n1022) );
  XOR2_X1 U1098 ( .A(KEYINPUT97), .B(G2446), .Z(n1017) );
  XNOR2_X1 U1099 ( .A(G1341), .B(G2430), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(n1017), .B(n1016), .ZN(n1018) );
  XOR2_X1 U1101 ( .A(n1018), .B(G2451), .Z(n1020) );
  XNOR2_X1 U1102 ( .A(G2438), .B(G2427), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(n1020), .B(n1019), .ZN(n1021) );
  XNOR2_X1 U1104 ( .A(n1022), .B(n1021), .ZN(n1023) );
  NAND2_X1 U1105 ( .A1(n1023), .A2(G14), .ZN(n1029) );
  NAND2_X1 U1106 ( .A1(n1029), .A2(G319), .ZN(n1026) );
  NOR2_X1 U1107 ( .A1(G229), .A2(G227), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(KEYINPUT49), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  NOR2_X1 U1110 ( .A1(G395), .A2(G397), .ZN(n1027) );
  NAND2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(G225) );
  INV_X1 U1112 ( .A(G225), .ZN(G308) );
  INV_X1 U1113 ( .A(G69), .ZN(G235) );
  INV_X1 U1114 ( .A(n1029), .ZN(G401) );
endmodule

