

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593;

  XOR2_X1 U324 ( .A(n398), .B(n306), .Z(n535) );
  INV_X1 U325 ( .A(n368), .ZN(n334) );
  XNOR2_X1 U326 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U327 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U328 ( .A(n410), .B(KEYINPUT54), .ZN(n411) );
  XNOR2_X1 U329 ( .A(n412), .B(n411), .ZN(n570) );
  NOR2_X1 U330 ( .A1(n535), .A2(n456), .ZN(n568) );
  XNOR2_X1 U331 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U332 ( .A(n460), .B(n459), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n293) );
  XNOR2_X1 U334 ( .A(G190GAT), .B(KEYINPUT17), .ZN(n292) );
  XNOR2_X1 U335 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U336 ( .A(n294), .B(G183GAT), .Z(n296) );
  XNOR2_X1 U337 ( .A(G169GAT), .B(G176GAT), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n398) );
  XOR2_X1 U339 ( .A(G43GAT), .B(G134GAT), .Z(n379) );
  XNOR2_X1 U340 ( .A(G99GAT), .B(G71GAT), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n297), .B(G120GAT), .ZN(n332) );
  XOR2_X1 U342 ( .A(n379), .B(n332), .Z(n299) );
  NAND2_X1 U343 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U345 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n301) );
  XNOR2_X1 U346 ( .A(KEYINPUT20), .B(KEYINPUT78), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U348 ( .A(n303), .B(n302), .Z(n305) );
  XOR2_X1 U349 ( .A(G113GAT), .B(G15GAT), .Z(n314) );
  XOR2_X1 U350 ( .A(KEYINPUT0), .B(G127GAT), .Z(n416) );
  XNOR2_X1 U351 ( .A(n314), .B(n416), .ZN(n304) );
  XNOR2_X1 U352 ( .A(n305), .B(n304), .ZN(n306) );
  INV_X1 U353 ( .A(KEYINPUT55), .ZN(n455) );
  XOR2_X1 U354 ( .A(G141GAT), .B(G50GAT), .Z(n308) );
  XNOR2_X1 U355 ( .A(G43GAT), .B(G36GAT), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U357 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n310) );
  XNOR2_X1 U358 ( .A(G169GAT), .B(G197GAT), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n322) );
  XNOR2_X1 U361 ( .A(G22GAT), .B(G1GAT), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n313), .B(G8GAT), .ZN(n358) );
  XOR2_X1 U363 ( .A(n314), .B(n358), .Z(n316) );
  NAND2_X1 U364 ( .A1(G229GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U366 ( .A(n317), .B(KEYINPUT29), .Z(n320) );
  XNOR2_X1 U367 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n318), .B(KEYINPUT7), .ZN(n380) );
  XNOR2_X1 U369 ( .A(n380), .B(KEYINPUT67), .ZN(n319) );
  XNOR2_X1 U370 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n575) );
  XOR2_X1 U372 ( .A(KEYINPUT32), .B(KEYINPUT71), .Z(n324) );
  XNOR2_X1 U373 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n339) );
  XNOR2_X1 U375 ( .A(G57GAT), .B(G64GAT), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n325), .B(KEYINPUT13), .ZN(n350) );
  NAND2_X1 U377 ( .A1(n350), .A2(KEYINPUT68), .ZN(n329) );
  INV_X1 U378 ( .A(n350), .ZN(n327) );
  INV_X1 U379 ( .A(KEYINPUT68), .ZN(n326) );
  NAND2_X1 U380 ( .A1(n327), .A2(n326), .ZN(n328) );
  NAND2_X1 U381 ( .A1(n329), .A2(n328), .ZN(n331) );
  AND2_X1 U382 ( .A1(G230GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n337) );
  XNOR2_X1 U384 ( .A(G176GAT), .B(n332), .ZN(n335) );
  XNOR2_X1 U385 ( .A(G85GAT), .B(G92GAT), .ZN(n333) );
  XNOR2_X1 U386 ( .A(n333), .B(KEYINPUT70), .ZN(n368) );
  XNOR2_X1 U387 ( .A(n339), .B(n338), .ZN(n344) );
  XOR2_X1 U388 ( .A(G148GAT), .B(G106GAT), .Z(n341) );
  XNOR2_X1 U389 ( .A(G204GAT), .B(G78GAT), .ZN(n340) );
  XNOR2_X1 U390 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U391 ( .A(KEYINPUT69), .B(n342), .Z(n442) );
  INV_X1 U392 ( .A(n442), .ZN(n343) );
  XNOR2_X1 U393 ( .A(n344), .B(n343), .ZN(n580) );
  XNOR2_X1 U394 ( .A(KEYINPUT41), .B(n580), .ZN(n540) );
  NOR2_X1 U395 ( .A1(n575), .A2(n540), .ZN(n345) );
  XNOR2_X1 U396 ( .A(n345), .B(KEYINPUT46), .ZN(n363) );
  XOR2_X1 U397 ( .A(KEYINPUT76), .B(G71GAT), .Z(n347) );
  XNOR2_X1 U398 ( .A(G15GAT), .B(G127GAT), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n362) );
  XOR2_X1 U400 ( .A(G155GAT), .B(G78GAT), .Z(n349) );
  XNOR2_X1 U401 ( .A(G183GAT), .B(G211GAT), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n354) );
  XOR2_X1 U403 ( .A(KEYINPUT77), .B(n350), .Z(n352) );
  NAND2_X1 U404 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U406 ( .A(n354), .B(n353), .Z(n360) );
  XOR2_X1 U407 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n356) );
  XNOR2_X1 U408 ( .A(KEYINPUT75), .B(KEYINPUT12), .ZN(n355) );
  XNOR2_X1 U409 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U411 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U412 ( .A(n362), .B(n361), .ZN(n584) );
  NOR2_X1 U413 ( .A1(n363), .A2(n584), .ZN(n365) );
  INV_X1 U414 ( .A(KEYINPUT112), .ZN(n364) );
  XNOR2_X1 U415 ( .A(n365), .B(n364), .ZN(n385) );
  XOR2_X1 U416 ( .A(KEYINPUT64), .B(KEYINPUT10), .Z(n367) );
  XNOR2_X1 U417 ( .A(KEYINPUT73), .B(KEYINPUT65), .ZN(n366) );
  XNOR2_X1 U418 ( .A(n367), .B(n366), .ZN(n372) );
  XOR2_X1 U419 ( .A(n368), .B(G190GAT), .Z(n370) );
  NAND2_X1 U420 ( .A1(G232GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U422 ( .A(n372), .B(n371), .ZN(n384) );
  XOR2_X1 U423 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n374) );
  XNOR2_X1 U424 ( .A(G218GAT), .B(G106GAT), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U426 ( .A(n375), .B(KEYINPUT72), .Z(n377) );
  XOR2_X1 U427 ( .A(G50GAT), .B(G162GAT), .Z(n438) );
  XNOR2_X1 U428 ( .A(G99GAT), .B(n438), .ZN(n376) );
  XNOR2_X1 U429 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U430 ( .A(G36GAT), .B(KEYINPUT74), .Z(n401) );
  XOR2_X1 U431 ( .A(n378), .B(n401), .Z(n382) );
  XNOR2_X1 U432 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U433 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U434 ( .A(n384), .B(n383), .ZN(n557) );
  NOR2_X1 U435 ( .A1(n385), .A2(n557), .ZN(n386) );
  XNOR2_X1 U436 ( .A(n386), .B(KEYINPUT47), .ZN(n392) );
  INV_X1 U437 ( .A(n557), .ZN(n476) );
  XNOR2_X1 U438 ( .A(KEYINPUT36), .B(n476), .ZN(n590) );
  INV_X1 U439 ( .A(n584), .ZN(n387) );
  NOR2_X1 U440 ( .A1(n590), .A2(n387), .ZN(n388) );
  XOR2_X1 U441 ( .A(KEYINPUT45), .B(n388), .Z(n389) );
  NOR2_X1 U442 ( .A1(n580), .A2(n389), .ZN(n390) );
  NAND2_X1 U443 ( .A1(n390), .A2(n575), .ZN(n391) );
  NAND2_X1 U444 ( .A1(n392), .A2(n391), .ZN(n393) );
  XNOR2_X1 U445 ( .A(n393), .B(KEYINPUT48), .ZN(n532) );
  XNOR2_X1 U446 ( .A(G211GAT), .B(KEYINPUT84), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n394), .B(KEYINPUT21), .ZN(n395) );
  XOR2_X1 U448 ( .A(n395), .B(KEYINPUT85), .Z(n397) );
  XNOR2_X1 U449 ( .A(G197GAT), .B(G218GAT), .ZN(n396) );
  XNOR2_X1 U450 ( .A(n397), .B(n396), .ZN(n450) );
  XNOR2_X1 U451 ( .A(n398), .B(n450), .ZN(n409) );
  XOR2_X1 U452 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n400) );
  XNOR2_X1 U453 ( .A(G64GAT), .B(KEYINPUT95), .ZN(n399) );
  XNOR2_X1 U454 ( .A(n400), .B(n399), .ZN(n405) );
  XOR2_X1 U455 ( .A(G92GAT), .B(n401), .Z(n403) );
  XNOR2_X1 U456 ( .A(G8GAT), .B(G204GAT), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U458 ( .A(n405), .B(n404), .Z(n407) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U460 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U461 ( .A(n409), .B(n408), .ZN(n498) );
  NAND2_X1 U462 ( .A1(n532), .A2(n498), .ZN(n412) );
  XOR2_X1 U463 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n410) );
  XOR2_X1 U464 ( .A(G85GAT), .B(G148GAT), .Z(n414) );
  XNOR2_X1 U465 ( .A(G113GAT), .B(G134GAT), .ZN(n413) );
  XNOR2_X1 U466 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U467 ( .A(n415), .B(G162GAT), .Z(n418) );
  XNOR2_X1 U468 ( .A(G29GAT), .B(n416), .ZN(n417) );
  XNOR2_X1 U469 ( .A(n418), .B(n417), .ZN(n431) );
  XOR2_X1 U470 ( .A(KEYINPUT4), .B(G57GAT), .Z(n420) );
  XNOR2_X1 U471 ( .A(G1GAT), .B(G120GAT), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U473 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n422) );
  XNOR2_X1 U474 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U476 ( .A(n424), .B(n423), .Z(n429) );
  XOR2_X1 U477 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n426) );
  NAND2_X1 U478 ( .A1(G225GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U479 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U480 ( .A(KEYINPUT89), .B(n427), .ZN(n428) );
  XNOR2_X1 U481 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n431), .B(n430), .ZN(n437) );
  XNOR2_X1 U483 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n432) );
  XNOR2_X1 U484 ( .A(n432), .B(KEYINPUT86), .ZN(n433) );
  XOR2_X1 U485 ( .A(n433), .B(KEYINPUT87), .Z(n435) );
  XNOR2_X1 U486 ( .A(G141GAT), .B(G155GAT), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n449) );
  INV_X1 U488 ( .A(n449), .ZN(n436) );
  XOR2_X1 U489 ( .A(n437), .B(n436), .Z(n520) );
  XOR2_X1 U490 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n440) );
  XNOR2_X1 U491 ( .A(n438), .B(KEYINPUT22), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U493 ( .A(n442), .B(n441), .Z(n444) );
  NAND2_X1 U494 ( .A1(G228GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U496 ( .A(KEYINPUT82), .B(KEYINPUT88), .Z(n446) );
  XNOR2_X1 U497 ( .A(G22GAT), .B(KEYINPUT83), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U499 ( .A(n448), .B(n447), .Z(n452) );
  XNOR2_X1 U500 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U501 ( .A(n452), .B(n451), .ZN(n468) );
  NAND2_X1 U502 ( .A1(n520), .A2(n468), .ZN(n453) );
  NOR2_X1 U503 ( .A1(n570), .A2(n453), .ZN(n454) );
  XOR2_X1 U504 ( .A(n455), .B(n454), .Z(n456) );
  NAND2_X1 U505 ( .A1(n568), .A2(n557), .ZN(n460) );
  XOR2_X1 U506 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n458) );
  INV_X1 U507 ( .A(G190GAT), .ZN(n457) );
  NOR2_X1 U508 ( .A1(n575), .A2(n580), .ZN(n492) );
  INV_X1 U509 ( .A(n535), .ZN(n500) );
  XNOR2_X1 U510 ( .A(n500), .B(KEYINPUT81), .ZN(n463) );
  XOR2_X1 U511 ( .A(n498), .B(KEYINPUT27), .Z(n465) );
  NOR2_X1 U512 ( .A1(n520), .A2(n465), .ZN(n533) );
  XOR2_X1 U513 ( .A(n468), .B(KEYINPUT28), .Z(n538) );
  INV_X1 U514 ( .A(n538), .ZN(n528) );
  NAND2_X1 U515 ( .A1(n533), .A2(n528), .ZN(n461) );
  XOR2_X1 U516 ( .A(KEYINPUT96), .B(n461), .Z(n462) );
  NAND2_X1 U517 ( .A1(n463), .A2(n462), .ZN(n475) );
  NOR2_X1 U518 ( .A1(n468), .A2(n500), .ZN(n464) );
  XOR2_X1 U519 ( .A(KEYINPUT26), .B(n464), .Z(n572) );
  NOR2_X1 U520 ( .A1(n465), .A2(n572), .ZN(n466) );
  XNOR2_X1 U521 ( .A(KEYINPUT97), .B(n466), .ZN(n471) );
  NAND2_X1 U522 ( .A1(n498), .A2(n500), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n468), .A2(n467), .ZN(n469) );
  XOR2_X1 U524 ( .A(KEYINPUT25), .B(n469), .Z(n470) );
  NAND2_X1 U525 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U526 ( .A(KEYINPUT98), .B(n472), .ZN(n473) );
  NAND2_X1 U527 ( .A1(n473), .A2(n520), .ZN(n474) );
  NAND2_X1 U528 ( .A1(n475), .A2(n474), .ZN(n488) );
  NAND2_X1 U529 ( .A1(n476), .A2(n584), .ZN(n477) );
  XOR2_X1 U530 ( .A(KEYINPUT16), .B(n477), .Z(n478) );
  AND2_X1 U531 ( .A1(n488), .A2(n478), .ZN(n507) );
  NAND2_X1 U532 ( .A1(n492), .A2(n507), .ZN(n486) );
  NOR2_X1 U533 ( .A1(n520), .A2(n486), .ZN(n479) );
  XOR2_X1 U534 ( .A(KEYINPUT34), .B(n479), .Z(n480) );
  XNOR2_X1 U535 ( .A(G1GAT), .B(n480), .ZN(G1324GAT) );
  INV_X1 U536 ( .A(n498), .ZN(n523) );
  NOR2_X1 U537 ( .A1(n523), .A2(n486), .ZN(n482) );
  XNOR2_X1 U538 ( .A(G8GAT), .B(KEYINPUT99), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(G1325GAT) );
  NOR2_X1 U540 ( .A1(n535), .A2(n486), .ZN(n484) );
  XNOR2_X1 U541 ( .A(KEYINPUT35), .B(KEYINPUT100), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U543 ( .A(G15GAT), .B(n485), .ZN(G1326GAT) );
  NOR2_X1 U544 ( .A1(n528), .A2(n486), .ZN(n487) );
  XOR2_X1 U545 ( .A(G22GAT), .B(n487), .Z(G1327GAT) );
  XNOR2_X1 U546 ( .A(KEYINPUT103), .B(KEYINPUT39), .ZN(n497) );
  XOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT101), .Z(n495) );
  XNOR2_X1 U548 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n491) );
  NOR2_X1 U549 ( .A1(n590), .A2(n584), .ZN(n489) );
  NAND2_X1 U550 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n518) );
  NAND2_X1 U552 ( .A1(n518), .A2(n492), .ZN(n493) );
  XOR2_X1 U553 ( .A(KEYINPUT38), .B(n493), .Z(n504) );
  INV_X1 U554 ( .A(n520), .ZN(n571) );
  NAND2_X1 U555 ( .A1(n504), .A2(n571), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(G1328GAT) );
  NAND2_X1 U558 ( .A1(n504), .A2(n498), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n499), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT104), .B(KEYINPUT40), .Z(n502) );
  NAND2_X1 U561 ( .A1(n504), .A2(n500), .ZN(n501) );
  XNOR2_X1 U562 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U563 ( .A(G43GAT), .B(n503), .Z(G1330GAT) );
  XOR2_X1 U564 ( .A(G50GAT), .B(KEYINPUT105), .Z(n506) );
  NAND2_X1 U565 ( .A1(n538), .A2(n504), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  INV_X1 U567 ( .A(n575), .ZN(n561) );
  NOR2_X1 U568 ( .A1(n540), .A2(n561), .ZN(n517) );
  NAND2_X1 U569 ( .A1(n517), .A2(n507), .ZN(n513) );
  NOR2_X1 U570 ( .A1(n520), .A2(n513), .ZN(n508) );
  XOR2_X1 U571 ( .A(G57GAT), .B(n508), .Z(n509) );
  XNOR2_X1 U572 ( .A(KEYINPUT42), .B(n509), .ZN(G1332GAT) );
  NOR2_X1 U573 ( .A1(n523), .A2(n513), .ZN(n510) );
  XOR2_X1 U574 ( .A(G64GAT), .B(n510), .Z(G1333GAT) );
  NOR2_X1 U575 ( .A1(n535), .A2(n513), .ZN(n511) );
  XOR2_X1 U576 ( .A(KEYINPUT106), .B(n511), .Z(n512) );
  XNOR2_X1 U577 ( .A(G71GAT), .B(n512), .ZN(G1334GAT) );
  NOR2_X1 U578 ( .A1(n528), .A2(n513), .ZN(n515) );
  XNOR2_X1 U579 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(n516) );
  XOR2_X1 U581 ( .A(G78GAT), .B(n516), .Z(G1335GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(KEYINPUT108), .ZN(n529) );
  NOR2_X1 U584 ( .A1(n520), .A2(n529), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n522), .B(KEYINPUT109), .ZN(G1336GAT) );
  NOR2_X1 U587 ( .A1(n529), .A2(n523), .ZN(n524) );
  XOR2_X1 U588 ( .A(G92GAT), .B(n524), .Z(n525) );
  XNOR2_X1 U589 ( .A(KEYINPUT110), .B(n525), .ZN(G1337GAT) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n527) );
  NOR2_X1 U591 ( .A1(n535), .A2(n529), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(G1338GAT) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(n530), .Z(n531) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NAND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U597 ( .A(KEYINPUT113), .B(n534), .Z(n550) );
  NOR2_X1 U598 ( .A1(n535), .A2(n550), .ZN(n536) );
  XOR2_X1 U599 ( .A(KEYINPUT114), .B(n536), .Z(n537) );
  NOR2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n561), .A2(n547), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n539), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n542) );
  INV_X1 U604 ( .A(n540), .ZN(n563) );
  NAND2_X1 U605 ( .A1(n547), .A2(n563), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U607 ( .A(G120GAT), .B(n543), .Z(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n545) );
  NAND2_X1 U609 ( .A1(n547), .A2(n584), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n546), .Z(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U613 ( .A1(n547), .A2(n557), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  XOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT117), .Z(n552) );
  NOR2_X1 U616 ( .A1(n572), .A2(n550), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n558), .A2(n561), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U620 ( .A1(n558), .A2(n563), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n584), .A2(n558), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(KEYINPUT118), .ZN(n560) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n561), .A2(n568), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT121), .Z(n565) );
  NAND2_X1 U631 ( .A1(n568), .A2(n563), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NAND2_X1 U635 ( .A1(n584), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n574) );
  INV_X1 U638 ( .A(n572), .ZN(n573) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n589) );
  NOR2_X1 U640 ( .A1(n589), .A2(n575), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n582) );
  INV_X1 U646 ( .A(n589), .ZN(n585) );
  NAND2_X1 U647 ( .A1(n585), .A2(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n587) );
  NAND2_X1 U651 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U652 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(G211GAT), .B(n588), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U655 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

