

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  NOR2_X1 U324 ( .A1(n530), .A2(n477), .ZN(n534) );
  XNOR2_X1 U325 ( .A(KEYINPUT25), .B(KEYINPUT97), .ZN(n383) );
  XNOR2_X1 U326 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U327 ( .A(G190GAT), .B(G218GAT), .Z(n349) );
  XNOR2_X1 U328 ( .A(n318), .B(KEYINPUT9), .ZN(n319) );
  XNOR2_X1 U329 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n471) );
  XNOR2_X1 U330 ( .A(n453), .B(n319), .ZN(n320) );
  XNOR2_X1 U331 ( .A(n472), .B(n471), .ZN(n550) );
  XNOR2_X1 U332 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U333 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U334 ( .A(n329), .B(n328), .Z(n547) );
  INV_X1 U335 ( .A(G134GAT), .ZN(n483) );
  XNOR2_X1 U336 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U337 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U338 ( .A(n486), .B(n485), .ZN(G1343GAT) );
  XNOR2_X1 U339 ( .A(n459), .B(n458), .ZN(G1330GAT) );
  XOR2_X1 U340 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n293) );
  XNOR2_X1 U341 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U343 ( .A(KEYINPUT19), .B(n294), .Z(n361) );
  XOR2_X1 U344 ( .A(G120GAT), .B(G71GAT), .Z(n440) );
  XOR2_X1 U345 ( .A(G127GAT), .B(KEYINPUT0), .Z(n296) );
  XNOR2_X1 U346 ( .A(G113GAT), .B(KEYINPUT81), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n390) );
  XOR2_X1 U348 ( .A(n440), .B(n390), .Z(n298) );
  XNOR2_X1 U349 ( .A(G99GAT), .B(G190GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n298), .B(n297), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n361), .B(n299), .ZN(n312) );
  XOR2_X1 U352 ( .A(G176GAT), .B(G134GAT), .Z(n301) );
  XNOR2_X1 U353 ( .A(G169GAT), .B(G43GAT), .ZN(n300) );
  XNOR2_X1 U354 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U355 ( .A(KEYINPUT65), .B(KEYINPUT84), .Z(n303) );
  XNOR2_X1 U356 ( .A(G15GAT), .B(KEYINPUT86), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U358 ( .A(n305), .B(n304), .Z(n310) );
  XOR2_X1 U359 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n307) );
  NAND2_X1 U360 ( .A1(G227GAT), .A2(G233GAT), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U362 ( .A(KEYINPUT83), .B(n308), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n556) );
  XNOR2_X1 U365 ( .A(KEYINPUT36), .B(KEYINPUT105), .ZN(n330) );
  XOR2_X1 U366 ( .A(KEYINPUT66), .B(KEYINPUT75), .Z(n314) );
  XNOR2_X1 U367 ( .A(KEYINPUT10), .B(KEYINPUT11), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n329) );
  XOR2_X1 U369 ( .A(KEYINPUT76), .B(KEYINPUT78), .Z(n316) );
  XOR2_X1 U370 ( .A(G134GAT), .B(KEYINPUT77), .Z(n389) );
  XNOR2_X1 U371 ( .A(n389), .B(n349), .ZN(n315) );
  XOR2_X1 U372 ( .A(n316), .B(n315), .Z(n321) );
  XNOR2_X1 U373 ( .A(G99GAT), .B(G85GAT), .ZN(n317) );
  XOR2_X1 U374 ( .A(n317), .B(G92GAT), .Z(n453) );
  NAND2_X1 U375 ( .A1(G232GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n327) );
  XNOR2_X1 U377 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n322), .B(G29GAT), .ZN(n323) );
  XOR2_X1 U379 ( .A(n323), .B(KEYINPUT7), .Z(n325) );
  XNOR2_X1 U380 ( .A(G43GAT), .B(G50GAT), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n432) );
  XOR2_X1 U382 ( .A(G162GAT), .B(G106GAT), .Z(n363) );
  XNOR2_X1 U383 ( .A(n432), .B(n363), .ZN(n326) );
  XNOR2_X1 U384 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U385 ( .A(KEYINPUT79), .B(n547), .ZN(n568) );
  XNOR2_X1 U386 ( .A(n330), .B(n568), .ZN(n588) );
  XOR2_X1 U387 ( .A(G78GAT), .B(G155GAT), .Z(n332) );
  XNOR2_X1 U388 ( .A(G22GAT), .B(G183GAT), .ZN(n331) );
  XNOR2_X1 U389 ( .A(n332), .B(n331), .ZN(n346) );
  XNOR2_X1 U390 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n333), .B(KEYINPUT69), .ZN(n448) );
  XOR2_X1 U392 ( .A(n448), .B(G71GAT), .Z(n335) );
  XOR2_X1 U393 ( .A(G15GAT), .B(G1GAT), .Z(n423) );
  XNOR2_X1 U394 ( .A(n423), .B(G127GAT), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U396 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n337) );
  NAND2_X1 U397 ( .A1(G231GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U399 ( .A(n339), .B(n338), .Z(n344) );
  XOR2_X1 U400 ( .A(KEYINPUT14), .B(G64GAT), .Z(n341) );
  XNOR2_X1 U401 ( .A(G8GAT), .B(G211GAT), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n342), .B(KEYINPUT15), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U405 ( .A(n346), .B(n345), .Z(n583) );
  INV_X1 U406 ( .A(n583), .ZN(n478) );
  XOR2_X1 U407 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n348) );
  XNOR2_X1 U408 ( .A(G204GAT), .B(KEYINPUT96), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n353) );
  XOR2_X1 U410 ( .A(n349), .B(G92GAT), .Z(n351) );
  XOR2_X1 U411 ( .A(G169GAT), .B(G8GAT), .Z(n427) );
  XNOR2_X1 U412 ( .A(G36GAT), .B(n427), .ZN(n350) );
  XNOR2_X1 U413 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U414 ( .A(n353), .B(n352), .Z(n359) );
  XNOR2_X1 U415 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n354), .B(G211GAT), .ZN(n362) );
  XNOR2_X1 U417 ( .A(G176GAT), .B(G64GAT), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n355), .B(KEYINPUT72), .ZN(n447) );
  XNOR2_X1 U419 ( .A(n362), .B(n447), .ZN(n357) );
  NAND2_X1 U420 ( .A1(G226GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n361), .B(n360), .ZN(n385) );
  INV_X1 U422 ( .A(n385), .ZN(n549) );
  NAND2_X1 U423 ( .A1(n549), .A2(n556), .ZN(n382) );
  XOR2_X1 U424 ( .A(n363), .B(n362), .Z(n365) );
  NAND2_X1 U425 ( .A1(G228GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n376) );
  XOR2_X1 U427 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n367) );
  XNOR2_X1 U428 ( .A(KEYINPUT24), .B(KEYINPUT91), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U430 ( .A(n368), .B(G218GAT), .Z(n370) );
  XOR2_X1 U431 ( .A(G141GAT), .B(G22GAT), .Z(n424) );
  XNOR2_X1 U432 ( .A(G50GAT), .B(n424), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n371), .B(KEYINPUT23), .ZN(n374) );
  XNOR2_X1 U435 ( .A(G78GAT), .B(G204GAT), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n372), .B(G148GAT), .ZN(n452) );
  XOR2_X1 U437 ( .A(n452), .B(KEYINPUT92), .Z(n373) );
  XNOR2_X1 U438 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n376), .B(n375), .ZN(n381) );
  XNOR2_X1 U440 ( .A(KEYINPUT90), .B(KEYINPUT88), .ZN(n377) );
  XNOR2_X1 U441 ( .A(n377), .B(G155GAT), .ZN(n378) );
  XOR2_X1 U442 ( .A(n378), .B(KEYINPUT89), .Z(n380) );
  XNOR2_X1 U443 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n379) );
  XOR2_X1 U444 ( .A(n380), .B(n379), .Z(n394) );
  XNOR2_X1 U445 ( .A(n381), .B(n394), .ZN(n552) );
  NAND2_X1 U446 ( .A1(n382), .A2(n552), .ZN(n384) );
  XOR2_X1 U447 ( .A(KEYINPUT27), .B(n385), .Z(n409) );
  NOR2_X1 U448 ( .A1(n552), .A2(n556), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n386), .B(KEYINPUT26), .ZN(n575) );
  NAND2_X1 U450 ( .A1(n409), .A2(n575), .ZN(n387) );
  NAND2_X1 U451 ( .A1(n388), .A2(n387), .ZN(n408) );
  XOR2_X1 U452 ( .A(n389), .B(G85GAT), .Z(n392) );
  XNOR2_X1 U453 ( .A(n390), .B(G162GAT), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U455 ( .A(n394), .B(n393), .Z(n407) );
  XOR2_X1 U456 ( .A(G148GAT), .B(G120GAT), .Z(n396) );
  XNOR2_X1 U457 ( .A(G29GAT), .B(G141GAT), .ZN(n395) );
  XNOR2_X1 U458 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U459 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n398) );
  XNOR2_X1 U460 ( .A(G57GAT), .B(KEYINPUT6), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U462 ( .A(n400), .B(n399), .Z(n405) );
  XOR2_X1 U463 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n402) );
  NAND2_X1 U464 ( .A1(G225GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U465 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(n403), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n523) );
  INV_X1 U469 ( .A(n523), .ZN(n573) );
  NAND2_X1 U470 ( .A1(n408), .A2(n573), .ZN(n413) );
  XOR2_X2 U471 ( .A(KEYINPUT28), .B(n552), .Z(n530) );
  NAND2_X1 U472 ( .A1(n523), .A2(n409), .ZN(n473) );
  NOR2_X1 U473 ( .A1(n530), .A2(n473), .ZN(n411) );
  INV_X1 U474 ( .A(n556), .ZN(n410) );
  NAND2_X1 U475 ( .A1(n411), .A2(n410), .ZN(n412) );
  NAND2_X1 U476 ( .A1(n413), .A2(n412), .ZN(n414) );
  XOR2_X1 U477 ( .A(KEYINPUT98), .B(n414), .Z(n489) );
  NOR2_X1 U478 ( .A1(n478), .A2(n489), .ZN(n416) );
  INV_X1 U479 ( .A(KEYINPUT106), .ZN(n415) );
  XNOR2_X1 U480 ( .A(n416), .B(n415), .ZN(n417) );
  NOR2_X1 U481 ( .A1(n588), .A2(n417), .ZN(n418) );
  XOR2_X1 U482 ( .A(KEYINPUT37), .B(n418), .Z(n419) );
  XNOR2_X1 U483 ( .A(n419), .B(KEYINPUT107), .ZN(n522) );
  XOR2_X1 U484 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n421) );
  NAND2_X1 U485 ( .A1(G229GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U486 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U487 ( .A(n422), .B(KEYINPUT30), .Z(n426) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U490 ( .A(n428), .B(n427), .Z(n430) );
  XNOR2_X1 U491 ( .A(G113GAT), .B(G197GAT), .ZN(n429) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U493 ( .A(n432), .B(n431), .ZN(n577) );
  XOR2_X1 U494 ( .A(KEYINPUT68), .B(n577), .Z(n558) );
  INV_X1 U495 ( .A(KEYINPUT33), .ZN(n433) );
  NAND2_X1 U496 ( .A1(KEYINPUT32), .A2(n433), .ZN(n436) );
  INV_X1 U497 ( .A(KEYINPUT32), .ZN(n434) );
  NAND2_X1 U498 ( .A1(n434), .A2(KEYINPUT33), .ZN(n435) );
  NAND2_X1 U499 ( .A1(n436), .A2(n435), .ZN(n438) );
  XNOR2_X1 U500 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n437) );
  XNOR2_X1 U501 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n442) );
  AND2_X1 U503 ( .A1(G230GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U504 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U505 ( .A(KEYINPUT74), .B(KEYINPUT31), .Z(n444) );
  XNOR2_X1 U506 ( .A(KEYINPUT70), .B(KEYINPUT73), .ZN(n443) );
  XOR2_X1 U507 ( .A(n444), .B(n443), .Z(n445) );
  XNOR2_X1 U508 ( .A(n446), .B(n445), .ZN(n450) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U510 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U511 ( .A(n452), .B(n451), .ZN(n454) );
  XNOR2_X1 U512 ( .A(n454), .B(n453), .ZN(n580) );
  NAND2_X1 U513 ( .A1(n558), .A2(n580), .ZN(n491) );
  NOR2_X1 U514 ( .A1(n522), .A2(n491), .ZN(n455) );
  XNOR2_X1 U515 ( .A(KEYINPUT38), .B(n455), .ZN(n507) );
  NAND2_X1 U516 ( .A1(n556), .A2(n507), .ZN(n459) );
  XOR2_X1 U517 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n457) );
  INV_X1 U518 ( .A(G43GAT), .ZN(n456) );
  INV_X1 U519 ( .A(KEYINPUT117), .ZN(n476) );
  INV_X1 U520 ( .A(n577), .ZN(n460) );
  XNOR2_X1 U521 ( .A(KEYINPUT41), .B(n580), .ZN(n539) );
  NAND2_X1 U522 ( .A1(n460), .A2(n539), .ZN(n461) );
  XNOR2_X1 U523 ( .A(KEYINPUT46), .B(n461), .ZN(n462) );
  NAND2_X1 U524 ( .A1(n462), .A2(n583), .ZN(n463) );
  XNOR2_X1 U525 ( .A(n463), .B(KEYINPUT115), .ZN(n464) );
  NAND2_X1 U526 ( .A1(n464), .A2(n547), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n465), .B(KEYINPUT47), .ZN(n470) );
  NOR2_X1 U528 ( .A1(n583), .A2(n588), .ZN(n466) );
  XNOR2_X1 U529 ( .A(n466), .B(KEYINPUT45), .ZN(n467) );
  NAND2_X1 U530 ( .A1(n467), .A2(n580), .ZN(n468) );
  NOR2_X1 U531 ( .A1(n558), .A2(n468), .ZN(n469) );
  NOR2_X1 U532 ( .A1(n470), .A2(n469), .ZN(n472) );
  NOR2_X1 U533 ( .A1(n473), .A2(n550), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(KEYINPUT116), .ZN(n537) );
  NAND2_X1 U535 ( .A1(n537), .A2(n556), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(n477) );
  NAND2_X1 U537 ( .A1(n534), .A2(n478), .ZN(n482) );
  XOR2_X1 U538 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n480) );
  INV_X1 U539 ( .A(G127GAT), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(G1342GAT) );
  NAND2_X1 U542 ( .A1(n534), .A2(n568), .ZN(n486) );
  XOR2_X1 U543 ( .A(KEYINPUT51), .B(KEYINPUT119), .Z(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT34), .B(KEYINPUT101), .Z(n494) );
  NOR2_X1 U545 ( .A1(n583), .A2(n568), .ZN(n487) );
  XOR2_X1 U546 ( .A(KEYINPUT16), .B(n487), .Z(n488) );
  NOR2_X1 U547 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT99), .B(n490), .ZN(n509) );
  NOR2_X1 U549 ( .A1(n509), .A2(n491), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n492), .B(KEYINPUT100), .ZN(n501) );
  NAND2_X1 U551 ( .A1(n523), .A2(n501), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U553 ( .A(G1GAT), .B(n495), .ZN(G1324GAT) );
  NAND2_X1 U554 ( .A1(n501), .A2(n549), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n496), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT35), .B(KEYINPUT103), .Z(n498) );
  NAND2_X1 U557 ( .A1(n556), .A2(n501), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n500) );
  XOR2_X1 U559 ( .A(G15GAT), .B(KEYINPUT102), .Z(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  NAND2_X1 U561 ( .A1(n501), .A2(n530), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n504) );
  NAND2_X1 U564 ( .A1(n523), .A2(n507), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U566 ( .A(n505), .B(G29GAT), .ZN(G1328GAT) );
  NAND2_X1 U567 ( .A1(n507), .A2(n549), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U569 ( .A1(n507), .A2(n530), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n508), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n511) );
  NAND2_X1 U572 ( .A1(n539), .A2(n577), .ZN(n521) );
  NOR2_X1 U573 ( .A1(n521), .A2(n509), .ZN(n516) );
  NAND2_X1 U574 ( .A1(n523), .A2(n516), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  XOR2_X1 U576 ( .A(G64GAT), .B(KEYINPUT109), .Z(n513) );
  NAND2_X1 U577 ( .A1(n516), .A2(n549), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1333GAT) );
  NAND2_X1 U579 ( .A1(n516), .A2(n556), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n514), .B(KEYINPUT110), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G71GAT), .B(n515), .ZN(G1334GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U583 ( .A1(n516), .A2(n530), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n518), .B(n517), .ZN(n520) );
  XOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT112), .Z(n519) );
  XNOR2_X1 U586 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  XOR2_X1 U587 ( .A(G85GAT), .B(KEYINPUT113), .Z(n525) );
  NOR2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n529), .A2(n523), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U591 ( .A1(n529), .A2(n549), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n526), .B(KEYINPUT114), .ZN(n527) );
  XNOR2_X1 U593 ( .A(G92GAT), .B(n527), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n529), .A2(n556), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U596 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U598 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NAND2_X1 U599 ( .A1(n534), .A2(n558), .ZN(n533) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n533), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U602 ( .A1(n534), .A2(n539), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  NAND2_X1 U604 ( .A1(n537), .A2(n575), .ZN(n546) );
  NOR2_X1 U605 ( .A1(n577), .A2(n546), .ZN(n538) );
  XOR2_X1 U606 ( .A(G141GAT), .B(n538), .Z(G1344GAT) );
  INV_X1 U607 ( .A(n539), .ZN(n560) );
  NOR2_X1 U608 ( .A1(n560), .A2(n546), .ZN(n544) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT121), .Z(n541) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n540) );
  XNOR2_X1 U611 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U612 ( .A(KEYINPUT120), .B(n542), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  NOR2_X1 U614 ( .A1(n583), .A2(n546), .ZN(n545) );
  XOR2_X1 U615 ( .A(G155GAT), .B(n545), .Z(G1346GAT) );
  NOR2_X1 U616 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U617 ( .A(G162GAT), .B(n548), .Z(G1347GAT) );
  NOR2_X1 U618 ( .A1(n550), .A2(n385), .ZN(n551) );
  XNOR2_X1 U619 ( .A(KEYINPUT54), .B(n551), .ZN(n574) );
  AND2_X1 U620 ( .A1(n552), .A2(n573), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n574), .A2(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n554), .B(KEYINPUT55), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n555), .B(KEYINPUT122), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n564) );
  INV_X1 U625 ( .A(n564), .ZN(n567) );
  AND2_X1 U626 ( .A1(n558), .A2(n567), .ZN(n559) );
  XOR2_X1 U627 ( .A(G169GAT), .B(n559), .Z(G1348GAT) );
  NOR2_X1 U628 ( .A1(n560), .A2(n564), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(n563), .ZN(G1349GAT) );
  NOR2_X1 U632 ( .A1(n583), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  NAND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(KEYINPUT58), .ZN(n570) );
  XNOR2_X1 U637 ( .A(G190GAT), .B(n570), .ZN(G1351GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n572) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n572), .B(n571), .ZN(n579) );
  AND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n587) );
  NOR2_X1 U643 ( .A1(n577), .A2(n587), .ZN(n578) );
  XOR2_X1 U644 ( .A(n579), .B(n578), .Z(G1352GAT) );
  NOR2_X1 U645 ( .A1(n580), .A2(n587), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n587), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n586) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(n590) );
  NOR2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U654 ( .A(n590), .B(n589), .Z(G1355GAT) );
endmodule

