//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  AND2_X1   g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT14), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT14), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n207), .B(new_n209), .C1(new_n205), .C2(new_n206), .ZN(new_n210));
  OR3_X1    g009(.A1(new_n203), .A2(new_n204), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT93), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n211), .A2(new_n212), .B1(new_n210), .B2(new_n203), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(new_n212), .B2(new_n211), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT17), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT16), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(G1gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(KEYINPUT95), .ZN(new_n221));
  INV_X1    g020(.A(G8gat), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n217), .A2(G1gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(KEYINPUT95), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n219), .B2(KEYINPUT94), .ZN(new_n226));
  AND2_X1   g025(.A1(new_n219), .A2(KEYINPUT94), .ZN(new_n227));
  OAI21_X1  g026(.A(G8gat), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n214), .A2(new_n229), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT18), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n214), .B(new_n229), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n233), .B(KEYINPUT96), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(KEYINPUT13), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n235), .A2(new_n236), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  AND2_X1   g039(.A1(new_n232), .A2(new_n234), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(KEYINPUT18), .A3(new_n233), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT11), .ZN(new_n245));
  INV_X1    g044(.A(G169gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G197gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT12), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT92), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n250), .ZN(new_n251));
  OR2_X1    g050(.A1(new_n251), .A2(KEYINPUT97), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n240), .A2(new_n242), .A3(new_n249), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(KEYINPUT97), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT6), .ZN(new_n257));
  NAND2_X1  g056(.A1(G225gat), .A2(G233gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT2), .ZN(new_n260));
  AND2_X1   g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g062(.A1(G141gat), .A2(G148gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT81), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT81), .ZN(new_n268));
  NAND2_X1  g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n263), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n260), .A2(new_n267), .A3(new_n269), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n261), .B2(new_n262), .ZN(new_n274));
  INV_X1    g073(.A(G155gat), .ZN(new_n275));
  INV_X1    g074(.A(G162gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(KEYINPUT80), .A3(new_n259), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n272), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(KEYINPUT3), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n281), .B1(G113gat), .B2(G120gat), .ZN(new_n282));
  AND2_X1   g081(.A1(G113gat), .A2(G120gat), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT68), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G113gat), .ZN(new_n285));
  INV_X1    g084(.A(G120gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n288));
  NAND2_X1  g087(.A1(G113gat), .A2(G120gat), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n281), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g090(.A1(G127gat), .A2(G134gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(G127gat), .A2(G134gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n287), .A2(new_n281), .A3(new_n289), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n294), .B1(new_n296), .B2(KEYINPUT68), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n259), .B1(new_n277), .B2(KEYINPUT2), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n264), .A2(new_n265), .A3(KEYINPUT81), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n268), .B1(new_n267), .B2(new_n269), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT3), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n272), .A2(new_n274), .A3(new_n278), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n280), .A2(new_n299), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n305), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n299), .A2(new_n308), .A3(KEYINPUT4), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n261), .A2(new_n262), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n264), .A2(new_n265), .ZN(new_n312));
  AOI22_X1  g111(.A1(KEYINPUT80), .A2(new_n311), .B1(new_n312), .B2(new_n260), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n270), .A2(new_n266), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n313), .A2(new_n274), .B1(new_n314), .B2(new_n300), .ZN(new_n315));
  XNOR2_X1  g114(.A(G127gat), .B(G134gat), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n316), .B1(new_n284), .B2(new_n290), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(new_n297), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n310), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n258), .B(new_n307), .C1(new_n309), .C2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT82), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n295), .A2(new_n298), .A3(new_n305), .A4(new_n303), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT4), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n315), .A2(new_n318), .A3(new_n310), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n326), .A2(KEYINPUT82), .A3(new_n258), .A4(new_n307), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT5), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n271), .A2(new_n279), .B1(new_n317), .B2(new_n297), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n258), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n322), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT83), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n322), .A2(KEYINPUT83), .A3(new_n327), .A4(new_n332), .ZN(new_n336));
  INV_X1    g135(.A(new_n320), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n335), .A2(new_n336), .B1(new_n328), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT0), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(G57gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n341), .B(G85gat), .Z(new_n342));
  AOI21_X1  g141(.A(KEYINPUT84), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n338), .A2(new_n342), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n257), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n337), .A2(new_n328), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT5), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n321), .B2(new_n320), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT83), .B1(new_n349), .B2(new_n327), .ZN(new_n350));
  AND4_X1   g149(.A1(KEYINPUT83), .A2(new_n322), .A3(new_n327), .A4(new_n332), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n346), .B(new_n342), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT84), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n257), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n346), .B1(new_n350), .B2(new_n351), .ZN(new_n355));
  INV_X1    g154(.A(new_n342), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n359));
  NAND2_X1  g158(.A1(G226gat), .A2(G233gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT23), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(G169gat), .B2(G176gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n363), .A2(new_n364), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G183gat), .A2(G190gat), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT24), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372));
  AND2_X1   g171(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(G190gat), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n368), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT28), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT27), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G183gat), .ZN(new_n378));
  INV_X1    g177(.A(G183gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT27), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT66), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT66), .B1(new_n379), .B2(KEYINPUT27), .ZN(new_n382));
  INV_X1    g181(.A(G190gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n376), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT27), .B(G183gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n376), .A2(G190gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT67), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT26), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n362), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n367), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n391), .B2(new_n362), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n394), .A2(new_n396), .B1(G183gat), .B2(G190gat), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n375), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT65), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n383), .ZN(new_n400));
  NAND3_X1  g199(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT64), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n400), .B(new_n401), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n369), .A2(new_n403), .A3(new_n370), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n399), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n371), .A2(KEYINPUT64), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(new_n403), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n374), .A2(new_n407), .A3(KEYINPUT65), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n363), .A2(new_n366), .A3(new_n367), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n406), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT25), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n361), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n374), .A2(new_n371), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n411), .A2(new_n417), .A3(new_n364), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n383), .B(new_n382), .C1(new_n386), .C2(KEYINPUT66), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n419), .A2(new_n376), .B1(new_n386), .B2(new_n387), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n394), .A2(new_n396), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(new_n369), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n418), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n374), .A2(new_n407), .A3(new_n408), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n410), .B1(new_n424), .B2(new_n399), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n364), .B1(new_n425), .B2(new_n409), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n361), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT75), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT75), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n429), .A3(new_n361), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n416), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G211gat), .A2(G218gat), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT22), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT74), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n432), .A2(KEYINPUT74), .A3(new_n433), .ZN(new_n437));
  INV_X1    g236(.A(G197gat), .ZN(new_n438));
  INV_X1    g237(.A(G204gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(G197gat), .A2(G204gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n436), .A2(new_n437), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G211gat), .B(G218gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n435), .A2(new_n434), .B1(new_n440), .B2(new_n441), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(new_n444), .A3(new_n437), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n359), .B1(new_n431), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n415), .B1(new_n423), .B2(new_n426), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n360), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n429), .B1(new_n414), .B2(new_n361), .ZN(new_n453));
  AOI211_X1 g252(.A(KEYINPUT75), .B(new_n360), .C1(new_n398), .C2(new_n413), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n449), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(KEYINPUT76), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n451), .A2(KEYINPUT77), .A3(new_n360), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT77), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n427), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n460), .B2(new_n416), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n449), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n450), .A2(new_n457), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G64gat), .B(G92gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n464), .B(G36gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT78), .B(G8gat), .ZN(new_n466));
  XOR2_X1   g265(.A(new_n465), .B(new_n466), .Z(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n463), .A2(KEYINPUT79), .A3(KEYINPUT30), .A4(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT79), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n450), .A2(new_n457), .A3(new_n462), .A4(new_n468), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT30), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(new_n472), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n450), .A2(new_n457), .A3(new_n462), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n467), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n345), .A2(new_n358), .A3(new_n474), .A4(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G78gat), .B(G106gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(KEYINPUT85), .ZN(new_n481));
  NAND2_X1  g280(.A1(G228gat), .A2(G233gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n443), .A2(new_n445), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n444), .B1(new_n447), .B2(new_n437), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n415), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n315), .B1(new_n485), .B2(new_n304), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n449), .B1(new_n415), .B2(new_n306), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n482), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT86), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n490), .B(new_n482), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G22gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n306), .A2(new_n415), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n456), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT29), .B1(new_n446), .B2(new_n448), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n308), .B1(new_n496), .B2(KEYINPUT3), .ZN(new_n497));
  INV_X1    g296(.A(new_n482), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT87), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n495), .A2(new_n497), .A3(KEYINPUT87), .A4(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n492), .A2(new_n493), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n493), .B1(new_n492), .B2(new_n503), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n481), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n492), .A2(new_n503), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G22gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n481), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n493), .A3(new_n503), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT31), .B(G50gat), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n512), .B1(new_n506), .B2(new_n511), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n479), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G227gat), .A2(G233gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n398), .A2(new_n413), .A3(new_n318), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n318), .B1(new_n398), .B2(new_n413), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT69), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI211_X1 g322(.A(KEYINPUT69), .B(new_n318), .C1(new_n398), .C2(new_n413), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G43gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(G71gat), .B(G99gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT33), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n525), .A2(KEYINPUT32), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT71), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n525), .A2(new_n533), .A3(KEYINPUT32), .A4(new_n530), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n525), .A2(KEYINPUT32), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT70), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT70), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n525), .A2(new_n538), .A3(KEYINPUT32), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n528), .B1(new_n525), .B2(new_n529), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n414), .A2(new_n299), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT69), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n521), .A2(new_n522), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n544), .A2(new_n518), .A3(new_n545), .A4(new_n520), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT72), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n546), .A2(new_n547), .A3(KEYINPUT34), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n547), .B1(new_n546), .B2(KEYINPUT34), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n546), .A2(KEYINPUT34), .ZN(new_n550));
  OR3_X1    g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n542), .A2(new_n551), .ZN(new_n552));
  NOR3_X1   g351(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(new_n535), .A3(new_n541), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(KEYINPUT73), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT73), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n557), .A3(new_n551), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n552), .A2(KEYINPUT36), .A3(new_n554), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT39), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n258), .B1(new_n326), .B2(new_n307), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n356), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT39), .B1(new_n330), .B2(new_n331), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g365(.A1(KEYINPUT89), .A2(KEYINPUT40), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n566), .B(new_n567), .Z(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n357), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n474), .A2(new_n478), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT88), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT88), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n474), .A2(new_n572), .A3(new_n478), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n569), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n471), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n476), .A2(KEYINPUT37), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT37), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n450), .A2(new_n457), .A3(new_n462), .A4(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n467), .A3(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT90), .B(KEYINPUT38), .Z(new_n580));
  AOI21_X1  g379(.A(new_n575), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n577), .B1(new_n461), .B2(new_n456), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n455), .A2(new_n449), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(new_n578), .A3(new_n467), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT91), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT91), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n584), .A2(new_n578), .A3(new_n587), .A4(new_n467), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n352), .A2(new_n353), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT6), .B1(new_n590), .B2(new_n357), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n338), .A2(KEYINPUT84), .A3(new_n342), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n344), .B1(new_n257), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n581), .B(new_n589), .C1(new_n591), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n515), .ZN(new_n595));
  OAI211_X1 g394(.A(new_n517), .B(new_n561), .C1(new_n574), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n506), .A2(new_n511), .ZN(new_n597));
  INV_X1    g396(.A(new_n512), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n599), .A2(new_n552), .A3(new_n600), .A4(new_n554), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT35), .B1(new_n479), .B2(new_n601), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n513), .A2(new_n514), .A3(KEYINPUT35), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n590), .A2(new_n357), .ZN(new_n604));
  AOI22_X1  g403(.A1(new_n604), .A2(new_n257), .B1(new_n354), .B2(new_n357), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n554), .A2(KEYINPUT73), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n553), .B1(new_n535), .B2(new_n541), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n558), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n603), .B(new_n605), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n571), .A2(new_n573), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n602), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n256), .B1(new_n596), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G85gat), .A2(G92gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT7), .ZN(new_n615));
  INV_X1    g414(.A(G99gat), .ZN(new_n616));
  INV_X1    g415(.A(G106gat), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT8), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT102), .B(G85gat), .Z(new_n619));
  OAI211_X1 g418(.A(new_n615), .B(new_n618), .C1(G92gat), .C2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G99gat), .B(G106gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n216), .A2(new_n231), .A3(new_n623), .ZN(new_n624));
  AND3_X1   g423(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n625), .B1(new_n214), .B2(new_n622), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n624), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n624), .B2(new_n626), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(G190gat), .B(G218gat), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n637), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(new_n634), .B2(new_n635), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(G57gat), .B(G64gat), .Z(new_n642));
  INV_X1    g441(.A(KEYINPUT9), .ZN(new_n643));
  INV_X1    g442(.A(G71gat), .ZN(new_n644));
  INV_X1    g443(.A(G78gat), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(G71gat), .B(G78gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT101), .Z(new_n650));
  AOI21_X1  g449(.A(new_n229), .B1(new_n650), .B2(KEYINPUT21), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(new_n379), .ZN(new_n652));
  NAND2_X1  g451(.A1(G231gat), .A2(G233gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT99), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT100), .ZN(new_n655));
  XOR2_X1   g454(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n652), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(KEYINPUT98), .B(KEYINPUT21), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n649), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(G127gat), .B(G155gat), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G211gat), .ZN(new_n663));
  OR2_X1    g462(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n658), .A2(new_n663), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n622), .B(new_n649), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT10), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n650), .A2(KEYINPUT10), .A3(new_n622), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(G230gat), .ZN(new_n672));
  INV_X1    g471(.A(G233gat), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(G230gat), .A2(G233gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n675), .B2(new_n667), .ZN(new_n676));
  XNOR2_X1  g475(.A(G120gat), .B(G148gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G176gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(new_n439), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n680), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n641), .A2(new_n666), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n613), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n685), .A2(new_n605), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(G1gat), .Z(G1324gat));
  INV_X1    g486(.A(new_n611), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  AND2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n691), .A2(KEYINPUT42), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(KEYINPUT42), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n692), .B(new_n693), .C1(new_n222), .C2(new_n689), .ZN(G1325gat));
  AND3_X1   g493(.A1(new_n559), .A2(KEYINPUT105), .A3(new_n560), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT105), .B1(new_n559), .B2(new_n560), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G15gat), .B1(new_n685), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n608), .A2(new_n609), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n699), .A2(G15gat), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n685), .B2(new_n700), .ZN(G1326gat));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n515), .ZN(new_n702));
  XNOR2_X1  g501(.A(KEYINPUT43), .B(G22gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT106), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n702), .B(new_n704), .ZN(G1327gat));
  INV_X1    g504(.A(new_n605), .ZN(new_n706));
  INV_X1    g505(.A(new_n641), .ZN(new_n707));
  INV_X1    g506(.A(new_n683), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n666), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n613), .A2(new_n205), .A3(new_n706), .A4(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT45), .Z(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n596), .A2(new_n612), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(new_n641), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n561), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n559), .A2(KEYINPUT105), .A3(new_n560), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n517), .B1(new_n574), .B2(new_n595), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n716), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n517), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n594), .A2(new_n515), .ZN(new_n724));
  INV_X1    g523(.A(new_n573), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n572), .B1(new_n474), .B2(new_n478), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n357), .B(new_n568), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n723), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(new_n697), .A3(KEYINPUT107), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n612), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n602), .B(KEYINPUT108), .C1(new_n610), .C2(new_n611), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n722), .A2(new_n729), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n641), .A2(new_n713), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n715), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n737), .A2(new_n256), .A3(new_n709), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n706), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n712), .B1(new_n739), .B2(G29gat), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT109), .Z(G1328gat));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742));
  AOI21_X1  g541(.A(G36gat), .B1(new_n742), .B2(KEYINPUT46), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n613), .A2(new_n611), .A3(new_n710), .A4(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n742), .B2(KEYINPUT46), .ZN(new_n745));
  OR3_X1    g544(.A1(new_n744), .A2(new_n742), .A3(KEYINPUT46), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n738), .A2(new_n611), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n745), .B(new_n746), .C1(new_n747), .C2(new_n206), .ZN(G1329gat));
  INV_X1    g547(.A(G43gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n738), .A2(new_n720), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(KEYINPUT111), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(KEYINPUT111), .B2(new_n750), .ZN(new_n752));
  INV_X1    g551(.A(new_n699), .ZN(new_n753));
  AND4_X1   g552(.A1(new_n749), .A2(new_n613), .A3(new_n753), .A4(new_n710), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT47), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n749), .B1(new_n738), .B2(new_n720), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n755), .B1(new_n758), .B2(new_n754), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(G1330gat));
  INV_X1    g559(.A(G50gat), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n738), .B2(new_n516), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT112), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n516), .A2(new_n761), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n710), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n762), .B1(new_n613), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g567(.A1(new_n641), .A2(new_n666), .ZN(new_n769));
  AND4_X1   g568(.A1(new_n256), .A2(new_n734), .A3(new_n769), .A4(new_n683), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n706), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n611), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT49), .B(G64gat), .Z(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n773), .B2(new_n775), .ZN(G1333gat));
  AOI21_X1  g575(.A(new_n644), .B1(new_n770), .B2(new_n720), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n699), .A2(G71gat), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n770), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g579(.A1(new_n770), .A2(new_n516), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g581(.A1(new_n256), .A2(new_n666), .A3(new_n683), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n728), .A2(new_n697), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n785), .A2(new_n716), .B1(new_n731), .B2(new_n732), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n735), .B1(new_n786), .B2(new_n729), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n784), .B1(new_n787), .B2(new_n715), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n619), .B1(new_n788), .B2(new_n605), .ZN(new_n789));
  INV_X1    g588(.A(new_n666), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n707), .A2(new_n255), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n734), .A2(KEYINPUT51), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT51), .B1(new_n734), .B2(new_n791), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n683), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n605), .A2(new_n619), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n789), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(KEYINPUT113), .Z(G1336gat));
  OAI21_X1  g597(.A(G92gat), .B1(new_n788), .B2(new_n688), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n734), .A2(new_n791), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(KEYINPUT114), .A3(new_n792), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n794), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n688), .A2(G92gat), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n683), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n799), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT52), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  INV_X1    g610(.A(new_n807), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n799), .B(new_n811), .C1(new_n795), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(G1337gat));
  NOR3_X1   g613(.A1(new_n788), .A2(new_n616), .A3(new_n697), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n795), .A2(new_n699), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n815), .B1(new_n816), .B2(new_n616), .ZN(G1338gat));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n737), .A2(new_n515), .A3(new_n783), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n819), .B2(new_n617), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n708), .A2(new_n515), .A3(G106gat), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n803), .A2(new_n805), .A3(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n516), .B(new_n784), .C1(new_n787), .C2(new_n715), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n823), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n820), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT53), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n821), .B1(new_n793), .B2(new_n794), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n827), .B(new_n828), .C1(new_n617), .C2(new_n819), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n826), .A2(KEYINPUT116), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1339gat));
  NAND3_X1  g633(.A1(new_n769), .A2(new_n256), .A3(new_n708), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n669), .A2(new_n670), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n672), .A2(new_n673), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(KEYINPUT54), .A3(new_n674), .ZN(new_n840));
  OR3_X1    g639(.A1(new_n837), .A2(KEYINPUT54), .A3(new_n838), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n841), .A3(new_n680), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(new_n681), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n844), .A2(KEYINPUT117), .A3(new_n681), .A4(new_n845), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n241), .A2(new_n233), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n237), .A2(new_n239), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n248), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n253), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n638), .B2(new_n640), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n850), .A2(new_n851), .A3(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n851), .B1(new_n850), .B2(new_n856), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n708), .A2(new_n855), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n850), .B2(new_n255), .ZN(new_n861));
  OAI22_X1  g660(.A1(new_n858), .A2(new_n859), .B1(new_n861), .B2(new_n641), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n836), .B1(new_n862), .B2(new_n666), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n863), .A2(new_n516), .A3(new_n699), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n611), .A2(new_n605), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(new_n285), .A3(new_n256), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n863), .A2(new_n601), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n865), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(G113gat), .B1(new_n870), .B2(new_n255), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n867), .A2(new_n871), .ZN(G1340gat));
  NOR3_X1   g671(.A1(new_n866), .A2(new_n286), .A3(new_n708), .ZN(new_n873));
  AOI21_X1  g672(.A(G120gat), .B1(new_n870), .B2(new_n683), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(G1341gat));
  OAI21_X1  g674(.A(G127gat), .B1(new_n866), .B2(new_n666), .ZN(new_n876));
  OR2_X1    g675(.A1(new_n666), .A2(G127gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n869), .B2(new_n877), .ZN(G1342gat));
  OAI21_X1  g677(.A(G134gat), .B1(new_n866), .B2(new_n707), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n869), .A2(G134gat), .A3(new_n707), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT119), .B1(new_n880), .B2(KEYINPUT56), .ZN(new_n883));
  OAI221_X1 g682(.A(new_n879), .B1(KEYINPUT56), .B2(new_n880), .C1(new_n882), .C2(new_n883), .ZN(G1343gat));
  NAND2_X1  g683(.A1(new_n850), .A2(new_n856), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT118), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n857), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n256), .A2(new_n846), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n707), .B1(new_n888), .B2(new_n860), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n836), .B1(new_n890), .B2(new_n666), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT57), .B1(new_n891), .B2(new_n515), .ZN(new_n892));
  INV_X1    g691(.A(new_n865), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n720), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n861), .A2(new_n641), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n790), .B1(new_n896), .B2(new_n887), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n895), .B(new_n516), .C1(new_n897), .C2(new_n836), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n892), .A2(new_n894), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G141gat), .B1(new_n899), .B2(new_n256), .ZN(new_n900));
  NOR4_X1   g699(.A1(new_n863), .A2(new_n515), .A3(new_n720), .A4(new_n893), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n256), .A2(G141gat), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n901), .A2(new_n902), .B1(new_n903), .B2(KEYINPUT58), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n903), .A2(KEYINPUT58), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n905), .B(new_n906), .Z(G1344gat));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT57), .B1(new_n863), .B2(new_n515), .ZN(new_n909));
  INV_X1    g708(.A(new_n846), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n856), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n790), .B1(new_n889), .B2(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n895), .B(new_n516), .C1(new_n912), .C2(new_n836), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n894), .A2(KEYINPUT122), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n909), .A2(new_n683), .A3(new_n913), .A4(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n894), .A2(KEYINPUT122), .ZN(new_n916));
  OAI21_X1  g715(.A(G148gat), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n892), .A2(new_n683), .A3(new_n894), .A4(new_n898), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n919), .A2(G148gat), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n917), .A2(KEYINPUT59), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(G148gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n901), .A2(new_n922), .A3(new_n683), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT121), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n908), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n923), .B(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n913), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n516), .B1(new_n897), .B2(new_n836), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(KEYINPUT57), .ZN(new_n930));
  INV_X1    g729(.A(new_n916), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n930), .A2(new_n683), .A3(new_n931), .A4(new_n914), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n919), .B1(new_n932), .B2(G148gat), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n918), .A2(new_n920), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n927), .B(KEYINPUT123), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n925), .A2(new_n935), .ZN(G1345gat));
  OAI21_X1  g735(.A(G155gat), .B1(new_n899), .B2(new_n666), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n901), .A2(new_n275), .A3(new_n790), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1346gat));
  NAND3_X1  g738(.A1(new_n901), .A2(new_n276), .A3(new_n641), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n899), .A2(new_n707), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(KEYINPUT124), .ZN(new_n942));
  OAI21_X1  g741(.A(G162gat), .B1(new_n941), .B2(KEYINPUT124), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(G1347gat));
  NOR2_X1   g743(.A1(new_n688), .A2(new_n706), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n868), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n246), .B1(new_n946), .B2(new_n256), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n864), .A2(G169gat), .A3(new_n255), .A4(new_n945), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(G1348gat));
  NAND2_X1  g748(.A1(new_n864), .A2(new_n945), .ZN(new_n950));
  OAI21_X1  g749(.A(G176gat), .B1(new_n950), .B2(new_n708), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n708), .A2(G176gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n946), .B2(new_n952), .ZN(G1349gat));
  INV_X1    g752(.A(KEYINPUT60), .ZN(new_n954));
  OAI21_X1  g753(.A(G183gat), .B1(new_n950), .B2(new_n666), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n868), .A2(new_n386), .A3(new_n790), .A4(new_n945), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n957), .B1(new_n955), .B2(new_n956), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n954), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(new_n960), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n962), .A2(KEYINPUT60), .A3(new_n958), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n961), .A2(new_n963), .ZN(G1350gat));
  NAND3_X1  g763(.A1(new_n864), .A2(new_n641), .A3(new_n945), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n965), .A2(new_n966), .A3(G190gat), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n966), .B1(new_n965), .B2(G190gat), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n641), .A2(new_n383), .ZN(new_n970));
  OAI22_X1  g769(.A1(new_n968), .A2(new_n969), .B1(new_n946), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(KEYINPUT126), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n973));
  OAI221_X1 g772(.A(new_n973), .B1(new_n946), .B2(new_n970), .C1(new_n968), .C2(new_n969), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1351gat));
  NAND2_X1  g774(.A1(new_n697), .A2(new_n945), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n929), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n977), .A2(new_n438), .A3(new_n255), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n909), .A2(new_n913), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n979), .A2(new_n256), .A3(new_n976), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n978), .B1(new_n980), .B2(new_n438), .ZN(G1352gat));
  NOR3_X1   g780(.A1(new_n979), .A2(new_n708), .A3(new_n976), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n982), .A2(new_n439), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n977), .A2(new_n439), .A3(new_n683), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n983), .B1(KEYINPUT62), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n985), .B1(KEYINPUT62), .B2(new_n984), .ZN(G1353gat));
  INV_X1    g785(.A(G211gat), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n977), .A2(new_n987), .A3(new_n790), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n979), .A2(new_n976), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(new_n790), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n990), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT63), .B1(new_n990), .B2(G211gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  AOI21_X1  g792(.A(G218gat), .B1(new_n977), .B2(new_n641), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT127), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n641), .A2(G218gat), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n995), .B1(new_n989), .B2(new_n996), .ZN(G1355gat));
endmodule


