

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  NOR2_X1 U323 ( .A1(n569), .A2(n389), .ZN(n469) );
  XNOR2_X1 U324 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U325 ( .A(n413), .B(n412), .Z(n563) );
  NOR2_X1 U326 ( .A1(n511), .A2(n481), .ZN(n448) );
  XOR2_X1 U327 ( .A(n427), .B(G92GAT), .Z(n291) );
  XOR2_X1 U328 ( .A(G29GAT), .B(G43GAT), .Z(n292) );
  XOR2_X1 U329 ( .A(n550), .B(n549), .Z(n293) );
  INV_X1 U330 ( .A(KEYINPUT19), .ZN(n302) );
  INV_X1 U331 ( .A(KEYINPUT97), .ZN(n395) );
  XNOR2_X1 U332 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n549) );
  XNOR2_X1 U333 ( .A(n303), .B(n302), .ZN(n305) );
  XNOR2_X1 U334 ( .A(n305), .B(n304), .ZN(n352) );
  XNOR2_X1 U335 ( .A(n444), .B(n443), .ZN(n446) );
  XNOR2_X1 U336 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U337 ( .A(n360), .B(n359), .ZN(n366) );
  XOR2_X1 U338 ( .A(n453), .B(n575), .Z(n540) );
  NOR2_X1 U339 ( .A1(n512), .A2(n502), .ZN(n508) );
  XNOR2_X1 U340 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n474) );
  XNOR2_X1 U341 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U342 ( .A(n475), .B(n474), .ZN(G1342GAT) );
  XNOR2_X1 U343 ( .A(n452), .B(n451), .ZN(G1330GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n295) );
  XNOR2_X1 U345 ( .A(G169GAT), .B(G120GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n313) );
  XOR2_X1 U347 ( .A(G99GAT), .B(G190GAT), .Z(n297) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G134GAT), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U350 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n299) );
  XNOR2_X1 U351 ( .A(G15GAT), .B(G71GAT), .ZN(n298) );
  XNOR2_X1 U352 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U353 ( .A(n301), .B(n300), .Z(n311) );
  XNOR2_X1 U354 ( .A(KEYINPUT82), .B(G183GAT), .ZN(n303) );
  XOR2_X1 U355 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n304) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n306), .B(G127GAT), .ZN(n339) );
  XOR2_X1 U358 ( .A(n339), .B(G176GAT), .Z(n308) );
  NAND2_X1 U359 ( .A1(G227GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n352), .B(n309), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n518) );
  INV_X1 U364 ( .A(n518), .ZN(n555) );
  XOR2_X1 U365 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n315) );
  XNOR2_X1 U366 ( .A(G64GAT), .B(KEYINPUT78), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n327) );
  XOR2_X1 U368 ( .A(G183GAT), .B(G78GAT), .Z(n317) );
  XNOR2_X1 U369 ( .A(G211GAT), .B(G155GAT), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n317), .B(n316), .ZN(n325) );
  XOR2_X1 U371 ( .A(KEYINPUT79), .B(KEYINPUT15), .Z(n319) );
  XNOR2_X1 U372 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U374 ( .A(KEYINPUT75), .B(G57GAT), .Z(n321) );
  XNOR2_X1 U375 ( .A(G8GAT), .B(G127GAT), .ZN(n320) );
  XNOR2_X1 U376 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U377 ( .A(n323), .B(n322), .Z(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U379 ( .A(n327), .B(n326), .ZN(n332) );
  XNOR2_X1 U380 ( .A(G22GAT), .B(G15GAT), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n328), .B(G1GAT), .ZN(n422) );
  XOR2_X1 U382 ( .A(G71GAT), .B(KEYINPUT13), .Z(n440) );
  XOR2_X1 U383 ( .A(n422), .B(n440), .Z(n330) );
  NAND2_X1 U384 ( .A1(G231GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U386 ( .A(n332), .B(n331), .Z(n579) );
  XOR2_X1 U387 ( .A(G155GAT), .B(KEYINPUT2), .Z(n334) );
  XNOR2_X1 U388 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n334), .B(n333), .ZN(n370) );
  XOR2_X1 U390 ( .A(n370), .B(G1GAT), .Z(n336) );
  NAND2_X1 U391 ( .A1(G225GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n338) );
  XOR2_X1 U393 ( .A(G120GAT), .B(G57GAT), .Z(n445) );
  INV_X1 U394 ( .A(n445), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n341) );
  XOR2_X1 U396 ( .A(G134GAT), .B(KEYINPUT73), .Z(n400) );
  XNOR2_X1 U397 ( .A(n339), .B(n400), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n349) );
  XOR2_X1 U399 ( .A(G85GAT), .B(G148GAT), .Z(n343) );
  XNOR2_X1 U400 ( .A(G29GAT), .B(G162GAT), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U402 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n345) );
  XNOR2_X1 U403 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U405 ( .A(n347), .B(n346), .Z(n348) );
  XOR2_X1 U406 ( .A(n349), .B(n348), .Z(n514) );
  INV_X1 U407 ( .A(n514), .ZN(n569) );
  XOR2_X1 U408 ( .A(KEYINPUT88), .B(KEYINPUT90), .Z(n354) );
  XOR2_X1 U409 ( .A(G64GAT), .B(G92GAT), .Z(n351) );
  XNOR2_X1 U410 ( .A(G204GAT), .B(G176GAT), .ZN(n350) );
  XNOR2_X1 U411 ( .A(n351), .B(n350), .ZN(n436) );
  XNOR2_X1 U412 ( .A(n352), .B(n436), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n360) );
  XOR2_X1 U414 ( .A(KEYINPUT89), .B(KEYINPUT75), .Z(n356) );
  XOR2_X1 U415 ( .A(G169GAT), .B(G8GAT), .Z(n423) );
  XOR2_X1 U416 ( .A(G36GAT), .B(G190GAT), .Z(n399) );
  XNOR2_X1 U417 ( .A(n423), .B(n399), .ZN(n355) );
  XNOR2_X1 U418 ( .A(n356), .B(n355), .ZN(n358) );
  AND2_X1 U419 ( .A1(G226GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U420 ( .A(G211GAT), .B(KEYINPUT86), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n361), .B(KEYINPUT21), .ZN(n362) );
  XOR2_X1 U422 ( .A(n362), .B(KEYINPUT87), .Z(n364) );
  XNOR2_X1 U423 ( .A(G197GAT), .B(G218GAT), .ZN(n363) );
  XOR2_X1 U424 ( .A(n364), .B(n363), .Z(n378) );
  INV_X1 U425 ( .A(n378), .ZN(n365) );
  XOR2_X1 U426 ( .A(n366), .B(n365), .Z(n495) );
  INV_X1 U427 ( .A(n495), .ZN(n548) );
  XOR2_X1 U428 ( .A(n548), .B(KEYINPUT27), .Z(n389) );
  XNOR2_X1 U429 ( .A(G106GAT), .B(G78GAT), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n367), .B(G148GAT), .ZN(n435) );
  XOR2_X1 U431 ( .A(KEYINPUT22), .B(n435), .Z(n369) );
  XOR2_X1 U432 ( .A(G50GAT), .B(G162GAT), .Z(n409) );
  XNOR2_X1 U433 ( .A(G22GAT), .B(n409), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n374) );
  XOR2_X1 U435 ( .A(n370), .B(G204GAT), .Z(n372) );
  NAND2_X1 U436 ( .A1(G228GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U438 ( .A(n374), .B(n373), .Z(n380) );
  XOR2_X1 U439 ( .A(KEYINPUT23), .B(KEYINPUT85), .Z(n376) );
  XNOR2_X1 U440 ( .A(KEYINPUT84), .B(KEYINPUT24), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U442 ( .A(n378), .B(n377), .Z(n379) );
  XNOR2_X1 U443 ( .A(n380), .B(n379), .ZN(n551) );
  XNOR2_X1 U444 ( .A(KEYINPUT28), .B(KEYINPUT65), .ZN(n381) );
  XOR2_X1 U445 ( .A(n551), .B(n381), .Z(n498) );
  NAND2_X1 U446 ( .A1(n469), .A2(n498), .ZN(n382) );
  XOR2_X1 U447 ( .A(KEYINPUT91), .B(n382), .Z(n383) );
  NOR2_X1 U448 ( .A1(n518), .A2(n383), .ZN(n394) );
  NAND2_X1 U449 ( .A1(n518), .A2(n548), .ZN(n384) );
  NAND2_X1 U450 ( .A1(n384), .A2(n551), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n385), .B(KEYINPUT93), .ZN(n386) );
  XOR2_X1 U452 ( .A(KEYINPUT25), .B(n386), .Z(n391) );
  NOR2_X1 U453 ( .A1(n551), .A2(n518), .ZN(n388) );
  XNOR2_X1 U454 ( .A(KEYINPUT26), .B(KEYINPUT92), .ZN(n387) );
  XOR2_X1 U455 ( .A(n388), .B(n387), .Z(n570) );
  NOR2_X1 U456 ( .A1(n570), .A2(n389), .ZN(n390) );
  NOR2_X1 U457 ( .A1(n391), .A2(n390), .ZN(n392) );
  NOR2_X1 U458 ( .A1(n514), .A2(n392), .ZN(n393) );
  NOR2_X1 U459 ( .A1(n394), .A2(n393), .ZN(n478) );
  NOR2_X1 U460 ( .A1(n579), .A2(n478), .ZN(n396) );
  XNOR2_X1 U461 ( .A(n396), .B(n395), .ZN(n414) );
  XOR2_X1 U462 ( .A(KEYINPUT11), .B(KEYINPUT71), .Z(n398) );
  XNOR2_X1 U463 ( .A(G218GAT), .B(G106GAT), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n398), .B(n397), .ZN(n413) );
  XNOR2_X1 U465 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U466 ( .A(G99GAT), .B(G85GAT), .Z(n441) );
  XNOR2_X1 U467 ( .A(n401), .B(n441), .ZN(n405) );
  XNOR2_X1 U468 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n402) );
  XNOR2_X1 U469 ( .A(n292), .B(n402), .ZN(n427) );
  NAND2_X1 U470 ( .A1(G232GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U471 ( .A(n291), .B(n403), .ZN(n404) );
  XOR2_X1 U472 ( .A(n405), .B(n404), .Z(n411) );
  XOR2_X1 U473 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n407) );
  XNOR2_X1 U474 ( .A(KEYINPUT72), .B(KEYINPUT10), .ZN(n406) );
  XNOR2_X1 U475 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U476 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U477 ( .A(n411), .B(n410), .ZN(n412) );
  INV_X1 U478 ( .A(n563), .ZN(n457) );
  XOR2_X1 U479 ( .A(KEYINPUT36), .B(n457), .Z(n583) );
  NAND2_X1 U480 ( .A1(n414), .A2(n583), .ZN(n415) );
  XOR2_X1 U481 ( .A(KEYINPUT37), .B(n415), .Z(n511) );
  XOR2_X1 U482 ( .A(G197GAT), .B(G141GAT), .Z(n417) );
  XNOR2_X1 U483 ( .A(G50GAT), .B(G36GAT), .ZN(n416) );
  XNOR2_X1 U484 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U485 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n419) );
  XNOR2_X1 U486 ( .A(G113GAT), .B(KEYINPUT30), .ZN(n418) );
  XNOR2_X1 U487 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U488 ( .A(n421), .B(n420), .ZN(n431) );
  XOR2_X1 U489 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U490 ( .A1(G229GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U492 ( .A(n426), .B(KEYINPUT68), .Z(n429) );
  XNOR2_X1 U493 ( .A(n427), .B(KEYINPUT67), .ZN(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U495 ( .A(n431), .B(n430), .Z(n501) );
  INV_X1 U496 ( .A(n501), .ZN(n572) );
  XOR2_X1 U497 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n433) );
  NAND2_X1 U498 ( .A1(G230GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U499 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U500 ( .A(n434), .B(KEYINPUT69), .Z(n438) );
  XNOR2_X1 U501 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U502 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U503 ( .A(n439), .B(KEYINPUT70), .ZN(n444) );
  XOR2_X1 U504 ( .A(n440), .B(KEYINPUT31), .Z(n442) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n575) );
  INV_X1 U506 ( .A(n575), .ZN(n465) );
  NAND2_X1 U507 ( .A1(n572), .A2(n465), .ZN(n481) );
  XOR2_X1 U508 ( .A(KEYINPUT38), .B(KEYINPUT98), .Z(n447) );
  XNOR2_X1 U509 ( .A(n448), .B(n447), .ZN(n497) );
  NOR2_X1 U510 ( .A1(n555), .A2(n497), .ZN(n452) );
  XNOR2_X1 U511 ( .A(KEYINPUT40), .B(KEYINPUT100), .ZN(n450) );
  INV_X1 U512 ( .A(G43GAT), .ZN(n449) );
  INV_X1 U513 ( .A(n498), .ZN(n522) );
  XNOR2_X1 U514 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n453) );
  NAND2_X1 U515 ( .A1(n572), .A2(n540), .ZN(n454) );
  XNOR2_X1 U516 ( .A(n454), .B(KEYINPUT46), .ZN(n455) );
  INV_X1 U517 ( .A(n579), .ZN(n476) );
  NAND2_X1 U518 ( .A1(n455), .A2(n476), .ZN(n456) );
  XNOR2_X1 U519 ( .A(n456), .B(KEYINPUT109), .ZN(n458) );
  NAND2_X1 U520 ( .A1(n458), .A2(n457), .ZN(n460) );
  XOR2_X1 U521 ( .A(KEYINPUT47), .B(KEYINPUT110), .Z(n459) );
  XNOR2_X1 U522 ( .A(n460), .B(n459), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n583), .A2(n579), .ZN(n462) );
  XOR2_X1 U524 ( .A(KEYINPUT45), .B(KEYINPUT111), .Z(n461) );
  XNOR2_X1 U525 ( .A(n462), .B(n461), .ZN(n463) );
  NOR2_X1 U526 ( .A1(n463), .A2(n572), .ZN(n464) );
  NAND2_X1 U527 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U528 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U529 ( .A(n468), .B(KEYINPUT48), .ZN(n547) );
  NAND2_X1 U530 ( .A1(n469), .A2(n547), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n470), .B(KEYINPUT112), .ZN(n534) );
  NOR2_X1 U532 ( .A1(n555), .A2(n534), .ZN(n471) );
  XNOR2_X1 U533 ( .A(n471), .B(KEYINPUT113), .ZN(n472) );
  NOR2_X1 U534 ( .A1(n522), .A2(n472), .ZN(n473) );
  XNOR2_X1 U535 ( .A(KEYINPUT114), .B(n473), .ZN(n531) );
  NAND2_X1 U536 ( .A1(n531), .A2(n579), .ZN(n475) );
  NOR2_X1 U537 ( .A1(n563), .A2(n476), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n477), .B(KEYINPUT16), .ZN(n480) );
  INV_X1 U539 ( .A(n478), .ZN(n479) );
  NAND2_X1 U540 ( .A1(n480), .A2(n479), .ZN(n502) );
  NOR2_X1 U541 ( .A1(n481), .A2(n502), .ZN(n488) );
  NAND2_X1 U542 ( .A1(n488), .A2(n514), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n482), .B(KEYINPUT34), .ZN(n483) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n548), .A2(n488), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT94), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U548 ( .A1(n488), .A2(n518), .ZN(n485) );
  XNOR2_X1 U549 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(n487), .ZN(G1326GAT) );
  XOR2_X1 U551 ( .A(G22GAT), .B(KEYINPUT95), .Z(n490) );
  NAND2_X1 U552 ( .A1(n488), .A2(n522), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(G1327GAT) );
  NOR2_X1 U554 ( .A1(n497), .A2(n569), .ZN(n494) );
  XOR2_X1 U555 ( .A(KEYINPUT96), .B(KEYINPUT99), .Z(n492) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n491) );
  XNOR2_X1 U557 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NOR2_X1 U559 ( .A1(n495), .A2(n497), .ZN(n496) );
  XOR2_X1 U560 ( .A(G36GAT), .B(n496), .Z(G1329GAT) );
  NOR2_X1 U561 ( .A1(n498), .A2(n497), .ZN(n500) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(KEYINPUT101), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1331GAT) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U565 ( .A(KEYINPUT102), .B(n540), .ZN(n558) );
  NAND2_X1 U566 ( .A1(n558), .A2(n501), .ZN(n512) );
  NAND2_X1 U567 ( .A1(n514), .A2(n508), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  XOR2_X1 U569 ( .A(G64GAT), .B(KEYINPUT103), .Z(n506) );
  NAND2_X1 U570 ( .A1(n508), .A2(n548), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n518), .A2(n508), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U575 ( .A1(n508), .A2(n522), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NOR2_X1 U577 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n513), .B(KEYINPUT104), .ZN(n523) );
  NAND2_X1 U579 ( .A1(n523), .A2(n514), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U581 ( .A(G92GAT), .B(KEYINPUT105), .Z(n517) );
  NAND2_X1 U582 ( .A1(n523), .A2(n548), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n517), .B(n516), .ZN(G1337GAT) );
  NAND2_X1 U584 ( .A1(n523), .A2(n518), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n521) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(KEYINPUT107), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n521), .B(n520), .ZN(n526) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(KEYINPUT106), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(G1339GAT) );
  XOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT115), .Z(n528) );
  NAND2_X1 U593 ( .A1(n572), .A2(n531), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n530) );
  NAND2_X1 U596 ( .A1(n558), .A2(n531), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(G134GAT), .B(KEYINPUT51), .Z(n533) );
  NAND2_X1 U599 ( .A1(n563), .A2(n531), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(G1343GAT) );
  XNOR2_X1 U601 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n536) );
  NOR2_X1 U602 ( .A1(n534), .A2(n570), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n572), .A2(n545), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n538) );
  XNOR2_X1 U606 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n537) );
  XNOR2_X1 U607 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(n539), .Z(n542) );
  NAND2_X1 U609 ( .A1(n545), .A2(n540), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(G1345GAT) );
  XOR2_X1 U611 ( .A(G155GAT), .B(KEYINPUT119), .Z(n544) );
  NAND2_X1 U612 ( .A1(n545), .A2(n579), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n544), .B(n543), .ZN(G1346GAT) );
  NAND2_X1 U614 ( .A1(n545), .A2(n563), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n546), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n550) );
  AND2_X1 U617 ( .A1(n569), .A2(n551), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n293), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT121), .ZN(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT55), .B(n554), .ZN(n556) );
  NOR2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n564) );
  NAND2_X1 U622 ( .A1(n564), .A2(n572), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U624 ( .A1(n564), .A2(n558), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(n561), .ZN(G1349GAT) );
  NAND2_X1 U628 ( .A1(n564), .A2(n579), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT58), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G190GAT), .B(n566), .ZN(G1351GAT) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n567), .B(KEYINPUT122), .ZN(n568) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(n568), .Z(n574) );
  NAND2_X1 U636 ( .A1(n569), .A2(n293), .ZN(n571) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n584) );
  NAND2_X1 U638 ( .A1(n584), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n577) );
  NAND2_X1 U641 ( .A1(n584), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n578), .Z(G1353GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n581) );
  NAND2_X1 U645 ( .A1(n584), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n588) );
  XOR2_X1 U649 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n586) );
  NAND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(G1355GAT) );
endmodule

