//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT0), .B(G128), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT64), .B1(new_n189), .B2(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(KEYINPUT64), .A3(G143), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n188), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  AND2_X1   g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  AND3_X1   g011(.A1(new_n191), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n187), .B1(new_n194), .B2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n191), .A2(new_n196), .A3(new_n197), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n189), .A2(KEYINPUT64), .A3(G143), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(new_n191), .B2(new_n190), .ZN(new_n202));
  OAI211_X1 g016(.A(KEYINPUT66), .B(new_n200), .C1(new_n202), .C2(new_n188), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n206), .A2(new_n208), .A3(new_n212), .A4(new_n209), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n199), .A2(new_n203), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT64), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n216), .B1(new_n195), .B2(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n195), .A2(G146), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n193), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT1), .B1(new_n195), .B2(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G128), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n224), .A2(new_n191), .A3(new_n196), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n205), .A2(G137), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n207), .A2(G134), .ZN(new_n229));
  OAI21_X1  g043(.A(G131), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n213), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n215), .A2(KEYINPUT30), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT30), .ZN(new_n233));
  INV_X1    g047(.A(new_n188), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n198), .B1(new_n219), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n214), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n213), .A2(new_n230), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(new_n222), .B2(new_n226), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n233), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  OR2_X1    g053(.A1(KEYINPUT65), .A2(G116), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT65), .A2(G116), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(G119), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G116), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(G119), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT2), .B(G113), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n247), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n242), .A3(new_n245), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n232), .A2(new_n239), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n251), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n215), .A2(new_n253), .A3(new_n231), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n255));
  INV_X1    g069(.A(G953), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT68), .A2(G953), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT67), .A2(G237), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT67), .A2(G237), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n257), .B(new_n258), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G210), .ZN(new_n262));
  OR3_X1    g076(.A1(new_n261), .A2(KEYINPUT27), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT27), .B1(new_n261), .B2(new_n262), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(G101), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n263), .B2(new_n264), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n252), .A2(new_n254), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT31), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT31), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n252), .A2(new_n271), .A3(new_n254), .A4(new_n268), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n254), .A2(KEYINPUT28), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT28), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n215), .A2(new_n231), .A3(new_n274), .A4(new_n253), .ZN(new_n275));
  OR2_X1    g089(.A1(new_n236), .A2(new_n238), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n273), .A2(new_n275), .B1(new_n251), .B2(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n270), .B(new_n272), .C1(new_n268), .C2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(G472), .A2(G902), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT32), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT32), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n272), .B1(new_n277), .B2(new_n268), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n269), .A2(KEYINPUT31), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n282), .B(new_n279), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n252), .A2(new_n254), .ZN(new_n286));
  INV_X1    g100(.A(new_n268), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT29), .B1(new_n277), .B2(new_n268), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n286), .A2(KEYINPUT69), .A3(new_n287), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n253), .B1(new_n215), .B2(new_n231), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n273), .B2(new_n275), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT70), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n268), .A2(KEYINPUT29), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n296), .B1(new_n295), .B2(new_n297), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n299), .A2(G902), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n281), .A2(new_n285), .B1(new_n301), .B2(G472), .ZN(new_n302));
  XNOR2_X1  g116(.A(KEYINPUT24), .B(G110), .ZN(new_n303));
  INV_X1    g117(.A(G119), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G128), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n223), .A2(G119), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT72), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n305), .B2(new_n306), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n303), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n312), .B1(new_n304), .B2(G128), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n313), .A2(new_n305), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n315));
  INV_X1    g129(.A(G110), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n223), .A2(KEYINPUT23), .A3(G119), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n314), .A2(new_n315), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n313), .A2(new_n317), .A3(new_n316), .A4(new_n305), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT76), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n311), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n311), .A2(new_n318), .A3(KEYINPUT77), .A4(new_n320), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT74), .A2(G125), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(KEYINPUT74), .A2(G125), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(G140), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G125), .ZN(new_n330));
  OR3_X1    g144(.A1(new_n330), .A2(KEYINPUT73), .A3(G140), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT73), .B1(new_n330), .B2(G140), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n329), .A2(new_n331), .A3(KEYINPUT16), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n328), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT75), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n334), .A2(new_n335), .A3(new_n336), .A4(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n328), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(new_n326), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n336), .A2(new_n337), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT75), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n333), .A2(new_n338), .A3(new_n342), .A4(G146), .ZN(new_n343));
  XNOR2_X1  g157(.A(G125), .B(G140), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n344), .B(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n189), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n325), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n314), .A2(new_n317), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G110), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n305), .A2(new_n306), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT72), .ZN(new_n354));
  INV_X1    g168(.A(new_n303), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n308), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n333), .A2(new_n338), .A3(new_n342), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n189), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(new_n359), .B2(new_n343), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  XOR2_X1   g175(.A(KEYINPUT68), .B(G953), .Z(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(G221), .A3(G234), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT22), .B(G137), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n350), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n365), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n348), .B1(new_n323), .B2(new_n324), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(new_n360), .ZN(new_n369));
  INV_X1    g183(.A(G902), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n372), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n366), .A2(new_n369), .A3(new_n370), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G234), .ZN(new_n378));
  OAI21_X1  g192(.A(G217), .B1(new_n378), .B2(G902), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(KEYINPUT71), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(G902), .B1(new_n378), .B2(G217), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n366), .A2(new_n369), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT80), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n302), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G469), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n222), .B2(new_n226), .ZN(new_n390));
  INV_X1    g204(.A(G104), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT3), .B1(new_n391), .B2(G107), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n393));
  INV_X1    g207(.A(G107), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(G104), .ZN(new_n395));
  INV_X1    g209(.A(G101), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n391), .A2(G107), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n392), .A2(new_n395), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n391), .A2(G107), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n394), .A2(G104), .ZN(new_n400));
  OAI21_X1  g214(.A(G101), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  AOI22_X1  g217(.A1(new_n220), .A2(G128), .B1(new_n191), .B2(new_n196), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n398), .B(new_n401), .C1(new_n404), .C2(new_n225), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n390), .A2(new_n403), .B1(new_n389), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n214), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n392), .A2(new_n395), .A3(new_n397), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(G101), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(G101), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(KEYINPUT4), .A3(new_n398), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n199), .A2(new_n203), .A3(new_n410), .A4(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n406), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n362), .A2(G227), .ZN(new_n415));
  XOR2_X1   g229(.A(G110), .B(G140), .Z(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n222), .A2(new_n402), .A3(new_n226), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n405), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n420), .A2(KEYINPUT12), .A3(new_n214), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT12), .B1(new_n420), .B2(new_n214), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n414), .B(new_n418), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n390), .A2(new_n403), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n405), .A2(new_n389), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AND4_X1   g241(.A1(new_n199), .A2(new_n203), .A3(new_n410), .A4(new_n412), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n214), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n418), .B1(new_n429), .B2(new_n414), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n388), .B(new_n370), .C1(new_n424), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(G469), .A2(G902), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n414), .B1(new_n421), .B2(new_n422), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n417), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n429), .A2(new_n414), .A3(new_n418), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(G469), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n431), .A2(new_n432), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT9), .B(G234), .ZN(new_n438));
  OAI21_X1  g252(.A(G221), .B1(new_n438), .B2(G902), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(G214), .B1(G237), .B2(G902), .ZN(new_n441));
  OAI21_X1  g255(.A(G210), .B1(G237), .B2(G902), .ZN(new_n442));
  XOR2_X1   g256(.A(new_n442), .B(KEYINPUT85), .Z(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G110), .B(G122), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n445), .B(KEYINPUT82), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT8), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n445), .B(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT8), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n242), .A2(KEYINPUT5), .A3(new_n245), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT5), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n244), .A2(KEYINPUT81), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n244), .A2(new_n454), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT81), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n453), .A2(G113), .A3(new_n455), .A4(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n459), .A2(new_n250), .A3(new_n403), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n403), .B1(new_n459), .B2(new_n250), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n452), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT83), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n464), .B(new_n452), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n227), .A2(new_n340), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n235), .A2(new_n334), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G224), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(G953), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n469), .A2(KEYINPUT84), .A3(KEYINPUT7), .A4(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT84), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT7), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n474), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n334), .B1(new_n222), .B2(new_n226), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n194), .A2(new_n198), .A3(new_n340), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n472), .A2(KEYINPUT84), .A3(KEYINPUT7), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n251), .A2(new_n412), .A3(new_n410), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n459), .A2(new_n250), .A3(new_n403), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n446), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n473), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n370), .B1(new_n466), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n482), .A2(new_n483), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n449), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(KEYINPUT6), .A3(new_n484), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n469), .B(new_n472), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n487), .A2(new_n491), .A3(new_n449), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n444), .B1(new_n486), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n473), .A2(new_n481), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(new_n484), .A3(new_n463), .A4(new_n465), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n489), .A2(new_n490), .A3(new_n492), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n496), .A2(new_n370), .A3(new_n443), .A4(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n440), .A2(new_n441), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  XOR2_X1   g315(.A(KEYINPUT91), .B(G475), .Z(new_n502));
  XNOR2_X1  g316(.A(G113), .B(G122), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n391), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT86), .B(G143), .ZN(new_n506));
  INV_X1    g320(.A(G214), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n506), .B1(new_n261), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT67), .B(G237), .ZN(new_n509));
  OR2_X1    g323(.A1(KEYINPUT86), .A2(G143), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n362), .A2(G214), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n212), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n508), .A2(new_n511), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n513), .B1(new_n514), .B2(G131), .ZN(new_n515));
  AOI211_X1 g329(.A(KEYINPUT87), .B(new_n212), .C1(new_n508), .C2(new_n511), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n505), .B(new_n512), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(G131), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT87), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n514), .A2(new_n513), .A3(G131), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(KEYINPUT17), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n359), .A2(new_n343), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n517), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n329), .A2(new_n332), .A3(new_n331), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G146), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n347), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT18), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(new_n212), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n527), .B1(new_n514), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n518), .A2(new_n528), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n524), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT92), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n504), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n530), .A2(new_n531), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n515), .A2(new_n516), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n522), .B1(new_n537), .B2(KEYINPUT17), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n538), .B2(new_n517), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT92), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n524), .A2(new_n504), .A3(new_n532), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT89), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT89), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n524), .A2(new_n532), .A3(new_n544), .A4(new_n504), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n502), .B1(new_n547), .B2(new_n370), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n525), .A2(KEYINPUT19), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n344), .B(KEYINPUT78), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n549), .B1(new_n550), .B2(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n343), .B1(new_n551), .B2(G146), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT88), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT88), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n555), .B(new_n343), .C1(new_n551), .C2(G146), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n504), .B1(new_n557), .B2(new_n532), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n544), .B1(new_n539), .B2(new_n504), .ZN(new_n560));
  INV_X1    g374(.A(new_n545), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT90), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(G475), .A2(G902), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n558), .B1(new_n543), .B2(new_n545), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT90), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n564), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT20), .ZN(new_n569));
  INV_X1    g383(.A(new_n565), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n566), .A2(KEYINPUT20), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n548), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G217), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n438), .A2(new_n574), .A3(G953), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT95), .B1(new_n195), .B2(G128), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n578), .A2(new_n223), .A3(G143), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n195), .A2(G128), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n205), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(G134), .A3(new_n581), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT13), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n580), .A2(new_n585), .A3(G134), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n580), .A2(new_n585), .A3(G134), .A4(new_n581), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G122), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(G116), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT93), .ZN(new_n592));
  AND2_X1   g406(.A1(KEYINPUT65), .A2(G116), .ZN(new_n593));
  NOR2_X1   g407(.A1(KEYINPUT65), .A2(G116), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(KEYINPUT94), .B1(new_n595), .B2(G122), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT94), .ZN(new_n597));
  NOR4_X1   g411(.A1(new_n593), .A2(new_n594), .A3(new_n597), .A4(new_n590), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n592), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G107), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n394), .B(new_n592), .C1(new_n596), .C2(new_n598), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n589), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n580), .A2(G134), .A3(new_n581), .ZN(new_n603));
  AOI21_X1  g417(.A(G134), .B1(new_n580), .B2(new_n581), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(new_n601), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT14), .B1(new_n596), .B2(new_n598), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n240), .A2(G122), .A3(new_n241), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n597), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n595), .A2(KEYINPUT94), .A3(G122), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT14), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n607), .A2(new_n592), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n606), .B1(G107), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n576), .B1(new_n602), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(G107), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n601), .A3(new_n605), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n600), .A2(new_n601), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n587), .A3(new_n588), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n619), .A3(new_n575), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT96), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n615), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n617), .A2(new_n619), .A3(KEYINPUT96), .A4(new_n575), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n370), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(G478), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n625), .A2(KEYINPUT15), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n626), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n622), .A2(new_n370), .A3(new_n623), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n256), .A2(G952), .ZN(new_n631));
  INV_X1    g445(.A(G237), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n631), .B1(new_n378), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  AOI211_X1 g448(.A(new_n370), .B(new_n362), .C1(G234), .C2(G237), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT21), .B(G898), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT97), .B1(new_n573), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n571), .B1(new_n568), .B2(KEYINPUT20), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n641));
  INV_X1    g455(.A(new_n638), .ZN(new_n642));
  NOR4_X1   g456(.A1(new_n640), .A2(new_n641), .A3(new_n548), .A4(new_n642), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n387), .B(new_n501), .C1(new_n639), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(KEYINPUT98), .B(G101), .Z(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G3));
  NAND2_X1  g460(.A1(new_n622), .A2(new_n623), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n620), .A2(KEYINPUT99), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n615), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n649), .B1(new_n651), .B2(new_n648), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n625), .A2(G902), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n652), .A2(new_n653), .B1(new_n625), .B2(new_n624), .ZN(new_n654));
  AOI21_X1  g468(.A(KEYINPUT90), .B1(new_n546), .B2(new_n559), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n563), .B(new_n558), .C1(new_n543), .C2(new_n545), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n655), .A2(new_n656), .A3(new_n570), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT20), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n572), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n502), .ZN(new_n660));
  AOI22_X1  g474(.A1(new_n540), .A2(new_n535), .B1(new_n543), .B2(new_n545), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n660), .B1(new_n661), .B2(G902), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n654), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n499), .A2(new_n441), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n637), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n278), .A2(new_n370), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(G472), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n667), .A2(new_n280), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n382), .A2(new_n385), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n668), .A2(new_n669), .A3(new_n440), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n663), .A2(new_n665), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G104), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT100), .B(KEYINPUT34), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n662), .A2(new_n630), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n564), .A2(new_n658), .A3(new_n567), .A4(new_n565), .ZN(new_n677));
  AOI211_X1 g491(.A(new_n637), .B(new_n676), .C1(new_n569), .C2(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n664), .B1(new_n678), .B2(KEYINPUT101), .ZN(new_n679));
  INV_X1    g493(.A(new_n637), .ZN(new_n680));
  INV_X1    g494(.A(new_n676), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n655), .A2(new_n656), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n658), .B1(new_n682), .B2(new_n565), .ZN(new_n683));
  NOR4_X1   g497(.A1(new_n655), .A2(new_n656), .A3(KEYINPUT20), .A4(new_n570), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n680), .B(new_n681), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n675), .B1(new_n679), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n664), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n685), .B2(new_n686), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n676), .B1(new_n569), .B2(new_n677), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT101), .B1(new_n691), .B2(new_n680), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n690), .A2(new_n692), .A3(KEYINPUT102), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n670), .B1(new_n688), .B2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT35), .B(G107), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G9));
  INV_X1    g510(.A(new_n668), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT103), .ZN(new_n698));
  INV_X1    g512(.A(new_n376), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n371), .B2(new_n372), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n380), .B1(new_n700), .B2(new_n375), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n350), .A2(new_n361), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n367), .A2(KEYINPUT36), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n383), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n698), .B1(new_n701), .B2(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n382), .A2(KEYINPUT103), .A3(new_n705), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n697), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n501), .B(new_n710), .C1(new_n639), .C2(new_n643), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT37), .B(G110), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G12));
  NOR3_X1   g527(.A1(new_n709), .A2(new_n500), .A3(new_n302), .ZN(new_n714));
  INV_X1    g528(.A(new_n635), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n716));
  OR3_X1    g530(.A1(new_n715), .A2(new_n716), .A3(G900), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n716), .B1(new_n715), .B2(G900), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n633), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n714), .A2(new_n691), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G128), .ZN(G30));
  XNOR2_X1  g535(.A(new_n719), .B(KEYINPUT39), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n440), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(KEYINPUT40), .Z(new_n724));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n499), .B(KEYINPUT38), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n701), .A2(new_n706), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n727), .A2(new_n630), .A3(new_n441), .A4(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n724), .B2(new_n725), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n659), .A2(new_n662), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n215), .A2(new_n253), .A3(new_n231), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n287), .B1(new_n732), .B2(new_n294), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n733), .A2(KEYINPUT105), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(KEYINPUT105), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n734), .A2(new_n269), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(G472), .B1(new_n736), .B2(G902), .ZN(new_n737));
  INV_X1    g551(.A(new_n285), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n282), .B1(new_n278), .B2(new_n279), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT106), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n281), .A2(new_n285), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n737), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n726), .A2(new_n730), .A3(new_n731), .A4(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G143), .ZN(G45));
  NAND3_X1  g561(.A1(new_n663), .A2(new_n719), .A3(new_n714), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G146), .ZN(G48));
  INV_X1    g563(.A(new_n654), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n750), .B(new_n665), .C1(new_n640), .C2(new_n548), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n406), .A2(new_n407), .A3(new_n413), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n407), .B1(new_n406), .B2(new_n413), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n417), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n423), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n370), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(G469), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n431), .ZN(new_n758));
  INV_X1    g572(.A(new_n439), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n387), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT108), .B1(new_n751), .B2(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n738), .A2(new_n739), .ZN(new_n764));
  INV_X1    g578(.A(G472), .ZN(new_n765));
  INV_X1    g579(.A(new_n298), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n766), .A2(G902), .A3(new_n299), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n765), .B1(new_n767), .B2(new_n293), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n669), .B1(new_n764), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n760), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n663), .A2(new_n763), .A3(new_n665), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n762), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(KEYINPUT41), .B(G113), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G15));
  OAI21_X1  g589(.A(KEYINPUT102), .B1(new_n690), .B2(new_n692), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n691), .A2(KEYINPUT101), .A3(new_n680), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n687), .A2(new_n777), .A3(new_n675), .A4(new_n689), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n761), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n243), .ZN(G18));
  NAND3_X1  g594(.A1(new_n760), .A2(new_n441), .A3(new_n499), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n709), .A3(new_n302), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n639), .B2(new_n643), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G119), .ZN(G21));
  NAND2_X1  g598(.A1(new_n689), .A2(new_n630), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n785), .B1(new_n659), .B2(new_n662), .ZN(new_n786));
  INV_X1    g600(.A(new_n295), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n787), .A2(new_n287), .B1(new_n269), .B2(KEYINPUT31), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n272), .B1(new_n788), .B2(new_n789), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n279), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n667), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n793), .A2(new_n770), .A3(new_n386), .A4(new_n637), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n786), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G122), .ZN(G24));
  NAND2_X1  g610(.A1(new_n382), .A2(new_n705), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n792), .A2(new_n797), .A3(new_n667), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n798), .A2(new_n781), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n731), .A2(new_n750), .A3(new_n719), .A4(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G125), .ZN(G27));
  XOR2_X1   g615(.A(KEYINPUT112), .B(KEYINPUT42), .Z(new_n802));
  OAI211_X1 g616(.A(new_n750), .B(new_n719), .C1(new_n640), .C2(new_n548), .ZN(new_n803));
  INV_X1    g617(.A(new_n441), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n494), .B2(new_n498), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n436), .A2(new_n432), .ZN(new_n807));
  AOI211_X1 g621(.A(G469), .B(G902), .C1(new_n754), .C2(new_n423), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n431), .A2(KEYINPUT110), .A3(new_n432), .A4(new_n436), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n805), .A2(new_n809), .A3(new_n439), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n759), .B1(new_n437), .B2(new_n806), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(KEYINPUT111), .A3(new_n805), .A4(new_n810), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n387), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n802), .B1(new_n803), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n769), .B1(new_n813), .B2(new_n815), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT42), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT112), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n663), .A2(new_n819), .A3(new_n719), .A4(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(new_n212), .ZN(G33));
  NAND3_X1  g638(.A1(new_n819), .A2(new_n691), .A3(new_n719), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G134), .ZN(G36));
  XNOR2_X1  g640(.A(new_n731), .B(KEYINPUT113), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(KEYINPUT43), .A3(new_n750), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT43), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n829), .B1(new_n731), .B2(new_n654), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n697), .A2(new_n797), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT114), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT44), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n805), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  INV_X1    g653(.A(new_n722), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n434), .A2(new_n435), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT45), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n388), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n432), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT46), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n431), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n439), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI211_X1 g664(.A(new_n840), .B(new_n850), .C1(new_n834), .C2(new_n835), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n838), .A2(new_n839), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n852), .B(G137), .ZN(G39));
  XNOR2_X1  g667(.A(new_n850), .B(KEYINPUT47), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n302), .A2(new_n386), .A3(new_n805), .ZN(new_n855));
  OR3_X1    g669(.A1(new_n854), .A2(new_n803), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(G140), .ZN(G42));
  NOR2_X1   g671(.A1(new_n745), .A2(new_n386), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n759), .B(new_n804), .C1(new_n758), .C2(KEYINPUT49), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(KEYINPUT49), .B2(new_n758), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n860), .A2(new_n727), .A3(new_n654), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n827), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n798), .ZN(new_n863));
  INV_X1    g677(.A(new_n805), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n770), .A2(new_n633), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n831), .A2(KEYINPUT121), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT121), .B1(new_n831), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n858), .A2(new_n865), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n869), .A2(new_n731), .A3(new_n750), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n793), .A2(new_n386), .A3(new_n633), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n831), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n757), .A2(new_n759), .A3(new_n431), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n864), .B1(new_n854), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n870), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n727), .A2(new_n441), .A3(new_n770), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n831), .A2(new_n871), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT50), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n868), .B(new_n875), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT51), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n872), .A2(new_n689), .A3(new_n760), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n750), .B1(new_n640), .B2(new_n548), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n885), .B(new_n631), .C1(new_n886), .C2(new_n869), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n387), .B1(new_n866), .B2(new_n867), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n888), .A2(KEYINPUT48), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(KEYINPUT48), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n884), .A2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n771), .B1(new_n688), .B2(new_n693), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n798), .B1(new_n813), .B2(new_n815), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n663), .A2(new_n719), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n709), .A2(new_n302), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n569), .A2(new_n677), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n627), .A2(new_n629), .A3(new_n719), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n662), .A2(new_n440), .A3(new_n805), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n897), .A2(new_n898), .A3(new_n899), .A4(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n901), .B1(new_n569), .B2(new_n677), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n897), .B1(new_n904), .B2(new_n898), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n896), .B(new_n825), .C1(new_n903), .C2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n823), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n662), .B(new_n630), .C1(new_n683), .C2(new_n571), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n886), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n670), .A2(new_n665), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n909), .A2(new_n910), .B1(new_n786), .B2(new_n794), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n644), .A2(new_n911), .A3(new_n783), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n773), .A2(new_n711), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n894), .A2(new_n907), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n799), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n681), .B(new_n719), .C1(new_n683), .C2(new_n684), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n301), .A2(G472), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n742), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n501), .A2(new_n918), .A3(new_n707), .A4(new_n708), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n803), .A2(new_n915), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT52), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n728), .A2(new_n814), .A3(new_n719), .A4(new_n810), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n923), .B1(new_n741), .B2(new_n744), .ZN(new_n924));
  INV_X1    g738(.A(new_n785), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n731), .A3(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n921), .A2(new_n922), .A3(new_n748), .A4(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n748), .A2(new_n800), .A3(new_n926), .A4(new_n720), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT52), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n893), .B1(new_n914), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n644), .A2(new_n911), .A3(new_n783), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n773), .A2(new_n711), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n779), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n920), .A2(KEYINPUT52), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n927), .A2(new_n929), .A3(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n934), .A2(new_n936), .A3(KEYINPUT53), .A4(new_n907), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT54), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n931), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT119), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT119), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n931), .A2(new_n937), .A3(new_n941), .A4(new_n938), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n927), .A2(new_n929), .A3(new_n935), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n893), .B1(new_n914), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT117), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT117), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n946), .B(new_n893), .C1(new_n914), .C2(new_n943), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n928), .B(new_n922), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n932), .A2(new_n933), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n948), .A2(new_n949), .A3(new_n894), .A4(new_n907), .ZN(new_n950));
  OAI21_X1  g764(.A(KEYINPUT118), .B1(new_n950), .B2(new_n893), .ZN(new_n951));
  AND4_X1   g765(.A1(new_n894), .A2(new_n907), .A3(new_n912), .A4(new_n913), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT118), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT53), .A4(new_n948), .ZN(new_n954));
  AOI22_X1  g768(.A1(new_n945), .A2(new_n947), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n940), .B(new_n942), .C1(new_n955), .C2(new_n938), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n883), .A2(KEYINPUT51), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n892), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g772(.A1(G952), .A2(G953), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n862), .B1(new_n958), .B2(new_n959), .ZN(G75));
  NOR2_X1   g774(.A1(new_n362), .A2(G952), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n370), .B1(new_n931), .B2(new_n937), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT56), .B1(new_n963), .B2(new_n443), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n489), .A2(new_n492), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(new_n490), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT55), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n962), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n964), .B2(new_n967), .ZN(G51));
  NAND2_X1  g783(.A1(new_n931), .A2(new_n937), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(KEYINPUT54), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n939), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n432), .B(KEYINPUT57), .Z(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n755), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n963), .B(new_n843), .C1(new_n842), .C2(new_n841), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n961), .B1(new_n975), .B2(new_n976), .ZN(G54));
  NAND3_X1  g791(.A1(new_n963), .A2(KEYINPUT58), .A3(G475), .ZN(new_n978));
  INV_X1    g792(.A(new_n682), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n980), .A2(new_n981), .A3(new_n961), .ZN(G60));
  NAND2_X1  g796(.A1(G478), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT59), .Z(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n652), .B1(new_n956), .B2(new_n985), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n652), .A2(new_n985), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n961), .B1(new_n972), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT122), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT122), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n945), .A2(new_n947), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n951), .A2(new_n954), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(KEYINPUT54), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n940), .A2(new_n942), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n984), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g811(.A(new_n991), .B(new_n988), .C1(new_n997), .C2(new_n652), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n990), .A2(new_n998), .ZN(G63));
  INV_X1    g813(.A(KEYINPUT61), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(KEYINPUT124), .ZN(new_n1001));
  XNOR2_X1  g815(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n574), .A2(new_n370), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n970), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n366), .A2(new_n369), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n961), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n970), .A2(new_n704), .A3(new_n1004), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1001), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1000), .A2(KEYINPUT124), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1009), .B(new_n1010), .Z(G66));
  OAI21_X1  g825(.A(G953), .B1(new_n636), .B2(new_n470), .ZN(new_n1012));
  INV_X1    g826(.A(new_n362), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1012), .B1(new_n934), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n965), .B1(G898), .B2(new_n362), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT125), .Z(new_n1016));
  XNOR2_X1  g830(.A(new_n1014), .B(new_n1016), .ZN(G69));
  INV_X1    g831(.A(new_n909), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n387), .A2(new_n440), .A3(new_n722), .A4(new_n805), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n921), .A2(new_n748), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n746), .ZN(new_n1021));
  OAI221_X1 g835(.A(new_n856), .B1(new_n1018), .B2(new_n1019), .C1(new_n1021), .C2(KEYINPUT62), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(KEYINPUT62), .ZN(new_n1023));
  OR2_X1    g837(.A1(new_n1023), .A2(KEYINPUT127), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(KEYINPUT127), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n852), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n232), .A2(new_n239), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT126), .Z(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(new_n551), .Z(new_n1030));
  NOR3_X1   g844(.A1(new_n1027), .A2(new_n1013), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(new_n1030), .ZN(new_n1032));
  INV_X1    g846(.A(new_n850), .ZN(new_n1033));
  NAND4_X1  g847(.A1(new_n1033), .A2(new_n387), .A3(new_n722), .A4(new_n786), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n856), .A2(new_n825), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1020), .ZN(new_n1036));
  NOR3_X1   g850(.A1(new_n1035), .A2(new_n823), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n852), .A2(new_n362), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1013), .A2(G900), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1032), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n362), .B1(G227), .B2(G900), .ZN(new_n1041));
  NOR3_X1   g855(.A1(new_n1031), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1043));
  NAND2_X1  g857(.A1(G227), .A2(G900), .ZN(new_n1044));
  AND4_X1   g858(.A1(new_n1013), .A2(new_n1043), .A3(new_n1044), .A4(new_n1030), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1042), .A2(new_n1045), .ZN(G72));
  NAND2_X1  g860(.A1(G472), .A2(G902), .ZN(new_n1047));
  XOR2_X1   g861(.A(new_n1047), .B(KEYINPUT63), .Z(new_n1048));
  NAND2_X1  g862(.A1(new_n852), .A2(new_n1026), .ZN(new_n1049));
  INV_X1    g863(.A(new_n934), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n287), .B1(new_n252), .B2(new_n254), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1053), .A2(new_n962), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n290), .A2(new_n269), .A3(new_n292), .ZN(new_n1055));
  AND3_X1   g869(.A1(new_n994), .A2(new_n1048), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g870(.A1(new_n852), .A2(new_n934), .A3(new_n1037), .ZN(new_n1057));
  AOI211_X1 g871(.A(new_n286), .B(new_n268), .C1(new_n1057), .C2(new_n1048), .ZN(new_n1058));
  NOR3_X1   g872(.A1(new_n1054), .A2(new_n1056), .A3(new_n1058), .ZN(G57));
endmodule


