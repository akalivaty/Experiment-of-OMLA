//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n562,
    new_n563, new_n564, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n592, new_n593, new_n596, new_n598,
    new_n599, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT65), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT66), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(KEYINPUT68), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n462), .A2(G2105), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n466), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n473), .A2(new_n474), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n468), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n466), .A2(G136), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT69), .Z(new_n483));
  AOI21_X1  g058(.A(new_n469), .B1(new_n463), .B2(new_n465), .ZN(new_n484));
  AOI211_X1 g059(.A(new_n481), .B(new_n483), .C1(G124), .C2(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(new_n484), .A2(G126), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n489), .A2(KEYINPUT70), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(new_n469), .A3(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT71), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n495), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n497), .A2(new_n470), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT3), .B1(new_n464), .B2(G2104), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n469), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n489), .A2(KEYINPUT70), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n490), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT5), .B(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n510), .A2(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT72), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n516), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n515), .A2(new_n520), .ZN(G166));
  INV_X1    g096(.A(new_n513), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n511), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n523), .B(new_n524), .C1(new_n528), .C2(KEYINPUT73), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n529), .A2(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n511), .A2(new_n533), .B1(new_n513), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n516), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(G171));
  AOI22_X1  g113(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n516), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n522), .A2(G43), .ZN(new_n541));
  INV_X1    g116(.A(new_n511), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G81), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND3_X1  g125(.A1(new_n522), .A2(KEYINPUT74), .A3(G53), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n552));
  AOI21_X1  g127(.A(KEYINPUT74), .B1(new_n522), .B2(G53), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n552), .B(new_n553), .Z(new_n554));
  AOI22_X1  g129(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(KEYINPUT75), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n516), .B1(new_n555), .B2(KEYINPUT75), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n556), .A2(new_n557), .B1(G91), .B2(new_n542), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G299));
  INV_X1    g134(.A(G171), .ZN(G301));
  INV_X1    g135(.A(G166), .ZN(G303));
  NAND2_X1  g136(.A1(new_n542), .A2(G87), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n522), .A2(G49), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(G288));
  AOI22_X1  g140(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(new_n516), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(KEYINPUT76), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(KEYINPUT76), .ZN(new_n569));
  AOI22_X1  g144(.A1(G86), .A2(new_n542), .B1(new_n522), .B2(G48), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G305));
  AOI22_X1  g146(.A1(G85), .A2(new_n542), .B1(new_n522), .B2(G47), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n516), .B2(new_n573), .ZN(G290));
  NAND2_X1  g149(.A1(G301), .A2(G868), .ZN(new_n575));
  AND3_X1   g150(.A1(new_n510), .A2(new_n509), .A3(G92), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT10), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(G79), .A2(G543), .ZN(new_n581));
  XOR2_X1   g156(.A(KEYINPUT5), .B(G543), .Z(new_n582));
  INV_X1    g157(.A(G66), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G651), .B1(new_n522), .B2(G54), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  OR2_X1    g161(.A1(new_n578), .A2(new_n579), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n575), .B1(new_n589), .B2(G868), .ZN(G284));
  OAI21_X1  g165(.A(new_n575), .B1(new_n589), .B2(G868), .ZN(G321));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(G299), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(new_n592), .B2(G168), .ZN(G297));
  OAI21_X1  g169(.A(new_n593), .B1(new_n592), .B2(G168), .ZN(G280));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n589), .B1(new_n596), .B2(G860), .ZN(G148));
  NAND2_X1  g172(.A1(new_n589), .A2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G868), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g175(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g176(.A1(new_n470), .A2(new_n467), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT12), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT13), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(G2100), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n466), .A2(G135), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n484), .A2(G123), .ZN(new_n607));
  OR2_X1    g182(.A1(G99), .A2(G2105), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n608), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(G2096), .Z(new_n611));
  NAND2_X1  g186(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT78), .ZN(G156));
  XNOR2_X1  g188(.A(G2427), .B(G2438), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2430), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT15), .B(G2435), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n616), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n617), .A2(KEYINPUT14), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(G1341), .B(G1348), .Z(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n619), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G2451), .B(G2454), .Z(new_n624));
  XNOR2_X1  g199(.A(G2443), .B(G2446), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n623), .A2(new_n626), .ZN(new_n628));
  AND3_X1   g203(.A1(new_n627), .A2(G14), .A3(new_n628), .ZN(G401));
  XNOR2_X1  g204(.A(G2067), .B(G2678), .ZN(new_n630));
  NOR2_X1   g205(.A1(G2072), .A2(G2078), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n442), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n633), .B2(KEYINPUT80), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(KEYINPUT80), .B2(new_n633), .ZN(new_n635));
  XOR2_X1   g210(.A(G2084), .B(G2090), .Z(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n632), .B(KEYINPUT17), .ZN(new_n638));
  INV_X1    g213(.A(new_n630), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n635), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n630), .A3(new_n636), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT18), .Z(new_n642));
  NAND3_X1  g217(.A1(new_n638), .A2(new_n639), .A3(new_n636), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n640), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT81), .ZN(new_n645));
  XOR2_X1   g220(.A(G2096), .B(G2100), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(G227));
  XOR2_X1   g222(.A(G1971), .B(G1976), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT19), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1956), .B(G2474), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1961), .B(G1966), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n649), .A2(new_n654), .A3(new_n652), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n649), .A2(new_n654), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n657));
  AOI211_X1 g232(.A(new_n653), .B(new_n655), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n656), .B2(new_n657), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1991), .B(G1996), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1981), .B(G1986), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G229));
  INV_X1    g241(.A(G305), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(G16), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(G6), .B2(G16), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT32), .B(G1981), .Z(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G22), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n674), .B1(G166), .B2(new_n673), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(G1971), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(G23), .ZN(new_n677));
  INV_X1    g252(.A(G288), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n677), .B1(new_n678), .B2(new_n673), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT33), .B(G1976), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND4_X1  g256(.A1(new_n671), .A2(new_n672), .A3(new_n676), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT85), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT84), .B(KEYINPUT34), .Z(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  MUX2_X1   g261(.A(G24), .B(G290), .S(G16), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1986), .ZN(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G25), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n466), .A2(G131), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n484), .A2(G119), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n469), .A2(G107), .ZN(new_n693));
  OAI21_X1  g268(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n691), .B(new_n692), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT83), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n690), .B1(new_n696), .B2(new_n689), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT35), .B(G1991), .Z(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n688), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n685), .A2(new_n686), .A3(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT36), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n689), .A2(G26), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT28), .Z(new_n706));
  NAND2_X1  g281(.A1(new_n466), .A2(G140), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT86), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n709));
  INV_X1    g284(.A(G116), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(G2105), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT87), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT87), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n712), .A2(new_n713), .B1(G128), .B2(new_n484), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n706), .B1(new_n715), .B2(G29), .ZN(new_n716));
  INV_X1    g291(.A(G2067), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT88), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT25), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n466), .A2(G139), .ZN(new_n722));
  AOI22_X1  g297(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n721), .B(new_n722), .C1(new_n469), .C2(new_n723), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT89), .Z(new_n725));
  MUX2_X1   g300(.A(G33), .B(new_n725), .S(G29), .Z(new_n726));
  XOR2_X1   g301(.A(KEYINPUT90), .B(G2072), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n673), .A2(G4), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(new_n589), .B2(new_n673), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n718), .B(new_n728), .C1(G1348), .C2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n730), .A2(G1348), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(G28), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n689), .B1(new_n733), .B2(G28), .ZN(new_n735));
  NOR2_X1   g310(.A1(KEYINPUT31), .A2(G11), .ZN(new_n736));
  AND2_X1   g311(.A1(KEYINPUT31), .A2(G11), .ZN(new_n737));
  OAI22_X1  g312(.A1(new_n734), .A2(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G19), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n545), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT92), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n610), .A2(new_n689), .ZN(new_n742));
  OAI22_X1  g317(.A1(new_n740), .A2(G1341), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n738), .B(new_n743), .C1(new_n741), .C2(new_n742), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT91), .B(KEYINPUT26), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G105), .B2(new_n467), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n466), .A2(G141), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n484), .A2(G129), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  MUX2_X1   g326(.A(G32), .B(new_n751), .S(G29), .Z(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT27), .B(G1996), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G2078), .ZN(new_n755));
  NOR2_X1   g330(.A1(G164), .A2(new_n689), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G27), .B2(new_n689), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n744), .B(new_n754), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n732), .B(new_n758), .C1(new_n755), .C2(new_n757), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G35), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G162), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2090), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n673), .A2(G21), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G168), .B2(new_n673), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(G1966), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT93), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n740), .A2(G1341), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  NOR2_X1   g345(.A1(G171), .A2(new_n673), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(G5), .B2(new_n673), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n769), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n770), .B2(new_n772), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT24), .ZN(new_n775));
  INV_X1    g350(.A(G34), .ZN(new_n776));
  AOI21_X1  g351(.A(G29), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n775), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G160), .B2(new_n689), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(G2084), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n765), .A2(G1966), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(G2084), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n774), .A2(new_n780), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n673), .A2(G20), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT23), .Z(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G299), .B2(G16), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT94), .B(G1956), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n731), .A2(new_n759), .A3(new_n768), .A4(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n704), .A2(new_n790), .ZN(G311));
  INV_X1    g366(.A(G311), .ZN(G150));
  NAND2_X1  g367(.A1(new_n589), .A2(G559), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT96), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT38), .ZN(new_n795));
  NAND2_X1  g370(.A1(G80), .A2(G543), .ZN(new_n796));
  INV_X1    g371(.A(G67), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n582), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT95), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n516), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n799), .B2(new_n798), .ZN(new_n801));
  AOI22_X1  g376(.A1(G93), .A2(new_n542), .B1(new_n522), .B2(G55), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(new_n544), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n795), .B(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT39), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT97), .ZN(new_n808));
  AOI21_X1  g383(.A(G860), .B1(new_n805), .B2(new_n806), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n803), .A2(G860), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT37), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(G145));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n505), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n489), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n500), .A2(new_n504), .A3(KEYINPUT98), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(new_n715), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n725), .B(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(new_n751), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n484), .A2(G130), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n469), .A2(G118), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G142), .B2(new_n466), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(new_n603), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n695), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n821), .A2(new_n828), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n477), .B(new_n610), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G162), .ZN(new_n833));
  AOI21_X1  g408(.A(G37), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n830), .A2(KEYINPUT99), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(KEYINPUT99), .ZN(new_n836));
  INV_X1    g411(.A(new_n833), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n836), .A2(new_n829), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n834), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g415(.A(new_n803), .B(new_n545), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n598), .B(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(G299), .A2(new_n588), .ZN(new_n843));
  NAND2_X1  g418(.A1(G299), .A2(new_n588), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT41), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n843), .A2(KEYINPUT41), .A3(new_n844), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n842), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n846), .A2(KEYINPUT100), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n847), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(KEYINPUT42), .ZN(new_n854));
  XOR2_X1   g429(.A(G305), .B(G290), .Z(new_n855));
  XNOR2_X1  g430(.A(G288), .B(G166), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n855), .B(new_n856), .Z(new_n857));
  INV_X1    g432(.A(KEYINPUT42), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n847), .B(new_n858), .C1(new_n851), .C2(new_n852), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n854), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n857), .B1(new_n854), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(G868), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n803), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(G868), .B2(new_n863), .ZN(G295));
  OAI21_X1  g439(.A(new_n862), .B1(G868), .B2(new_n863), .ZN(G331));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n841), .A2(G301), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n804), .A2(G171), .ZN(new_n868));
  AOI21_X1  g443(.A(G168), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n867), .A3(G168), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n849), .A2(new_n870), .A3(new_n850), .A4(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT102), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n871), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n844), .B(new_n843), .C1(new_n875), .C2(new_n869), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n872), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(new_n857), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT103), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n874), .A2(new_n877), .A3(new_n880), .A4(new_n857), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n857), .ZN(new_n883));
  AND3_X1   g458(.A1(new_n872), .A2(new_n876), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(G37), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(KEYINPUT43), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n883), .B1(new_n872), .B2(new_n876), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(G37), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n884), .B1(new_n890), .B2(KEYINPUT101), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n889), .B2(G37), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n888), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n866), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n888), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(KEYINPUT44), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n886), .A2(KEYINPUT43), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n888), .B1(new_n882), .B2(new_n885), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n902), .A2(new_n898), .A3(KEYINPUT104), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n895), .B1(new_n901), .B2(new_n903), .ZN(G397));
  OAI211_X1 g479(.A(G40), .B(new_n468), .C1(new_n475), .C2(new_n476), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n489), .B1(new_n505), .B2(new_n814), .ZN(new_n908));
  AOI211_X1 g483(.A(new_n907), .B(G1384), .C1(new_n908), .C2(new_n817), .ZN(new_n909));
  INV_X1    g484(.A(G1384), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT108), .B1(new_n818), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT50), .ZN(new_n913));
  OAI211_X1 g488(.A(KEYINPUT113), .B(new_n906), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT113), .ZN(new_n915));
  AOI22_X1  g490(.A1(new_n496), .A2(new_n499), .B1(new_n503), .B2(KEYINPUT4), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n816), .B1(new_n916), .B2(KEYINPUT98), .ZN(new_n917));
  INV_X1    g492(.A(new_n817), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n910), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n907), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n818), .A2(KEYINPUT108), .A3(new_n910), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n913), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n915), .B1(new_n922), .B2(new_n905), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n507), .A2(new_n910), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n924), .A2(KEYINPUT50), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n914), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G1956), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(G299), .B(KEYINPUT57), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n924), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n818), .A2(KEYINPUT45), .A3(new_n910), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n933), .A2(new_n934), .A3(new_n906), .ZN(new_n935));
  XNOR2_X1  g510(.A(KEYINPUT56), .B(G2072), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n929), .A2(new_n931), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n931), .B1(new_n929), .B2(new_n938), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n920), .A2(new_n913), .A3(new_n921), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n905), .B1(new_n924), .B2(KEYINPUT50), .ZN(new_n942));
  AOI21_X1  g517(.A(G1348), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n920), .A2(new_n906), .A3(new_n921), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n944), .A2(G2067), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n946), .A2(new_n588), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n939), .B1(new_n940), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n920), .A2(new_n921), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n905), .B1(new_n949), .B2(KEYINPUT50), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n925), .B1(new_n950), .B2(KEYINPUT113), .ZN(new_n951));
  AOI21_X1  g526(.A(G1956), .B1(new_n951), .B2(new_n923), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n930), .B1(new_n952), .B2(new_n937), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(KEYINPUT61), .A3(new_n939), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT117), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n953), .A2(KEYINPUT117), .A3(new_n939), .A4(KEYINPUT61), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT60), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n943), .A2(new_n945), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT119), .B1(new_n960), .B2(new_n588), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n941), .A2(new_n942), .ZN(new_n962));
  INV_X1    g537(.A(G1348), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n912), .A2(new_n717), .A3(new_n906), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(KEYINPUT60), .A3(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT119), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n967), .A3(new_n589), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n961), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT118), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n960), .A2(new_n970), .A3(new_n588), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n964), .A2(KEYINPUT60), .A3(new_n588), .A4(new_n965), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT118), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OAI22_X1  g549(.A1(new_n969), .A2(new_n974), .B1(KEYINPUT60), .B2(new_n946), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT61), .ZN(new_n976));
  AOI211_X1 g551(.A(new_n930), .B(new_n937), .C1(new_n927), .C2(new_n928), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n976), .B1(new_n940), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  XOR2_X1   g554(.A(KEYINPUT58), .B(G1341), .Z(new_n980));
  AOI22_X1  g555(.A1(new_n935), .A2(new_n979), .B1(new_n944), .B2(new_n980), .ZN(new_n981));
  OAI22_X1  g556(.A1(new_n981), .A2(new_n544), .B1(KEYINPUT115), .B2(KEYINPUT59), .ZN(new_n982));
  NAND2_X1  g557(.A1(KEYINPUT115), .A2(KEYINPUT59), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT116), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n982), .B(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n975), .A2(new_n978), .A3(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n948), .B1(new_n958), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(G286), .A2(G8), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT120), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT45), .B1(new_n920), .B2(new_n921), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n991), .B2(new_n905), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n932), .B1(new_n909), .B2(new_n911), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n993), .A2(KEYINPUT114), .A3(new_n906), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n910), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n992), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1966), .ZN(new_n997));
  INV_X1    g572(.A(G2084), .ZN(new_n998));
  INV_X1    g573(.A(new_n962), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n996), .A2(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G8), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n989), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n996), .A2(new_n997), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n999), .A2(new_n998), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n989), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT51), .B1(new_n1006), .B2(KEYINPUT121), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1002), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G303), .A2(G8), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n933), .A2(new_n934), .A3(new_n906), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT107), .B(G1971), .Z(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1017), .B1(new_n927), .B2(G2090), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1014), .B1(new_n1018), .B2(G8), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n678), .A2(G1976), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n944), .A2(KEYINPUT110), .A3(G8), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT110), .B1(new_n944), .B2(G8), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT52), .ZN(new_n1024));
  AND2_X1   g599(.A1(G305), .A2(G1981), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT111), .B(G1981), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1025), .B1(new_n667), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1028), .B2(KEYINPUT49), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n1030));
  OAI221_X1 g605(.A(new_n1029), .B1(new_n1027), .B2(new_n1030), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1017), .B1(new_n962), .B2(G2090), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1032), .A2(G8), .A3(new_n1014), .ZN(new_n1033));
  INV_X1    g608(.A(G1976), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT52), .B1(G288), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1020), .B(new_n1035), .C1(new_n1021), .C2(new_n1022), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1024), .A2(new_n1031), .A3(new_n1033), .A4(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1019), .A2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n989), .B(new_n1008), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n933), .A2(new_n934), .A3(new_n755), .A4(new_n906), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n962), .A2(new_n770), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n919), .A2(new_n932), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1041), .A2(G2078), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(G40), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n473), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1043), .A2(new_n468), .A3(new_n934), .A4(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1042), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G171), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n992), .A2(new_n994), .A3(new_n1044), .A4(new_n995), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1042), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1049), .B(KEYINPUT54), .C1(G171), .C2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1010), .A2(new_n1038), .A3(new_n1039), .A4(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT122), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1054), .B1(new_n1051), .B2(G171), .ZN(new_n1055));
  AOI211_X1 g630(.A(KEYINPUT122), .B(G301), .C1(new_n1050), .C2(new_n1042), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1042), .A2(G301), .A3(new_n1047), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT123), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT54), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n987), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(G288), .A2(G1976), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1031), .A2(new_n1063), .B1(new_n667), .B2(new_n1026), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1024), .A2(new_n1031), .A3(new_n1036), .ZN(new_n1067));
  OAI22_X1  g642(.A1(new_n1064), .A2(new_n1066), .B1(new_n1067), .B2(new_n1033), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1000), .A2(new_n1001), .A3(G286), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1038), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT63), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1037), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1032), .A2(G8), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1071), .B1(new_n1074), .B2(new_n1013), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1069), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1068), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(KEYINPUT62), .B1(new_n1010), .B2(new_n1039), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1006), .B1(new_n1005), .B2(G8), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1009), .B1(new_n1000), .B2(new_n989), .ZN(new_n1081));
  OAI211_X1 g656(.A(KEYINPUT62), .B(new_n1039), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1057), .A2(new_n1019), .A3(new_n1037), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1079), .A2(KEYINPUT124), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT124), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1057), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1082), .A2(new_n1086), .A3(new_n1038), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1087), .B2(new_n1078), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1062), .A2(new_n1077), .A3(new_n1084), .A4(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1043), .A2(new_n905), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n715), .A2(G2067), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n708), .A2(new_n717), .A3(new_n714), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1093), .B(KEYINPUT106), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n751), .B(new_n979), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n695), .B(new_n699), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g673(.A1(G290), .A2(G1986), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1099), .A2(KEYINPUT105), .ZN(new_n1100));
  NAND2_X1  g675(.A1(G290), .A2(G1986), .ZN(new_n1101));
  XOR2_X1   g676(.A(new_n1100), .B(new_n1101), .Z(new_n1102));
  OAI21_X1  g677(.A(new_n1090), .B1(new_n1098), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1089), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1090), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1096), .A2(new_n696), .A3(new_n699), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(new_n1092), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT125), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT46), .B1(new_n1090), .B2(new_n979), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n751), .B1(KEYINPUT46), .B2(new_n979), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1094), .A2(new_n1113), .ZN(new_n1114));
  OAI22_X1  g689(.A1(new_n1111), .A2(new_n1112), .B1(new_n1114), .B2(new_n1105), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT47), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1098), .A2(new_n1090), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1090), .A2(new_n1099), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT48), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1118), .A2(KEYINPUT48), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1117), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1108), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1104), .A2(new_n1122), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g698(.A1(new_n887), .A2(new_n894), .ZN(new_n1125));
  NOR3_X1   g699(.A1(G227), .A2(G401), .A3(new_n459), .ZN(new_n1126));
  OR2_X1    g700(.A1(new_n1126), .A2(KEYINPUT127), .ZN(new_n1127));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT127), .ZN(new_n1128));
  NAND4_X1  g702(.A1(new_n839), .A2(new_n665), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  NOR2_X1   g703(.A1(new_n1125), .A2(new_n1129), .ZN(G308));
  OR2_X1    g704(.A1(new_n1125), .A2(new_n1129), .ZN(G225));
endmodule


