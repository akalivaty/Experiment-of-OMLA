

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n739), .A2(n738), .ZN(n741) );
  AND2_X1 U549 ( .A1(n734), .A2(G1996), .ZN(n705) );
  NOR2_X1 U550 ( .A1(n855), .A2(n708), .ZN(n710) );
  INV_X1 U551 ( .A(KEYINPUT28), .ZN(n727) );
  INV_X1 U552 ( .A(KEYINPUT96), .ZN(n740) );
  NOR2_X1 U553 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U554 ( .A1(n701), .A2(n700), .ZN(n712) );
  BUF_X1 U555 ( .A(n712), .Z(n761) );
  NOR2_X1 U556 ( .A1(G2105), .A2(G2104), .ZN(n513) );
  NOR2_X1 U557 ( .A1(G543), .A2(G651), .ZN(n630) );
  NAND2_X1 U558 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U559 ( .A(n522), .B(KEYINPUT65), .ZN(G160) );
  AND2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n993) );
  NAND2_X1 U561 ( .A1(n993), .A2(G113), .ZN(n521) );
  XOR2_X2 U562 ( .A(KEYINPUT17), .B(n513), .Z(n998) );
  NAND2_X1 U563 ( .A1(G137), .A2(n998), .ZN(n515) );
  INV_X1 U564 ( .A(G2105), .ZN(n516) );
  NOR2_X1 U565 ( .A1(G2104), .A2(n516), .ZN(n994) );
  NAND2_X1 U566 ( .A1(G125), .A2(n994), .ZN(n514) );
  NAND2_X1 U567 ( .A1(n515), .A2(n514), .ZN(n519) );
  AND2_X1 U568 ( .A1(n516), .A2(G2104), .ZN(n997) );
  NAND2_X1 U569 ( .A1(G101), .A2(n997), .ZN(n517) );
  XNOR2_X1 U570 ( .A(KEYINPUT23), .B(n517), .ZN(n518) );
  NOR2_X1 U571 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U572 ( .A1(G85), .A2(n630), .ZN(n524) );
  XOR2_X1 U573 ( .A(KEYINPUT0), .B(G543), .Z(n639) );
  INV_X1 U574 ( .A(G651), .ZN(n525) );
  NOR2_X1 U575 ( .A1(n639), .A2(n525), .ZN(n628) );
  NAND2_X1 U576 ( .A1(G72), .A2(n628), .ZN(n523) );
  NAND2_X1 U577 ( .A1(n524), .A2(n523), .ZN(n531) );
  NOR2_X1 U578 ( .A1(G543), .A2(n525), .ZN(n526) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n526), .Z(n643) );
  NAND2_X1 U580 ( .A1(G60), .A2(n643), .ZN(n529) );
  NOR2_X1 U581 ( .A1(n639), .A2(G651), .ZN(n527) );
  XNOR2_X1 U582 ( .A(KEYINPUT64), .B(n527), .ZN(n644) );
  NAND2_X1 U583 ( .A1(G47), .A2(n644), .ZN(n528) );
  NAND2_X1 U584 ( .A1(n529), .A2(n528), .ZN(n530) );
  OR2_X1 U585 ( .A1(n531), .A2(n530), .ZN(G290) );
  XOR2_X1 U586 ( .A(G2443), .B(G2446), .Z(n533) );
  XNOR2_X1 U587 ( .A(G2427), .B(G2451), .ZN(n532) );
  XNOR2_X1 U588 ( .A(n533), .B(n532), .ZN(n539) );
  XOR2_X1 U589 ( .A(G2430), .B(G2454), .Z(n535) );
  XNOR2_X1 U590 ( .A(G1348), .B(G1341), .ZN(n534) );
  XNOR2_X1 U591 ( .A(n535), .B(n534), .ZN(n537) );
  XOR2_X1 U592 ( .A(G2435), .B(G2438), .Z(n536) );
  XNOR2_X1 U593 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U594 ( .A(n539), .B(n538), .Z(n540) );
  AND2_X1 U595 ( .A1(G14), .A2(n540), .ZN(G401) );
  AND2_X1 U596 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U597 ( .A1(G123), .A2(n994), .ZN(n541) );
  XNOR2_X1 U598 ( .A(n541), .B(KEYINPUT18), .ZN(n549) );
  NAND2_X1 U599 ( .A1(G111), .A2(n993), .ZN(n542) );
  XNOR2_X1 U600 ( .A(n542), .B(KEYINPUT76), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n997), .A2(G99), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n547) );
  NAND2_X1 U603 ( .A1(G135), .A2(n998), .ZN(n545) );
  XNOR2_X1 U604 ( .A(KEYINPUT75), .B(n545), .ZN(n546) );
  NOR2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n982) );
  XNOR2_X1 U607 ( .A(G2096), .B(n982), .ZN(n550) );
  OR2_X1 U608 ( .A1(G2100), .A2(n550), .ZN(G156) );
  INV_X1 U609 ( .A(G82), .ZN(G220) );
  INV_X1 U610 ( .A(G108), .ZN(G238) );
  NAND2_X1 U611 ( .A1(G90), .A2(n630), .ZN(n552) );
  NAND2_X1 U612 ( .A1(G77), .A2(n628), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U614 ( .A(KEYINPUT9), .B(n553), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n644), .A2(G52), .ZN(n555) );
  NAND2_X1 U616 ( .A1(G64), .A2(n643), .ZN(n554) );
  AND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U618 ( .A1(n557), .A2(n556), .ZN(G301) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n558), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U621 ( .A(G223), .ZN(n823) );
  NAND2_X1 U622 ( .A1(n823), .A2(G567), .ZN(n559) );
  XOR2_X1 U623 ( .A(KEYINPUT11), .B(n559), .Z(G234) );
  NAND2_X1 U624 ( .A1(G81), .A2(n630), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT69), .B(n560), .Z(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(KEYINPUT12), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G68), .A2(n628), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT13), .B(n564), .Z(n569) );
  XOR2_X1 U630 ( .A(KEYINPUT68), .B(KEYINPUT14), .Z(n566) );
  NAND2_X1 U631 ( .A1(G56), .A2(n643), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT67), .B(n567), .Z(n568) );
  NOR2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(KEYINPUT70), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G43), .A2(n644), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n855) );
  INV_X1 U638 ( .A(G860), .ZN(n604) );
  OR2_X1 U639 ( .A1(n855), .A2(n604), .ZN(G153) );
  NAND2_X1 U640 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U641 ( .A1(G66), .A2(n643), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G92), .A2(n630), .ZN(n574) );
  NAND2_X1 U643 ( .A1(G79), .A2(n628), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U645 ( .A1(G54), .A2(n644), .ZN(n575) );
  XNOR2_X1 U646 ( .A(KEYINPUT71), .B(n575), .ZN(n576) );
  NOR2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U649 ( .A(n580), .B(KEYINPUT15), .ZN(n958) );
  OR2_X1 U650 ( .A1(n958), .A2(G868), .ZN(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U652 ( .A1(G51), .A2(n644), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n643), .A2(G63), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U655 ( .A(KEYINPUT6), .B(n585), .ZN(n591) );
  NAND2_X1 U656 ( .A1(n630), .A2(G89), .ZN(n586) );
  XNOR2_X1 U657 ( .A(n586), .B(KEYINPUT4), .ZN(n588) );
  NAND2_X1 U658 ( .A1(G76), .A2(n628), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U660 ( .A(n589), .B(KEYINPUT5), .Z(n590) );
  NOR2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U662 ( .A(KEYINPUT7), .B(n592), .Z(n593) );
  XNOR2_X1 U663 ( .A(KEYINPUT72), .B(n593), .ZN(G168) );
  XOR2_X1 U664 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U665 ( .A1(G65), .A2(n643), .ZN(n595) );
  NAND2_X1 U666 ( .A1(G53), .A2(n644), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U668 ( .A1(G91), .A2(n630), .ZN(n597) );
  NAND2_X1 U669 ( .A1(G78), .A2(n628), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U671 ( .A1(n599), .A2(n598), .ZN(n1017) );
  INV_X1 U672 ( .A(G868), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n1017), .A2(n601), .ZN(n600) );
  XNOR2_X1 U674 ( .A(n600), .B(KEYINPUT73), .ZN(n603) );
  NOR2_X1 U675 ( .A1(G286), .A2(n601), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n603), .A2(n602), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n604), .A2(G559), .ZN(n605) );
  NAND2_X1 U678 ( .A1(n605), .A2(n958), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n855), .ZN(n607) );
  XNOR2_X1 U681 ( .A(KEYINPUT74), .B(n607), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G868), .A2(n958), .ZN(n608) );
  NOR2_X1 U683 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U684 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U685 ( .A1(n958), .A2(G559), .ZN(n655) );
  XNOR2_X1 U686 ( .A(n855), .B(n655), .ZN(n611) );
  NOR2_X1 U687 ( .A1(n611), .A2(G860), .ZN(n618) );
  NAND2_X1 U688 ( .A1(G93), .A2(n630), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G80), .A2(n628), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U691 ( .A1(G67), .A2(n643), .ZN(n615) );
  NAND2_X1 U692 ( .A1(G55), .A2(n644), .ZN(n614) );
  NAND2_X1 U693 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n657) );
  XNOR2_X1 U695 ( .A(n618), .B(n657), .ZN(G145) );
  NAND2_X1 U696 ( .A1(G88), .A2(n630), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n619), .B(KEYINPUT82), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G75), .A2(n628), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G62), .A2(n643), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G50), .A2(n644), .ZN(n622) );
  XNOR2_X1 U702 ( .A(KEYINPUT81), .B(n622), .ZN(n623) );
  NOR2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U704 ( .A1(n626), .A2(n625), .ZN(G303) );
  INV_X1 U705 ( .A(G303), .ZN(G166) );
  NAND2_X1 U706 ( .A1(G48), .A2(n644), .ZN(n627) );
  XNOR2_X1 U707 ( .A(KEYINPUT80), .B(n627), .ZN(n638) );
  NAND2_X1 U708 ( .A1(n628), .A2(G73), .ZN(n629) );
  XNOR2_X1 U709 ( .A(KEYINPUT2), .B(n629), .ZN(n635) );
  NAND2_X1 U710 ( .A1(G86), .A2(n630), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G61), .A2(n643), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U713 ( .A(KEYINPUT78), .B(n633), .Z(n634) );
  NAND2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U715 ( .A(KEYINPUT79), .B(n636), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U717 ( .A1(G74), .A2(G651), .ZN(n641) );
  NAND2_X1 U718 ( .A1(G87), .A2(n639), .ZN(n640) );
  NAND2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U720 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n644), .A2(G49), .ZN(n645) );
  XOR2_X1 U722 ( .A(KEYINPUT77), .B(n645), .Z(n646) );
  NAND2_X1 U723 ( .A1(n647), .A2(n646), .ZN(G288) );
  XNOR2_X1 U724 ( .A(G166), .B(G305), .ZN(n648) );
  XNOR2_X1 U725 ( .A(n648), .B(G288), .ZN(n651) );
  XOR2_X1 U726 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n649) );
  XNOR2_X1 U727 ( .A(G290), .B(n649), .ZN(n650) );
  XOR2_X1 U728 ( .A(n651), .B(n650), .Z(n653) );
  XNOR2_X1 U729 ( .A(n1017), .B(n657), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n654), .B(n855), .ZN(n957) );
  XOR2_X1 U732 ( .A(n957), .B(n655), .Z(n656) );
  NAND2_X1 U733 ( .A1(G868), .A2(n656), .ZN(n659) );
  OR2_X1 U734 ( .A1(n657), .A2(G868), .ZN(n658) );
  NAND2_X1 U735 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U736 ( .A1(G2084), .A2(G2078), .ZN(n660) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n661), .ZN(n662) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n662), .ZN(n663) );
  NAND2_X1 U740 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U741 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U742 ( .A(KEYINPUT66), .B(G132), .Z(G219) );
  NAND2_X1 U743 ( .A1(G120), .A2(G69), .ZN(n664) );
  XNOR2_X1 U744 ( .A(KEYINPUT84), .B(n664), .ZN(n665) );
  NOR2_X1 U745 ( .A1(G238), .A2(n665), .ZN(n666) );
  NAND2_X1 U746 ( .A1(G57), .A2(n666), .ZN(n955) );
  NAND2_X1 U747 ( .A1(n955), .A2(G567), .ZN(n671) );
  NOR2_X1 U748 ( .A1(G219), .A2(G220), .ZN(n667) );
  XOR2_X1 U749 ( .A(KEYINPUT22), .B(n667), .Z(n668) );
  NOR2_X1 U750 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U751 ( .A1(G96), .A2(n669), .ZN(n956) );
  NAND2_X1 U752 ( .A1(n956), .A2(G2106), .ZN(n670) );
  NAND2_X1 U753 ( .A1(n671), .A2(n670), .ZN(n1016) );
  NAND2_X1 U754 ( .A1(G661), .A2(G483), .ZN(n672) );
  XOR2_X1 U755 ( .A(KEYINPUT85), .B(n672), .Z(n673) );
  NOR2_X1 U756 ( .A1(n1016), .A2(n673), .ZN(n826) );
  NAND2_X1 U757 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U758 ( .A1(G114), .A2(n993), .ZN(n675) );
  NAND2_X1 U759 ( .A1(G126), .A2(n994), .ZN(n674) );
  NAND2_X1 U760 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U761 ( .A(KEYINPUT86), .B(n676), .ZN(n680) );
  NAND2_X1 U762 ( .A1(G102), .A2(n997), .ZN(n678) );
  NAND2_X1 U763 ( .A1(G138), .A2(n998), .ZN(n677) );
  NAND2_X1 U764 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U765 ( .A1(n680), .A2(n679), .ZN(G164) );
  NOR2_X1 U766 ( .A1(G164), .A2(G1384), .ZN(n700) );
  NAND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n699) );
  NOR2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n818) );
  NAND2_X1 U769 ( .A1(G117), .A2(n993), .ZN(n682) );
  NAND2_X1 U770 ( .A1(G129), .A2(n994), .ZN(n681) );
  NAND2_X1 U771 ( .A1(n682), .A2(n681), .ZN(n685) );
  NAND2_X1 U772 ( .A1(n997), .A2(G105), .ZN(n683) );
  XOR2_X1 U773 ( .A(KEYINPUT38), .B(n683), .Z(n684) );
  NOR2_X1 U774 ( .A1(n685), .A2(n684), .ZN(n687) );
  NAND2_X1 U775 ( .A1(n998), .A2(G141), .ZN(n686) );
  NAND2_X1 U776 ( .A1(n687), .A2(n686), .ZN(n1004) );
  NAND2_X1 U777 ( .A1(G1996), .A2(n1004), .ZN(n688) );
  XOR2_X1 U778 ( .A(KEYINPUT89), .B(n688), .Z(n696) );
  NAND2_X1 U779 ( .A1(G107), .A2(n993), .ZN(n690) );
  NAND2_X1 U780 ( .A1(G119), .A2(n994), .ZN(n689) );
  NAND2_X1 U781 ( .A1(n690), .A2(n689), .ZN(n694) );
  NAND2_X1 U782 ( .A1(G95), .A2(n997), .ZN(n692) );
  NAND2_X1 U783 ( .A1(G131), .A2(n998), .ZN(n691) );
  NAND2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n693) );
  OR2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n990) );
  NAND2_X1 U786 ( .A1(G1991), .A2(n990), .ZN(n695) );
  NAND2_X1 U787 ( .A1(n696), .A2(n695), .ZN(n916) );
  NAND2_X1 U788 ( .A1(n818), .A2(n916), .ZN(n807) );
  XNOR2_X1 U789 ( .A(G1986), .B(G290), .ZN(n843) );
  NAND2_X1 U790 ( .A1(n843), .A2(n818), .ZN(n697) );
  XOR2_X1 U791 ( .A(KEYINPUT87), .B(n697), .Z(n698) );
  NAND2_X1 U792 ( .A1(n807), .A2(n698), .ZN(n795) );
  INV_X1 U793 ( .A(n699), .ZN(n701) );
  NAND2_X1 U794 ( .A1(G8), .A2(n761), .ZN(n788) );
  NOR2_X1 U795 ( .A1(G1981), .A2(G305), .ZN(n702) );
  XOR2_X1 U796 ( .A(n702), .B(KEYINPUT24), .Z(n703) );
  NOR2_X1 U797 ( .A1(n788), .A2(n703), .ZN(n793) );
  INV_X1 U798 ( .A(n712), .ZN(n734) );
  XNOR2_X1 U799 ( .A(KEYINPUT26), .B(KEYINPUT93), .ZN(n704) );
  XNOR2_X1 U800 ( .A(n705), .B(n704), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n761), .A2(G1341), .ZN(n706) );
  NAND2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U803 ( .A1(n958), .A2(n710), .ZN(n709) );
  XNOR2_X1 U804 ( .A(n709), .B(KEYINPUT95), .ZN(n719) );
  NAND2_X1 U805 ( .A1(n958), .A2(n710), .ZN(n717) );
  INV_X1 U806 ( .A(KEYINPUT90), .ZN(n711) );
  XOR2_X1 U807 ( .A(n712), .B(n711), .Z(n733) );
  INV_X1 U808 ( .A(n733), .ZN(n721) );
  NAND2_X1 U809 ( .A1(G2067), .A2(n721), .ZN(n713) );
  XNOR2_X1 U810 ( .A(n713), .B(KEYINPUT94), .ZN(n715) );
  NAND2_X1 U811 ( .A1(G1348), .A2(n761), .ZN(n714) );
  NAND2_X1 U812 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U813 ( .A1(n717), .A2(n716), .ZN(n718) );
  NAND2_X1 U814 ( .A1(n719), .A2(n718), .ZN(n725) );
  NAND2_X1 U815 ( .A1(n721), .A2(G2072), .ZN(n720) );
  XNOR2_X1 U816 ( .A(n720), .B(KEYINPUT27), .ZN(n723) );
  INV_X1 U817 ( .A(G1956), .ZN(n872) );
  NOR2_X1 U818 ( .A1(n721), .A2(n872), .ZN(n722) );
  NOR2_X1 U819 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n726), .A2(n1017), .ZN(n724) );
  NAND2_X1 U821 ( .A1(n725), .A2(n724), .ZN(n730) );
  NOR2_X1 U822 ( .A1(n726), .A2(n1017), .ZN(n728) );
  XNOR2_X1 U823 ( .A(n728), .B(n727), .ZN(n729) );
  NAND2_X1 U824 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U825 ( .A(n731), .B(KEYINPUT29), .ZN(n739) );
  XNOR2_X1 U826 ( .A(G2078), .B(KEYINPUT25), .ZN(n732) );
  XNOR2_X1 U827 ( .A(n732), .B(KEYINPUT91), .ZN(n939) );
  NOR2_X1 U828 ( .A1(n939), .A2(n733), .ZN(n736) );
  NOR2_X1 U829 ( .A1(n734), .A2(G1961), .ZN(n735) );
  NOR2_X1 U830 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U831 ( .A(KEYINPUT92), .B(n737), .ZN(n742) );
  NOR2_X1 U832 ( .A1(G301), .A2(n742), .ZN(n738) );
  XNOR2_X1 U833 ( .A(n741), .B(n740), .ZN(n751) );
  NAND2_X1 U834 ( .A1(G301), .A2(n742), .ZN(n743) );
  XNOR2_X1 U835 ( .A(n743), .B(KEYINPUT97), .ZN(n748) );
  NOR2_X1 U836 ( .A1(G2084), .A2(n761), .ZN(n755) );
  NOR2_X1 U837 ( .A1(G1966), .A2(n788), .ZN(n752) );
  NOR2_X1 U838 ( .A1(n755), .A2(n752), .ZN(n744) );
  NAND2_X1 U839 ( .A1(G8), .A2(n744), .ZN(n745) );
  XNOR2_X1 U840 ( .A(KEYINPUT30), .B(n745), .ZN(n746) );
  NOR2_X1 U841 ( .A1(G168), .A2(n746), .ZN(n747) );
  NOR2_X1 U842 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U843 ( .A(KEYINPUT31), .B(n749), .Z(n750) );
  NAND2_X1 U844 ( .A1(n751), .A2(n750), .ZN(n760) );
  INV_X1 U845 ( .A(n760), .ZN(n753) );
  XNOR2_X1 U846 ( .A(n754), .B(KEYINPUT98), .ZN(n757) );
  NAND2_X1 U847 ( .A1(n755), .A2(G8), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n757), .A2(n756), .ZN(n784) );
  NAND2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n837) );
  INV_X1 U850 ( .A(n788), .ZN(n758) );
  NAND2_X1 U851 ( .A1(n837), .A2(n758), .ZN(n775) );
  INV_X1 U852 ( .A(n775), .ZN(n759) );
  AND2_X1 U853 ( .A1(n784), .A2(n759), .ZN(n772) );
  NAND2_X1 U854 ( .A1(n760), .A2(G286), .ZN(n766) );
  NOR2_X1 U855 ( .A1(G1971), .A2(n788), .ZN(n763) );
  NOR2_X1 U856 ( .A1(G2090), .A2(n761), .ZN(n762) );
  NOR2_X1 U857 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n764), .A2(G303), .ZN(n765) );
  NAND2_X1 U859 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U860 ( .A1(n767), .A2(G8), .ZN(n768) );
  XNOR2_X1 U861 ( .A(n768), .B(KEYINPUT32), .ZN(n783) );
  NOR2_X1 U862 ( .A1(G1976), .A2(G288), .ZN(n774) );
  NAND2_X1 U863 ( .A1(n774), .A2(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U864 ( .A1(n769), .A2(n788), .ZN(n779) );
  INV_X1 U865 ( .A(n779), .ZN(n770) );
  AND2_X1 U866 ( .A1(n783), .A2(n770), .ZN(n771) );
  NAND2_X1 U867 ( .A1(n772), .A2(n771), .ZN(n781) );
  INV_X1 U868 ( .A(KEYINPUT33), .ZN(n777) );
  NOR2_X1 U869 ( .A1(G1971), .A2(G303), .ZN(n773) );
  NOR2_X1 U870 ( .A1(n774), .A2(n773), .ZN(n838) );
  OR2_X1 U871 ( .A1(n775), .A2(n838), .ZN(n776) );
  AND2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n778) );
  OR2_X1 U873 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U875 ( .A(G1981), .B(G305), .Z(n847) );
  NAND2_X1 U876 ( .A1(n782), .A2(n847), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n784), .A2(n783), .ZN(n787) );
  NOR2_X1 U878 ( .A1(G2090), .A2(G303), .ZN(n785) );
  NAND2_X1 U879 ( .A1(G8), .A2(n785), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U883 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n806) );
  NAND2_X1 U885 ( .A1(G104), .A2(n997), .ZN(n797) );
  NAND2_X1 U886 ( .A1(G140), .A2(n998), .ZN(n796) );
  NAND2_X1 U887 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U888 ( .A(KEYINPUT34), .B(n798), .ZN(n804) );
  NAND2_X1 U889 ( .A1(G116), .A2(n993), .ZN(n800) );
  NAND2_X1 U890 ( .A1(G128), .A2(n994), .ZN(n799) );
  NAND2_X1 U891 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U892 ( .A(KEYINPUT88), .B(n801), .Z(n802) );
  XNOR2_X1 U893 ( .A(KEYINPUT35), .B(n802), .ZN(n803) );
  NOR2_X1 U894 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U895 ( .A(KEYINPUT36), .B(n805), .ZN(n986) );
  XNOR2_X1 U896 ( .A(G2067), .B(KEYINPUT37), .ZN(n816) );
  NOR2_X1 U897 ( .A1(n986), .A2(n816), .ZN(n906) );
  NAND2_X1 U898 ( .A1(n906), .A2(n818), .ZN(n815) );
  NAND2_X1 U899 ( .A1(n806), .A2(n815), .ZN(n821) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n1004), .ZN(n909) );
  INV_X1 U901 ( .A(n807), .ZN(n810) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n808) );
  NOR2_X1 U903 ( .A1(G1991), .A2(n990), .ZN(n903) );
  NOR2_X1 U904 ( .A1(n808), .A2(n903), .ZN(n809) );
  NOR2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U906 ( .A1(n909), .A2(n811), .ZN(n812) );
  XOR2_X1 U907 ( .A(n812), .B(KEYINPUT99), .Z(n813) );
  XNOR2_X1 U908 ( .A(KEYINPUT39), .B(n813), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n986), .A2(n816), .ZN(n913) );
  NAND2_X1 U911 ( .A1(n817), .A2(n913), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U914 ( .A(n822), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U915 ( .A(G301), .ZN(G171) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U918 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(G188) );
  XOR2_X1 U921 ( .A(G96), .B(KEYINPUT100), .Z(G221) );
  XNOR2_X1 U922 ( .A(G69), .B(KEYINPUT101), .ZN(G235) );
  NAND2_X1 U924 ( .A1(G136), .A2(n998), .ZN(n833) );
  NAND2_X1 U925 ( .A1(G100), .A2(n997), .ZN(n828) );
  NAND2_X1 U926 ( .A1(G112), .A2(n993), .ZN(n827) );
  NAND2_X1 U927 ( .A1(n828), .A2(n827), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n994), .A2(G124), .ZN(n829) );
  XOR2_X1 U929 ( .A(KEYINPUT44), .B(n829), .Z(n830) );
  NOR2_X1 U930 ( .A1(n831), .A2(n830), .ZN(n832) );
  NAND2_X1 U931 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n834), .B(KEYINPUT105), .ZN(G162) );
  XNOR2_X1 U933 ( .A(KEYINPUT56), .B(G16), .ZN(n861) );
  XNOR2_X1 U934 ( .A(n872), .B(n1017), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n835), .B(KEYINPUT121), .ZN(n845) );
  INV_X1 U936 ( .A(G1971), .ZN(n836) );
  NOR2_X1 U937 ( .A1(G166), .A2(n836), .ZN(n840) );
  NAND2_X1 U938 ( .A1(n838), .A2(n837), .ZN(n839) );
  NOR2_X1 U939 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U940 ( .A(KEYINPUT122), .B(n841), .Z(n842) );
  NOR2_X1 U941 ( .A1(n843), .A2(n842), .ZN(n844) );
  NAND2_X1 U942 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U943 ( .A(KEYINPUT123), .B(n846), .ZN(n859) );
  XNOR2_X1 U944 ( .A(G1966), .B(G168), .ZN(n848) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U946 ( .A(KEYINPUT57), .B(n849), .ZN(n854) );
  XOR2_X1 U947 ( .A(n958), .B(G1348), .Z(n850) );
  XNOR2_X1 U948 ( .A(KEYINPUT120), .B(n850), .ZN(n852) );
  XNOR2_X1 U949 ( .A(G1961), .B(G301), .ZN(n851) );
  NOR2_X1 U950 ( .A1(n852), .A2(n851), .ZN(n853) );
  NAND2_X1 U951 ( .A1(n854), .A2(n853), .ZN(n857) );
  XNOR2_X1 U952 ( .A(G1341), .B(n855), .ZN(n856) );
  NOR2_X1 U953 ( .A1(n857), .A2(n856), .ZN(n858) );
  NAND2_X1 U954 ( .A1(n859), .A2(n858), .ZN(n860) );
  NAND2_X1 U955 ( .A1(n861), .A2(n860), .ZN(n929) );
  XNOR2_X1 U956 ( .A(G1986), .B(G24), .ZN(n866) );
  XNOR2_X1 U957 ( .A(G1971), .B(G22), .ZN(n863) );
  XNOR2_X1 U958 ( .A(G1976), .B(G23), .ZN(n862) );
  NOR2_X1 U959 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U960 ( .A(KEYINPUT125), .B(n864), .ZN(n865) );
  NOR2_X1 U961 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U962 ( .A(KEYINPUT58), .B(n867), .ZN(n871) );
  XNOR2_X1 U963 ( .A(G1966), .B(G21), .ZN(n869) );
  XNOR2_X1 U964 ( .A(G5), .B(G1961), .ZN(n868) );
  NOR2_X1 U965 ( .A1(n869), .A2(n868), .ZN(n870) );
  NAND2_X1 U966 ( .A1(n871), .A2(n870), .ZN(n883) );
  XNOR2_X1 U967 ( .A(G20), .B(n872), .ZN(n876) );
  XNOR2_X1 U968 ( .A(G1341), .B(G19), .ZN(n874) );
  XNOR2_X1 U969 ( .A(G1981), .B(G6), .ZN(n873) );
  NOR2_X1 U970 ( .A1(n874), .A2(n873), .ZN(n875) );
  NAND2_X1 U971 ( .A1(n876), .A2(n875), .ZN(n880) );
  XOR2_X1 U972 ( .A(KEYINPUT124), .B(G4), .Z(n878) );
  XNOR2_X1 U973 ( .A(G1348), .B(KEYINPUT59), .ZN(n877) );
  XNOR2_X1 U974 ( .A(n878), .B(n877), .ZN(n879) );
  NOR2_X1 U975 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U976 ( .A(KEYINPUT60), .B(n881), .Z(n882) );
  NOR2_X1 U977 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U978 ( .A(KEYINPUT61), .B(n884), .Z(n885) );
  NOR2_X1 U979 ( .A1(G16), .A2(n885), .ZN(n886) );
  XOR2_X1 U980 ( .A(KEYINPUT126), .B(n886), .Z(n887) );
  NAND2_X1 U981 ( .A1(G11), .A2(n887), .ZN(n927) );
  INV_X1 U982 ( .A(G29), .ZN(n924) );
  XOR2_X1 U983 ( .A(G164), .B(G2078), .Z(n899) );
  NAND2_X1 U984 ( .A1(G103), .A2(n997), .ZN(n896) );
  XNOR2_X1 U985 ( .A(KEYINPUT47), .B(KEYINPUT107), .ZN(n891) );
  NAND2_X1 U986 ( .A1(G115), .A2(n993), .ZN(n889) );
  NAND2_X1 U987 ( .A1(G127), .A2(n994), .ZN(n888) );
  NAND2_X1 U988 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n891), .B(n890), .ZN(n894) );
  NAND2_X1 U990 ( .A1(n998), .A2(G139), .ZN(n892) );
  XOR2_X1 U991 ( .A(KEYINPUT106), .B(n892), .Z(n893) );
  NOR2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n895) );
  NAND2_X1 U993 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n897), .B(KEYINPUT108), .ZN(n989) );
  XNOR2_X1 U995 ( .A(G2072), .B(n989), .ZN(n898) );
  NOR2_X1 U996 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U997 ( .A(KEYINPUT50), .B(n900), .Z(n919) );
  XNOR2_X1 U998 ( .A(G160), .B(G2084), .ZN(n901) );
  NAND2_X1 U999 ( .A1(n901), .A2(n982), .ZN(n902) );
  NOR2_X1 U1000 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n904), .B(KEYINPUT111), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(n906), .A2(n905), .ZN(n907) );
  XOR2_X1 U1003 ( .A(KEYINPUT112), .B(n907), .Z(n912) );
  XOR2_X1 U1004 ( .A(G2090), .B(G162), .Z(n908) );
  NOR2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(KEYINPUT51), .B(n910), .ZN(n911) );
  NOR2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(n914) );
  NAND2_X1 U1008 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1010 ( .A(KEYINPUT113), .B(n917), .ZN(n918) );
  NOR2_X1 U1011 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1012 ( .A(n920), .B(KEYINPUT114), .Z(n921) );
  XNOR2_X1 U1013 ( .A(KEYINPUT52), .B(n921), .ZN(n922) );
  NOR2_X1 U1014 ( .A1(KEYINPUT55), .A2(n922), .ZN(n923) );
  NOR2_X1 U1015 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1016 ( .A(KEYINPUT115), .B(n925), .Z(n926) );
  NOR2_X1 U1017 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1018 ( .A1(n929), .A2(n928), .ZN(n953) );
  XNOR2_X1 U1019 ( .A(G33), .B(G2072), .ZN(n930) );
  XNOR2_X1 U1020 ( .A(n930), .B(KEYINPUT117), .ZN(n938) );
  XNOR2_X1 U1021 ( .A(G1996), .B(G32), .ZN(n932) );
  XNOR2_X1 U1022 ( .A(G1991), .B(G25), .ZN(n931) );
  NOR2_X1 U1023 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1024 ( .A1(G28), .A2(n933), .ZN(n936) );
  XNOR2_X1 U1025 ( .A(KEYINPUT116), .B(G2067), .ZN(n934) );
  XNOR2_X1 U1026 ( .A(G26), .B(n934), .ZN(n935) );
  NOR2_X1 U1027 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1028 ( .A1(n938), .A2(n937), .ZN(n941) );
  XNOR2_X1 U1029 ( .A(G27), .B(n939), .ZN(n940) );
  NOR2_X1 U1030 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1031 ( .A(KEYINPUT53), .B(n942), .Z(n945) );
  XOR2_X1 U1032 ( .A(G34), .B(KEYINPUT54), .Z(n943) );
  XNOR2_X1 U1033 ( .A(G2084), .B(n943), .ZN(n944) );
  NAND2_X1 U1034 ( .A1(n945), .A2(n944), .ZN(n947) );
  XNOR2_X1 U1035 ( .A(G35), .B(G2090), .ZN(n946) );
  NOR2_X1 U1036 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1037 ( .A(KEYINPUT55), .B(n948), .Z(n950) );
  XNOR2_X1 U1038 ( .A(KEYINPUT118), .B(G29), .ZN(n949) );
  NOR2_X1 U1039 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1040 ( .A(KEYINPUT119), .B(n951), .Z(n952) );
  NOR2_X1 U1041 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1042 ( .A(KEYINPUT62), .B(n954), .ZN(G311) );
  XNOR2_X1 U1043 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1044 ( .A(G120), .ZN(G236) );
  NOR2_X1 U1045 ( .A1(n956), .A2(n955), .ZN(G325) );
  INV_X1 U1046 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1047 ( .A(G286), .B(n957), .ZN(n960) );
  XNOR2_X1 U1048 ( .A(G171), .B(n958), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(n960), .B(n959), .ZN(n961) );
  NOR2_X1 U1050 ( .A1(G37), .A2(n961), .ZN(G397) );
  XNOR2_X1 U1051 ( .A(G1976), .B(G2474), .ZN(n971) );
  XOR2_X1 U1052 ( .A(G1986), .B(G1971), .Z(n963) );
  XNOR2_X1 U1053 ( .A(G1966), .B(G1961), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(n963), .B(n962), .ZN(n967) );
  XOR2_X1 U1055 ( .A(KEYINPUT104), .B(KEYINPUT41), .Z(n965) );
  XNOR2_X1 U1056 ( .A(G1996), .B(G1991), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n965), .B(n964), .ZN(n966) );
  XOR2_X1 U1058 ( .A(n967), .B(n966), .Z(n969) );
  XNOR2_X1 U1059 ( .A(G1956), .B(G1981), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n969), .B(n968), .ZN(n970) );
  XNOR2_X1 U1061 ( .A(n971), .B(n970), .ZN(G229) );
  XOR2_X1 U1062 ( .A(KEYINPUT103), .B(G2678), .Z(n973) );
  XNOR2_X1 U1063 ( .A(G2072), .B(G2090), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(n973), .B(n972), .ZN(n977) );
  XOR2_X1 U1065 ( .A(KEYINPUT43), .B(KEYINPUT102), .Z(n975) );
  XNOR2_X1 U1066 ( .A(G2067), .B(KEYINPUT42), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n975), .B(n974), .ZN(n976) );
  XOR2_X1 U1068 ( .A(n977), .B(n976), .Z(n979) );
  XNOR2_X1 U1069 ( .A(G2096), .B(G2100), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(n979), .B(n978), .ZN(n981) );
  XOR2_X1 U1071 ( .A(G2084), .B(G2078), .Z(n980) );
  XNOR2_X1 U1072 ( .A(n981), .B(n980), .ZN(G227) );
  XNOR2_X1 U1073 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(n982), .B(KEYINPUT109), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(n984), .B(n983), .ZN(n988) );
  XOR2_X1 U1076 ( .A(G160), .B(G162), .Z(n985) );
  XNOR2_X1 U1077 ( .A(n986), .B(n985), .ZN(n987) );
  XNOR2_X1 U1078 ( .A(n988), .B(n987), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(n990), .B(n989), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(n992), .B(n991), .ZN(n1008) );
  NAND2_X1 U1081 ( .A1(G118), .A2(n993), .ZN(n996) );
  NAND2_X1 U1082 ( .A1(G130), .A2(n994), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n1003) );
  NAND2_X1 U1084 ( .A1(G106), .A2(n997), .ZN(n1000) );
  NAND2_X1 U1085 ( .A1(G142), .A2(n998), .ZN(n999) );
  NAND2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1087 ( .A(n1001), .B(KEYINPUT45), .Z(n1002) );
  NOR2_X1 U1088 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1089 ( .A(n1005), .B(n1004), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(G164), .B(n1006), .ZN(n1007) );
  XNOR2_X1 U1091 ( .A(n1008), .B(n1007), .ZN(n1009) );
  NOR2_X1 U1092 ( .A1(G37), .A2(n1009), .ZN(G395) );
  NOR2_X1 U1093 ( .A1(G229), .A2(G227), .ZN(n1010) );
  XNOR2_X1 U1094 ( .A(KEYINPUT49), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1095 ( .A1(G397), .A2(n1011), .ZN(n1015) );
  NOR2_X1 U1096 ( .A1(n1016), .A2(G401), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(KEYINPUT110), .B(n1012), .Z(n1013) );
  NOR2_X1 U1098 ( .A1(G395), .A2(n1013), .ZN(n1014) );
  NAND2_X1 U1099 ( .A1(n1015), .A2(n1014), .ZN(G225) );
  INV_X1 U1100 ( .A(G225), .ZN(G308) );
  INV_X1 U1101 ( .A(n1016), .ZN(G319) );
  INV_X1 U1102 ( .A(G57), .ZN(G237) );
  INV_X1 U1103 ( .A(n1017), .ZN(G299) );
endmodule

