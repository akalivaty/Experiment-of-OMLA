//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT5), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT82), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G155gat), .ZN(new_n206));
  INV_X1    g005(.A(G162gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n205), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT83), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G141gat), .ZN(new_n213));
  INV_X1    g012(.A(G141gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G148gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n217));
  AOI22_X1  g016(.A1(new_n210), .A2(new_n211), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n205), .A2(new_n208), .A3(KEYINPUT83), .A4(new_n209), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT84), .B(G141gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n213), .B1(new_n220), .B2(new_n212), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n203), .B1(new_n208), .B2(KEYINPUT2), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n218), .A2(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G134gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G127gat), .ZN(new_n225));
  INV_X1    g024(.A(G127gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G134gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(KEYINPUT1), .ZN(new_n230));
  INV_X1    g029(.A(G120gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G113gat), .ZN(new_n232));
  INV_X1    g031(.A(G113gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G120gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G127gat), .B(G134gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n230), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n210), .A2(new_n211), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n216), .A2(new_n217), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n219), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n221), .A2(new_n222), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n239), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n241), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n202), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  AND3_X1   g050(.A1(new_n230), .A2(new_n238), .A3(KEYINPUT70), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT70), .B1(new_n230), .B2(new_n238), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT4), .B1(new_n254), .B2(new_n246), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n223), .A2(new_n240), .A3(new_n256), .ZN(new_n257));
  AND3_X1   g056(.A1(new_n255), .A2(KEYINPUT85), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n240), .B1(new_n246), .B2(KEYINPUT3), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT3), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n223), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT85), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n263), .B(KEYINPUT4), .C1(new_n254), .C2(new_n246), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n264), .A3(new_n249), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n251), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n256), .B1(new_n254), .B2(new_n246), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n223), .A2(new_n240), .A3(KEYINPUT4), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n267), .A2(new_n202), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n250), .B1(new_n259), .B2(new_n261), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G1gat), .B(G29gat), .Z(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G57gat), .B(G85gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n255), .A2(KEYINPUT85), .A3(new_n257), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(new_n264), .A3(new_n270), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n283), .A2(new_n251), .B1(new_n269), .B2(new_n270), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(new_n277), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n266), .A2(new_n277), .A3(new_n271), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n280), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT87), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n285), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT6), .B1(new_n284), .B2(new_n277), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT87), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n281), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT81), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n294), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT26), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(KEYINPUT28), .A3(new_n301), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n299), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G226gat), .ZN(new_n308));
  INV_X1    g107(.A(G233gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312));
  NOR4_X1   g111(.A1(new_n312), .A2(KEYINPUT66), .A3(G169gat), .A4(G176gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT66), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n294), .B2(KEYINPUT23), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT67), .B1(new_n294), .B2(KEYINPUT23), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT67), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n318), .B(new_n312), .C1(G169gat), .C2(G176gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n296), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT24), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT65), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n322), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT64), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT64), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n330), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT65), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n327), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT25), .B1(new_n321), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT25), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(new_n294), .B2(KEYINPUT23), .ZN(new_n338));
  AND4_X1   g137(.A1(new_n317), .A2(new_n338), .A3(new_n296), .A4(new_n319), .ZN(new_n339));
  OR2_X1    g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT68), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n340), .B(new_n328), .C1(new_n333), .C2(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n325), .A2(KEYINPUT68), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT69), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n340), .A2(new_n328), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n325), .A2(KEYINPUT68), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT69), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n333), .A2(new_n341), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n339), .A2(new_n344), .A3(new_n349), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n307), .B(new_n311), .C1(new_n336), .C2(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n317), .A2(new_n338), .A3(new_n296), .A4(new_n319), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n342), .A2(new_n343), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(new_n347), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n344), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n317), .A2(new_n296), .A3(new_n319), .ZN(new_n356));
  INV_X1    g155(.A(new_n315), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n294), .A2(new_n314), .A3(KEYINPUT23), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n335), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n337), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n306), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n310), .A2(KEYINPUT29), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n351), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT77), .ZN(new_n365));
  XNOR2_X1  g164(.A(G211gat), .B(G218gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(G211gat), .A2(G218gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT22), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G197gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT75), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT75), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G197gat), .ZN(new_n373));
  AND3_X1   g172(.A1(new_n371), .A2(new_n373), .A3(G204gat), .ZN(new_n374));
  AOI21_X1  g173(.A(G204gat), .B1(new_n371), .B2(new_n373), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n366), .B(new_n369), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(G204gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n372), .A2(G197gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n370), .A2(KEYINPUT75), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n371), .A2(new_n373), .A3(G204gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n366), .B1(new_n384), .B2(new_n369), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n369), .B1(new_n374), .B2(new_n375), .ZN(new_n387));
  INV_X1    g186(.A(new_n366), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(KEYINPUT76), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n365), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(new_n388), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n392), .A2(new_n377), .A3(new_n376), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(KEYINPUT77), .A3(new_n389), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n364), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n389), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n351), .B(new_n397), .C1(new_n362), .C2(new_n363), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(G8gat), .B(G36gat), .Z(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(KEYINPUT79), .ZN(new_n401));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n293), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  AOI211_X1 g205(.A(KEYINPUT81), .B(new_n403), .C1(new_n396), .C2(new_n398), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n398), .ZN(new_n411));
  INV_X1    g210(.A(new_n363), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n344), .A2(new_n354), .B1(new_n360), .B2(new_n337), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n412), .B1(new_n413), .B2(new_n306), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n414), .A2(new_n351), .B1(new_n391), .B2(new_n394), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT78), .B1(new_n411), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n403), .B(KEYINPUT80), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT78), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n396), .A2(new_n418), .A3(new_n398), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n416), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n399), .A2(KEYINPUT30), .A3(new_n404), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n410), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n292), .A2(new_n422), .ZN(new_n423));
  OAI22_X1  g222(.A1(new_n413), .A2(new_n306), .B1(new_n252), .B2(new_n253), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n254), .B(new_n307), .C1(new_n336), .C2(new_n350), .ZN(new_n425));
  INV_X1    g224(.A(G227gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(new_n309), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT32), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT33), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  XOR2_X1   g230(.A(G15gat), .B(G43gat), .Z(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT71), .ZN(new_n433));
  XNOR2_X1  g232(.A(G71gat), .B(G99gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(new_n431), .A3(new_n436), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n435), .A2(KEYINPUT72), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n435), .A2(KEYINPUT72), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(KEYINPUT33), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(KEYINPUT32), .A3(new_n428), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n427), .B1(new_n424), .B2(new_n425), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT73), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT34), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n446), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n443), .A2(new_n447), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n437), .A2(new_n450), .A3(new_n446), .A4(new_n441), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT29), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n393), .A2(new_n453), .A3(new_n389), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n260), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n246), .ZN(new_n456));
  INV_X1    g255(.A(G228gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(new_n309), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n261), .A2(new_n453), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n391), .A2(new_n394), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n392), .A2(new_n462), .A3(new_n376), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n384), .A2(KEYINPUT88), .A3(new_n366), .A4(new_n369), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n463), .A2(new_n453), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n223), .B1(new_n465), .B2(new_n260), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n453), .A2(new_n261), .B1(new_n393), .B2(new_n389), .ZN(new_n467));
  OAI22_X1  g266(.A1(new_n466), .A2(new_n467), .B1(new_n457), .B2(new_n309), .ZN(new_n468));
  INV_X1    g267(.A(G22gat), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n461), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n469), .B1(new_n461), .B2(new_n468), .ZN(new_n471));
  OAI21_X1  g270(.A(G78gat), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n461), .A2(new_n468), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(G22gat), .ZN(new_n474));
  INV_X1    g273(.A(G78gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n461), .A2(new_n468), .A3(new_n469), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT31), .B(G50gat), .ZN(new_n478));
  INV_X1    g277(.A(G106gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n472), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n480), .B1(new_n472), .B2(new_n477), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n423), .A2(new_n452), .A3(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT35), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n472), .A2(new_n477), .ZN(new_n486));
  INV_X1    g285(.A(new_n480), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n477), .A3(new_n480), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n285), .A2(KEYINPUT6), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n490), .B1(new_n285), .B2(new_n287), .ZN(new_n491));
  AND4_X1   g290(.A1(new_n485), .A2(new_n488), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n442), .A2(new_n448), .A3(KEYINPUT74), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT74), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n449), .A2(new_n451), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n422), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n484), .A2(KEYINPUT35), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT95), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n416), .A2(KEYINPUT37), .A3(new_n419), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT94), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n499), .A2(new_n500), .A3(new_n403), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n499), .B2(new_n403), .ZN(new_n502));
  XOR2_X1   g301(.A(KEYINPUT93), .B(KEYINPUT37), .Z(new_n503));
  NAND2_X1  g302(.A1(new_n399), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NOR3_X1   g304(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT38), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n498), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n499), .A2(new_n403), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n505), .B1(new_n509), .B2(KEYINPUT94), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n499), .A2(new_n500), .A3(new_n403), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n512), .A2(KEYINPUT95), .A3(KEYINPUT38), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n364), .A2(new_n389), .A3(new_n393), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n514), .B(KEYINPUT37), .C1(new_n364), .C2(new_n395), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n504), .A2(new_n515), .A3(new_n507), .A4(new_n417), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n516), .A2(new_n406), .A3(new_n408), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n491), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n508), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n262), .A2(new_n267), .A3(new_n268), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n520), .A2(new_n250), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT39), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n278), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n250), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT90), .B1(new_n248), .B2(new_n250), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT90), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n241), .A2(new_n247), .A3(new_n526), .A4(new_n249), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n524), .A2(new_n528), .A3(KEYINPUT39), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n523), .A2(KEYINPUT40), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n285), .B1(new_n530), .B2(KEYINPUT92), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT30), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n420), .A2(new_n421), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT40), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n524), .A2(new_n528), .A3(KEYINPUT39), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n277), .B1(new_n524), .B2(KEYINPUT39), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT91), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT91), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n540), .B(new_n535), .C1(new_n536), .C2(new_n537), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n539), .B(new_n541), .C1(KEYINPUT92), .C2(new_n530), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n488), .A2(new_n489), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI22_X1  g344(.A1(new_n292), .A2(new_n422), .B1(new_n481), .B2(new_n482), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT36), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n495), .A2(new_n547), .A3(new_n493), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n449), .A2(new_n451), .A3(KEYINPUT36), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n519), .A2(new_n545), .B1(new_n551), .B2(KEYINPUT89), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT89), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n546), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n497), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G113gat), .B(G141gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(G197gat), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT11), .B(G169gat), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n559), .B(KEYINPUT12), .Z(new_n560));
  NAND2_X1  g359(.A1(G229gat), .A2(G233gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G15gat), .B(G22gat), .ZN(new_n563));
  OR2_X1    g362(.A1(new_n563), .A2(G1gat), .ZN(new_n564));
  AOI21_X1  g363(.A(G8gat), .B1(new_n564), .B2(KEYINPUT100), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT16), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n563), .B1(new_n566), .B2(G1gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n565), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G43gat), .B(G50gat), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(KEYINPUT15), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT14), .ZN(new_n572));
  OR3_X1    g371(.A1(new_n572), .A2(G29gat), .A3(G36gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(G29gat), .B2(G36gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(KEYINPUT15), .ZN(new_n577));
  NAND2_X1  g376(.A1(G29gat), .A2(G36gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT98), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n580), .A2(KEYINPUT99), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(KEYINPUT99), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT97), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n575), .A2(new_n584), .B1(G29gat), .B2(G36gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n573), .A2(KEYINPUT96), .A3(new_n574), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n577), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g386(.A1(new_n581), .A2(new_n582), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT17), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n587), .A2(new_n583), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n569), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT101), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n588), .A2(new_n590), .ZN(new_n596));
  INV_X1    g395(.A(new_n569), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  OAI211_X1 g398(.A(new_n595), .B(new_n569), .C1(new_n592), .C2(new_n593), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n562), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT18), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n596), .B(new_n597), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n561), .B(KEYINPUT13), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(new_n601), .B2(KEYINPUT18), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n560), .B1(new_n603), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n599), .A2(new_n600), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(new_n561), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT18), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n560), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n612), .A2(new_n613), .A3(new_n602), .A4(new_n606), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n608), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n555), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G190gat), .B(G218gat), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT109), .ZN(new_n619));
  NAND2_X1  g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n621), .A2(KEYINPUT41), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n619), .B(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT7), .ZN(new_n626));
  INV_X1    g425(.A(G85gat), .ZN(new_n627));
  OAI21_X1  g426(.A(G92gat), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G92gat), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n628), .A2(new_n630), .B1(new_n626), .B2(new_n627), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT8), .ZN(new_n632));
  NAND2_X1  g431(.A1(G99gat), .A2(G106gat), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT107), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(new_n634), .B2(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G99gat), .B(G106gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT108), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT108), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n631), .A2(new_n636), .A3(new_n641), .A4(new_n638), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n593), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n644), .B2(new_n591), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n596), .A2(new_n643), .B1(KEYINPUT41), .B2(new_n621), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n625), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n645), .A2(new_n647), .A3(new_n625), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n624), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(new_n623), .A3(new_n648), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT106), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G155gat), .ZN(new_n656));
  XOR2_X1   g455(.A(G183gat), .B(G211gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(G71gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(new_n475), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n661), .A2(KEYINPUT102), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(new_n660), .B2(new_n475), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n662), .B(new_n664), .C1(G71gat), .C2(G78gat), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n661), .A2(KEYINPUT9), .ZN(new_n667));
  XOR2_X1   g466(.A(G57gat), .B(G64gat), .Z(new_n668));
  AOI22_X1  g467(.A1(new_n665), .A2(new_n666), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n669), .B1(new_n666), .B2(new_n665), .ZN(new_n670));
  XNOR2_X1  g469(.A(G71gat), .B(G78gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT105), .ZN(new_n672));
  INV_X1    g471(.A(G57gat), .ZN(new_n673));
  INV_X1    g472(.A(G64gat), .ZN(new_n674));
  OR3_X1    g473(.A1(new_n673), .A2(new_n674), .A3(KEYINPUT104), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n673), .B2(KEYINPUT104), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n672), .A2(new_n667), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT21), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(G231gat), .A2(G233gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n678), .A2(new_n679), .A3(new_n681), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G127gat), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n569), .B1(new_n678), .B2(new_n679), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n683), .A2(new_n226), .A3(new_n684), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n659), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n691), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n689), .A3(new_n658), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n651), .A2(new_n653), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT111), .ZN(new_n698));
  INV_X1    g497(.A(G230gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n309), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n643), .A2(new_n678), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n678), .A2(new_n639), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT10), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n643), .A2(KEYINPUT10), .A3(new_n677), .A4(new_n670), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n700), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n703), .A2(new_n699), .A3(new_n309), .ZN(new_n708));
  XNOR2_X1  g507(.A(G120gat), .B(G148gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(G176gat), .B(G204gat), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n709), .B(new_n710), .Z(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OR3_X1    g511(.A1(new_n707), .A2(new_n708), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n712), .B1(new_n707), .B2(new_n708), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(KEYINPUT110), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n716));
  OAI211_X1 g515(.A(new_n716), .B(new_n712), .C1(new_n707), .C2(new_n708), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n697), .A2(new_n698), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n718), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT111), .B1(new_n720), .B2(new_n696), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n292), .A2(KEYINPUT112), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n292), .A2(KEYINPUT112), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n617), .A2(new_n722), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(G1gat), .ZN(G1324gat));
  NAND3_X1  g527(.A1(new_n617), .A2(new_n422), .A3(new_n722), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT113), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n518), .B1(new_n731), .B2(KEYINPUT95), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n506), .A2(new_n498), .A3(new_n507), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n545), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n551), .A2(KEYINPUT89), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(new_n554), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n292), .A2(new_n422), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n488), .A2(new_n452), .A3(new_n489), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT35), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n492), .A2(new_n496), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n615), .ZN(new_n743));
  INV_X1    g542(.A(new_n722), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n746), .A3(new_n422), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n747), .A3(G8gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT16), .B(G8gat), .Z(new_n749));
  NAND4_X1  g548(.A1(new_n745), .A2(KEYINPUT42), .A3(new_n422), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n730), .A2(new_n747), .ZN(new_n751));
  AOI211_X1 g550(.A(KEYINPUT114), .B(KEYINPUT42), .C1(new_n751), .C2(new_n749), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n746), .B1(new_n745), .B2(new_n422), .ZN(new_n754));
  INV_X1    g553(.A(new_n422), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n743), .A2(KEYINPUT113), .A3(new_n755), .A4(new_n744), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n749), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n753), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n748), .B(new_n750), .C1(new_n752), .C2(new_n759), .ZN(G1325gat));
  INV_X1    g559(.A(G15gat), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n495), .A2(new_n493), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n743), .A2(new_n550), .A3(new_n744), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n761), .B2(new_n764), .ZN(G1326gat));
  NAND2_X1  g564(.A1(new_n745), .A2(new_n544), .ZN(new_n766));
  XNOR2_X1  g565(.A(KEYINPUT43), .B(G22gat), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1327gat));
  NAND2_X1  g567(.A1(new_n651), .A2(new_n653), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n720), .A2(new_n770), .A3(new_n695), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n617), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n726), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n772), .A2(G29gat), .A3(new_n773), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT45), .Z(new_n775));
  AOI21_X1  g574(.A(new_n770), .B1(new_n736), .B2(new_n741), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT115), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n779), .B(KEYINPUT44), .C1(new_n555), .C2(new_n770), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n483), .B1(new_n542), .B2(new_n534), .ZN(new_n781));
  INV_X1    g580(.A(new_n518), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n512), .A2(KEYINPUT38), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n783), .B2(new_n498), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n781), .B1(new_n784), .B2(new_n513), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n741), .B1(new_n785), .B2(new_n551), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n777), .A3(new_n769), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n778), .A2(new_n780), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n720), .A2(new_n695), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n615), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n726), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G29gat), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n775), .A2(new_n794), .ZN(G1328gat));
  NOR2_X1   g594(.A1(new_n755), .A2(G36gat), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n617), .A2(new_n771), .A3(new_n796), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(KEYINPUT116), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(KEYINPUT116), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n798), .A2(KEYINPUT46), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT46), .B1(new_n798), .B2(new_n799), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n792), .A2(new_n422), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G36gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1329gat));
  INV_X1    g604(.A(new_n550), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n806), .A3(new_n791), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G43gat), .ZN(new_n808));
  INV_X1    g607(.A(G43gat), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n617), .A2(new_n809), .A3(new_n762), .A4(new_n771), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT47), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(KEYINPUT47), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1330gat));
  NOR3_X1   g614(.A1(new_n772), .A2(G50gat), .A3(new_n483), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n788), .A2(new_n544), .A3(new_n791), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(G50gat), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT48), .ZN(G1331gat));
  AOI21_X1  g618(.A(new_n551), .B1(new_n519), .B2(new_n545), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n497), .ZN(new_n821));
  NOR4_X1   g620(.A1(new_n821), .A2(new_n615), .A3(new_n696), .A4(new_n718), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n726), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n422), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n825), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n826));
  XOR2_X1   g625(.A(KEYINPUT49), .B(G64gat), .Z(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n825), .B2(new_n827), .ZN(G1333gat));
  AOI21_X1  g627(.A(new_n660), .B1(new_n822), .B2(new_n806), .ZN(new_n829));
  AOI21_X1  g628(.A(G71gat), .B1(new_n495), .B2(new_n493), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n822), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g631(.A1(new_n822), .A2(new_n544), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(G78gat), .ZN(G1335gat));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n836), .B(new_n769), .C1(new_n820), .C2(new_n497), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n615), .A2(new_n695), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n836), .B1(new_n786), .B2(new_n769), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT117), .B1(new_n821), .B2(new_n770), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n842), .A2(KEYINPUT51), .A3(new_n838), .A4(new_n837), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n844), .A2(new_n627), .A3(new_n720), .A4(new_n726), .ZN(new_n845));
  INV_X1    g644(.A(new_n838), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n846), .A2(new_n718), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n788), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n726), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n845), .B1(new_n849), .B2(new_n627), .ZN(G1336gat));
  NOR2_X1   g649(.A1(new_n755), .A2(new_n629), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n788), .A2(new_n847), .A3(new_n851), .ZN(new_n852));
  OR2_X1    g651(.A1(KEYINPUT118), .A2(KEYINPUT52), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n720), .A2(new_n422), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n841), .B2(new_n843), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n852), .B(new_n853), .C1(new_n855), .C2(G92gat), .ZN(new_n856));
  NAND2_X1  g655(.A1(KEYINPUT118), .A2(KEYINPUT52), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT119), .Z(new_n858));
  XNOR2_X1  g657(.A(new_n856), .B(new_n858), .ZN(G1337gat));
  NAND2_X1  g658(.A1(new_n848), .A2(new_n806), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(G99gat), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n720), .A2(new_n762), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(G99gat), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n844), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(G1338gat));
  NAND3_X1  g664(.A1(new_n788), .A2(new_n544), .A3(new_n847), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G106gat), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n844), .A2(new_n479), .A3(new_n544), .A4(new_n720), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT53), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n867), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(G1339gat));
  NAND4_X1  g672(.A1(new_n697), .A2(new_n608), .A3(new_n614), .A4(new_n718), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT120), .ZN(new_n875));
  INV_X1    g674(.A(new_n695), .ZN(new_n876));
  OAI22_X1  g675(.A1(new_n609), .A2(new_n561), .B1(new_n604), .B2(new_n605), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n559), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n614), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n707), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n705), .A2(new_n700), .A3(new_n706), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n711), .B1(new_n707), .B2(new_n880), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT55), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n883), .A2(KEYINPUT55), .A3(new_n884), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n887), .A2(new_n713), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n769), .B1(new_n879), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n770), .B1(new_n879), .B2(new_n718), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n608), .B2(new_n614), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n876), .B(new_n890), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n738), .ZN(new_n895));
  AND4_X1   g694(.A1(new_n755), .A2(new_n894), .A3(new_n895), .A4(new_n726), .ZN(new_n896));
  AOI21_X1  g695(.A(G113gat), .B1(new_n896), .B2(new_n615), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n544), .B1(new_n875), .B2(new_n893), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n496), .A3(new_n726), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n899), .A2(new_n233), .A3(new_n616), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n897), .A2(new_n900), .ZN(G1340gat));
  AOI21_X1  g700(.A(G120gat), .B1(new_n896), .B2(new_n720), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n899), .A2(new_n231), .A3(new_n718), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(G1341gat));
  NAND3_X1  g703(.A1(new_n896), .A2(new_n226), .A3(new_n695), .ZN(new_n905));
  OAI21_X1  g704(.A(G127gat), .B1(new_n899), .B2(new_n876), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1342gat));
  NAND3_X1  g706(.A1(new_n896), .A2(new_n224), .A3(new_n769), .ZN(new_n908));
  XOR2_X1   g707(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n909));
  XNOR2_X1  g708(.A(new_n908), .B(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G134gat), .B1(new_n899), .B2(new_n770), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1343gat));
  NOR3_X1   g711(.A1(new_n773), .A2(new_n422), .A3(new_n806), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n483), .B1(new_n875), .B2(new_n893), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT57), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n914), .A2(KEYINPUT57), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n220), .B1(new_n918), .B2(new_n616), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT58), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n894), .A2(new_n544), .ZN(new_n922));
  INV_X1    g721(.A(new_n913), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n616), .A2(G141gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n919), .A2(new_n920), .A3(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n220), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT57), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n922), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n923), .B1(new_n930), .B2(new_n915), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n931), .B2(new_n615), .ZN(new_n932));
  INV_X1    g731(.A(new_n926), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT58), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n927), .A2(new_n934), .ZN(G1344gat));
  NAND3_X1  g734(.A1(new_n924), .A2(new_n212), .A3(new_n720), .ZN(new_n936));
  AOI211_X1 g735(.A(KEYINPUT59), .B(new_n212), .C1(new_n931), .C2(new_n720), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n722), .A2(new_n616), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n483), .B1(new_n939), .B2(new_n893), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n915), .B1(KEYINPUT57), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(new_n720), .A3(new_n913), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n938), .B1(new_n942), .B2(G148gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n936), .B1(new_n937), .B2(new_n943), .ZN(G1345gat));
  OAI21_X1  g743(.A(G155gat), .B1(new_n918), .B2(new_n876), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n924), .A2(new_n206), .A3(new_n695), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1346gat));
  NAND3_X1  g746(.A1(new_n924), .A2(new_n207), .A3(new_n769), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n769), .B(new_n913), .C1(new_n916), .C2(new_n917), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT123), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G162gat), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n949), .A2(KEYINPUT123), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(G1347gat));
  NOR2_X1   g752(.A1(new_n726), .A2(new_n755), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n898), .A2(new_n762), .A3(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(G169gat), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n955), .A2(new_n956), .A3(new_n616), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT124), .B1(new_n894), .B2(new_n773), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n958), .A2(new_n755), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n894), .A2(KEYINPUT124), .A3(new_n773), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n895), .A3(new_n960), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n961), .A2(new_n616), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n957), .B1(new_n962), .B2(new_n956), .ZN(G1348gat));
  OR2_X1    g762(.A1(new_n961), .A2(new_n718), .ZN(new_n964));
  INV_X1    g763(.A(G176gat), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n898), .A2(new_n954), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n862), .A2(new_n965), .ZN(new_n967));
  AOI22_X1  g766(.A1(new_n964), .A2(new_n965), .B1(new_n966), .B2(new_n967), .ZN(G1349gat));
  OAI21_X1  g767(.A(G183gat), .B1(new_n955), .B2(new_n876), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n695), .A2(new_n300), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n961), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(KEYINPUT60), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT60), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n973), .B(new_n969), .C1(new_n961), .C2(new_n970), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1350gat));
  NOR2_X1   g774(.A1(new_n770), .A2(G190gat), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n959), .A2(new_n895), .A3(new_n960), .A4(new_n976), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n898), .A2(new_n762), .A3(new_n769), .A4(new_n954), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT61), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n978), .A2(new_n979), .A3(G190gat), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n979), .B1(new_n978), .B2(G190gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(KEYINPUT125), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT125), .ZN(new_n984));
  OAI211_X1 g783(.A(new_n977), .B(new_n984), .C1(new_n980), .C2(new_n981), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(new_n985), .ZN(G1351gat));
  NOR2_X1   g785(.A1(new_n806), .A2(new_n483), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n959), .A2(new_n960), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n615), .A2(new_n370), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n988), .A2(KEYINPUT126), .A3(new_n989), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n726), .A2(new_n755), .A3(new_n806), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n941), .A2(new_n615), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n992), .B1(new_n994), .B2(G197gat), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n990), .B1(new_n991), .B2(new_n995), .ZN(G1352gat));
  NAND3_X1  g795(.A1(new_n941), .A2(new_n720), .A3(new_n993), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n941), .A2(KEYINPUT127), .A3(new_n720), .A4(new_n993), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n999), .A2(G204gat), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n720), .A2(new_n379), .ZN(new_n1002));
  OR3_X1    g801(.A1(new_n988), .A2(KEYINPUT62), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g802(.A(KEYINPUT62), .B1(new_n988), .B2(new_n1002), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(G1353gat));
  NAND3_X1  g804(.A1(new_n941), .A2(new_n695), .A3(new_n993), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n1006), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1007));
  AOI21_X1  g806(.A(KEYINPUT63), .B1(new_n1006), .B2(G211gat), .ZN(new_n1008));
  OR2_X1    g807(.A1(new_n876), .A2(G211gat), .ZN(new_n1009));
  OAI22_X1  g808(.A1(new_n1007), .A2(new_n1008), .B1(new_n988), .B2(new_n1009), .ZN(G1354gat));
  NAND3_X1  g809(.A1(new_n941), .A2(new_n769), .A3(new_n993), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1011), .A2(G218gat), .ZN(new_n1012));
  OR2_X1    g811(.A1(new_n770), .A2(G218gat), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1012), .B1(new_n988), .B2(new_n1013), .ZN(G1355gat));
endmodule


