//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT16), .ZN(new_n193));
  OR3_X1    g007(.A1(new_n191), .A2(KEYINPUT16), .A3(G140), .ZN(new_n194));
  AOI21_X1  g008(.A(G146), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n194), .A3(G146), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(KEYINPUT69), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT69), .ZN(new_n199));
  AND4_X1   g013(.A1(new_n199), .A2(new_n193), .A3(G146), .A4(new_n194), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n202), .B(G119), .C1(KEYINPUT68), .C2(KEYINPUT23), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G128), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n207), .B1(new_n205), .B2(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n203), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G119), .B(G128), .ZN(new_n210));
  XOR2_X1   g024(.A(KEYINPUT24), .B(G110), .Z(new_n211));
  AOI22_X1  g025(.A1(new_n209), .A2(G110), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n198), .A2(new_n201), .A3(new_n212), .ZN(new_n213));
  OAI22_X1  g027(.A1(new_n209), .A2(G110), .B1(new_n210), .B2(new_n211), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n190), .A2(new_n192), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n197), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G953), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(G221), .A3(G234), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n221), .B(KEYINPUT70), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G137), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n219), .B(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G902), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n188), .B1(new_n227), .B2(KEYINPUT25), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n228), .B1(KEYINPUT25), .B2(new_n227), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n188), .A2(new_n226), .ZN(new_n230));
  XOR2_X1   g044(.A(new_n230), .B(KEYINPUT71), .Z(new_n231));
  NAND2_X1  g045(.A1(new_n225), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G143), .B(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT0), .B(G128), .Z(new_n237));
  OAI21_X1  g051(.A(new_n236), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G131), .ZN(new_n239));
  INV_X1    g053(.A(G134), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT64), .B1(new_n240), .B2(G137), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT11), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  OAI211_X1 g057(.A(KEYINPUT64), .B(new_n243), .C1(new_n240), .C2(G137), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n245), .A2(G134), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  AND4_X1   g061(.A1(new_n239), .A2(new_n242), .A3(new_n244), .A4(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n246), .B1(new_n241), .B2(KEYINPUT11), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n239), .B1(new_n249), .B2(new_n244), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT65), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n248), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n242), .A2(new_n244), .A3(new_n247), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G131), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n249), .A2(new_n239), .A3(new_n244), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT65), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n238), .B1(new_n252), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n216), .A2(G143), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n202), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(new_n259), .A3(new_n260), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n258), .A2(KEYINPUT1), .A3(G146), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n240), .A2(G137), .ZN(new_n267));
  OAI21_X1  g081(.A(G131), .B1(new_n267), .B2(new_n246), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n255), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n257), .A2(KEYINPUT30), .A3(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT2), .B(G113), .Z(new_n271));
  INV_X1    g085(.A(G116), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n205), .ZN(new_n273));
  NAND2_X1  g087(.A1(G116), .A2(G119), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT2), .B(G113), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n273), .A3(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT30), .ZN(new_n280));
  INV_X1    g094(.A(new_n238), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(new_n254), .B2(new_n255), .ZN(new_n282));
  INV_X1    g096(.A(new_n269), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n270), .A2(new_n279), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT31), .ZN(new_n286));
  XNOR2_X1  g100(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n287));
  NOR2_X1   g101(.A1(G237), .A2(G953), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G210), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n287), .B(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(G101), .ZN(new_n291));
  XOR2_X1   g105(.A(new_n290), .B(new_n291), .Z(new_n292));
  OAI21_X1  g106(.A(new_n251), .B1(new_n248), .B2(new_n250), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n254), .A2(KEYINPUT65), .A3(new_n255), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n283), .B1(new_n295), .B2(new_n238), .ZN(new_n296));
  INV_X1    g110(.A(new_n279), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n292), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n285), .A2(new_n286), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT67), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n285), .A2(new_n301), .A3(new_n298), .A4(new_n286), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n285), .A2(new_n298), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n257), .A2(new_n297), .A3(new_n269), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n296), .A2(KEYINPUT28), .A3(new_n297), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI22_X1  g124(.A1(KEYINPUT31), .A2(new_n304), .B1(new_n310), .B2(new_n292), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n303), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(G472), .A2(G902), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT32), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT32), .ZN(new_n315));
  INV_X1    g129(.A(new_n313), .ZN(new_n316));
  AOI211_X1 g130(.A(new_n315), .B(new_n316), .C1(new_n303), .C2(new_n311), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n292), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n310), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n319), .B1(new_n296), .B2(new_n297), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n285), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT29), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n257), .A2(new_n269), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(new_n279), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n307), .A2(new_n309), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(KEYINPUT29), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n226), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(G472), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n233), .B1(new_n318), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT87), .ZN(new_n331));
  NOR2_X1   g145(.A1(G475), .A2(G902), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT85), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n193), .A2(G146), .A3(new_n194), .ZN(new_n335));
  NOR3_X1   g149(.A1(new_n335), .A2(new_n195), .A3(new_n199), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n334), .B1(new_n336), .B2(new_n200), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT17), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n288), .A2(G214), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(new_n258), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n288), .B(G214), .C1(KEYINPUT83), .C2(G143), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n341), .A2(new_n239), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n239), .B1(new_n341), .B2(new_n342), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n341), .A2(new_n342), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT17), .B1(new_n346), .B2(new_n239), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n198), .A2(new_n201), .A3(KEYINPUT85), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n337), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(G113), .B(G122), .ZN(new_n351));
  INV_X1    g165(.A(G104), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT18), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n346), .B1(new_n354), .B2(new_n239), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n341), .A2(new_n342), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT18), .A3(G131), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n215), .B(new_n216), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n350), .A2(new_n353), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT84), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n361), .A2(KEYINPUT19), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(KEYINPUT19), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n190), .B(new_n192), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n215), .B2(new_n363), .ZN(new_n365));
  OAI221_X1 g179(.A(new_n197), .B1(new_n365), .B2(G146), .C1(new_n344), .C2(new_n343), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n359), .ZN(new_n367));
  INV_X1    g181(.A(new_n353), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n333), .B1(new_n360), .B2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n370), .A2(KEYINPUT86), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n372));
  AOI211_X1 g186(.A(new_n372), .B(new_n333), .C1(new_n360), .C2(new_n369), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n360), .A2(new_n369), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n372), .B(new_n374), .C1(new_n376), .C2(new_n333), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n350), .A2(new_n353), .A3(new_n359), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n353), .B1(new_n350), .B2(new_n359), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n226), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G475), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n331), .B1(new_n375), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G475), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n350), .A2(new_n359), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(new_n368), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n360), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n384), .B1(new_n387), .B2(new_n226), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n370), .A2(KEYINPUT86), .A3(KEYINPUT20), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n374), .B1(new_n370), .B2(KEYINPUT86), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n391), .B1(KEYINPUT86), .B2(new_n370), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(KEYINPUT87), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(KEYINPUT9), .B(G234), .ZN(new_n394));
  INV_X1    g208(.A(G217), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n394), .A2(new_n395), .A3(G953), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n272), .A2(G122), .ZN(new_n397));
  INV_X1    g211(.A(G122), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(G116), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(G107), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(KEYINPUT88), .B1(new_n202), .B2(G143), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n258), .A3(G128), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n202), .A2(G143), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n240), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n240), .B1(new_n406), .B2(new_n407), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT14), .B1(new_n398), .B2(G116), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT90), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n397), .B1(new_n413), .B2(new_n399), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI221_X1 g229(.A(new_n402), .B1(new_n409), .B2(new_n410), .C1(new_n415), .C2(new_n401), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n400), .B(new_n401), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT13), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n407), .B1(new_n406), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n406), .A2(new_n418), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT89), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT89), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n406), .A2(new_n422), .A3(new_n418), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n419), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n408), .B(new_n417), .C1(new_n424), .C2(new_n240), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n396), .B1(new_n416), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n416), .A2(new_n425), .A3(new_n396), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT92), .A3(new_n226), .ZN(new_n430));
  INV_X1    g244(.A(G478), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT15), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(KEYINPUT91), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(KEYINPUT91), .B2(new_n432), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(G902), .B1(new_n427), .B2(new_n428), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(KEYINPUT92), .A3(new_n434), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(G234), .A2(G237), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n440), .A2(G952), .A3(new_n220), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT21), .B(G898), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT93), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n440), .A2(G902), .A3(G953), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n442), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n439), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n383), .A2(new_n393), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G214), .B1(G237), .B2(G902), .ZN(new_n451));
  OAI21_X1  g265(.A(G210), .B1(G237), .B2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G110), .B(G122), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT77), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(KEYINPUT8), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT5), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n273), .B2(new_n274), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n205), .A3(G116), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G113), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n276), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(KEYINPUT3), .B1(new_n352), .B2(G107), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n463), .A2(new_n401), .A3(G104), .ZN(new_n464));
  INV_X1    g278(.A(G101), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n352), .A2(G107), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n462), .A2(new_n464), .A3(new_n465), .A4(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n352), .A2(G107), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n401), .A2(G104), .ZN(new_n469));
  OAI21_X1  g283(.A(G101), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n461), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n467), .A2(new_n470), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n458), .A2(new_n460), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n276), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n461), .A2(new_n471), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT81), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n456), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n462), .A2(new_n464), .A3(new_n466), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n481), .A2(KEYINPUT73), .A3(G101), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT73), .B1(new_n481), .B2(G101), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n467), .A2(KEYINPUT4), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT4), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n481), .A2(new_n486), .A3(G101), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n279), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n455), .B(new_n475), .C1(new_n485), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT79), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n236), .B(G125), .C1(new_n234), .C2(new_n237), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n262), .A2(new_n191), .A3(new_n264), .A4(new_n265), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G224), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(G953), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n491), .A2(new_n490), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n494), .A2(KEYINPUT7), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n491), .A2(new_n492), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT7), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(new_n496), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n480), .A2(new_n489), .A3(new_n499), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n226), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n481), .A2(G101), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT73), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n481), .A2(KEYINPUT73), .A3(G101), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n507), .A2(KEYINPUT4), .A3(new_n508), .A4(new_n467), .ZN(new_n509));
  INV_X1    g323(.A(new_n488), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n478), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n455), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT78), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n489), .B(KEYINPUT6), .C1(new_n511), .C2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n516));
  INV_X1    g330(.A(new_n498), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n496), .B1(new_n517), .B2(new_n493), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n475), .B1(new_n485), .B2(new_n488), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT6), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n520), .A2(new_n513), .A3(new_n521), .A4(new_n512), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n515), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT80), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n515), .A2(new_n519), .A3(KEYINPUT80), .A4(new_n522), .ZN(new_n526));
  AOI211_X1 g340(.A(new_n453), .B(new_n504), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  INV_X1    g342(.A(new_n504), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n452), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n451), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT82), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g347(.A(KEYINPUT82), .B(new_n451), .C1(new_n527), .C2(new_n530), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n450), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n220), .A2(G227), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(G140), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT72), .B(G110), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT10), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n471), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n473), .A2(KEYINPUT10), .A3(new_n266), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n238), .A2(new_n487), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n543), .B(new_n544), .C1(new_n485), .C2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT74), .B1(new_n546), .B2(new_n295), .ZN(new_n547));
  INV_X1    g361(.A(new_n295), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n473), .A2(KEYINPUT10), .A3(new_n266), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT10), .B1(new_n473), .B2(new_n266), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n509), .A2(new_n238), .A3(new_n487), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT74), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n548), .A2(new_n551), .A3(new_n552), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n473), .A2(new_n266), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n471), .A2(new_n264), .A3(new_n265), .A4(new_n262), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT12), .B1(new_n248), .B2(new_n250), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n295), .A2(new_n559), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT12), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n563), .A2(KEYINPUT75), .A3(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT75), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n293), .A2(new_n294), .B1(new_n557), .B2(new_n558), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n566), .B1(new_n567), .B2(KEYINPUT12), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n562), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n540), .B1(new_n556), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n555), .A2(KEYINPUT76), .A3(new_n539), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n546), .A2(new_n295), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n540), .B1(new_n547), .B2(new_n554), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n574), .A2(KEYINPUT76), .ZN(new_n575));
  OAI211_X1 g389(.A(G469), .B(new_n570), .C1(new_n573), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n555), .A2(new_n539), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n547), .A2(new_n554), .B1(new_n295), .B2(new_n546), .ZN(new_n578));
  OAI22_X1  g392(.A1(new_n577), .A2(new_n569), .B1(new_n578), .B2(new_n539), .ZN(new_n579));
  INV_X1    g393(.A(G469), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n226), .ZN(new_n581));
  NAND2_X1  g395(.A1(G469), .A2(G902), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n576), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(G221), .B1(new_n394), .B2(G902), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n330), .A2(new_n535), .A3(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n383), .A2(new_n393), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n437), .A2(G478), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT33), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n429), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT33), .B1(new_n427), .B2(new_n428), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n431), .A2(G902), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n528), .A2(new_n529), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n453), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n528), .A2(new_n452), .A3(new_n529), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(KEYINPUT94), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n451), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n604), .B1(new_n527), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n603), .A2(new_n447), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n589), .B1(new_n599), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n451), .B1(new_n602), .B2(KEYINPUT94), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n527), .A2(new_n530), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(KEYINPUT94), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n597), .B1(new_n383), .B2(new_n393), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n611), .A2(new_n612), .A3(KEYINPUT95), .A4(new_n447), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n312), .A2(new_n313), .ZN(new_n615));
  INV_X1    g429(.A(G472), .ZN(new_n616));
  AOI21_X1  g430(.A(G902), .B1(new_n303), .B2(new_n311), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n618), .A2(new_n585), .A3(new_n233), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT96), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT34), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G104), .ZN(G6));
  NAND3_X1  g437(.A1(new_n390), .A2(new_n439), .A3(new_n392), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n607), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G107), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  NOR2_X1   g442(.A1(new_n618), .A2(new_n585), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n533), .A2(new_n534), .ZN(new_n630));
  INV_X1    g444(.A(new_n450), .ZN(new_n631));
  INV_X1    g445(.A(new_n224), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(new_n219), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n231), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n229), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n629), .A2(new_n630), .A3(new_n631), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT37), .B(G110), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G12));
  NAND2_X1  g453(.A1(new_n615), .A2(new_n315), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n312), .A2(KEYINPUT32), .A3(new_n313), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n329), .A3(new_n641), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n642), .A2(new_n586), .A3(new_n636), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n375), .A2(new_n382), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT97), .B(G900), .Z(new_n646));
  AOI21_X1  g460(.A(new_n441), .B1(new_n646), .B2(new_n445), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n644), .A2(new_n645), .A3(new_n439), .A4(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT98), .B1(new_n624), .B2(new_n647), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n611), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT99), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n611), .A2(new_n650), .A3(new_n649), .A4(KEYINPUT99), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n643), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT100), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  XNOR2_X1  g471(.A(new_n610), .B(KEYINPUT101), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n658), .A2(KEYINPUT38), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(KEYINPUT38), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n285), .A2(new_n305), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n319), .ZN(new_n663));
  AOI21_X1  g477(.A(G902), .B1(new_n321), .B2(new_n325), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n616), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n314), .A2(new_n317), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n647), .B(KEYINPUT39), .Z(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n585), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT40), .ZN(new_n674));
  INV_X1    g488(.A(new_n439), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n383), .B2(new_n393), .ZN(new_n676));
  INV_X1    g490(.A(new_n636), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n676), .A2(new_n451), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n661), .A2(new_n670), .A3(new_n674), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  NAND3_X1  g494(.A1(new_n611), .A2(new_n612), .A3(new_n648), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n643), .A2(new_n682), .A3(KEYINPUT103), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n642), .A2(new_n586), .A3(new_n636), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n684), .B1(new_n685), .B2(new_n681), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  INV_X1    g502(.A(new_n233), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT104), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n580), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n555), .A2(new_n572), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT75), .B1(new_n563), .B2(new_n564), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n567), .A2(new_n566), .A3(KEYINPUT12), .ZN(new_n694));
  OAI22_X1  g508(.A1(new_n693), .A2(new_n694), .B1(new_n560), .B2(new_n561), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n540), .A2(new_n692), .B1(new_n695), .B2(new_n574), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n691), .B1(new_n696), .B2(G902), .ZN(new_n697));
  INV_X1    g511(.A(new_n691), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n579), .A2(new_n226), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n697), .A2(new_n699), .A3(new_n584), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n642), .A2(new_n689), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n608), .B2(new_n613), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g519(.A(KEYINPUT41), .B(G113), .Z(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT106), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n705), .B(new_n707), .ZN(G15));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n611), .A2(new_n644), .A3(new_n439), .A4(new_n447), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n709), .B1(new_n702), .B2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n330), .A2(new_n625), .A3(KEYINPUT107), .A4(new_n701), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT108), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n272), .ZN(G18));
  NOR3_X1   g529(.A1(new_n527), .A2(new_n530), .A3(new_n605), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n716), .A2(new_n700), .A3(new_n609), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n642), .A3(new_n631), .A4(new_n636), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  NOR2_X1   g533(.A1(new_n617), .A2(new_n616), .ZN(new_n720));
  AOI22_X1  g534(.A1(KEYINPUT31), .A2(new_n304), .B1(new_n326), .B2(new_n292), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n316), .B1(new_n303), .B2(new_n721), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n720), .A2(new_n722), .A3(new_n233), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n700), .A2(new_n448), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(new_n676), .A3(new_n611), .A4(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NAND2_X1  g540(.A1(new_n303), .A2(new_n721), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n313), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n728), .B(new_n636), .C1(new_n616), .C2(new_n617), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT109), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n312), .A2(new_n226), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G472), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT109), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n636), .A4(new_n728), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n375), .A2(new_n382), .A3(new_n331), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT87), .B1(new_n390), .B2(new_n392), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n598), .B(new_n648), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n692), .A2(new_n540), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n695), .A2(new_n574), .ZN(new_n740));
  AOI211_X1 g554(.A(G902), .B(new_n691), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n698), .B1(new_n579), .B2(new_n226), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n603), .A2(new_n743), .A3(new_n606), .A4(new_n584), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n735), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT110), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n735), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  AOI211_X1 g565(.A(new_n647), .B(new_n597), .C1(new_n383), .C2(new_n393), .ZN(new_n752));
  AND4_X1   g566(.A1(new_n584), .A2(new_n610), .A3(new_n583), .A4(new_n451), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n752), .A2(new_n753), .A3(new_n642), .A4(new_n689), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(KEYINPUT42), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n756), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n330), .A2(new_n752), .A3(new_n758), .A4(new_n753), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G131), .ZN(G33));
  NAND4_X1  g575(.A1(new_n330), .A2(new_n649), .A3(new_n650), .A4(new_n753), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT112), .B(G134), .Z(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G36));
  OAI21_X1  g578(.A(new_n570), .B1(new_n573), .B2(new_n575), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n766));
  OR2_X1    g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT114), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n765), .A2(new_n766), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(KEYINPUT113), .A3(G469), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT113), .B1(new_n769), .B2(G469), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n582), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(KEYINPUT46), .B(new_n582), .C1(new_n771), .C2(new_n772), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n581), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n584), .A3(new_n671), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n590), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n598), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n781), .A2(KEYINPUT43), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(KEYINPUT43), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n677), .B1(new_n732), .B2(new_n615), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(KEYINPUT44), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n527), .A2(new_n530), .A3(new_n604), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(KEYINPUT115), .Z(new_n791));
  NAND3_X1  g605(.A1(new_n786), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n779), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  NAND2_X1  g609(.A1(new_n777), .A2(new_n584), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT47), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n777), .A2(new_n798), .A3(new_n584), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n790), .A2(new_n233), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n738), .A2(new_n642), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  AND2_X1   g617(.A1(new_n723), .A2(new_n441), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n782), .A2(new_n783), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n799), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n798), .B1(new_n777), .B2(new_n584), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n743), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n584), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n791), .B(new_n806), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n670), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n701), .A2(new_n441), .A3(new_n790), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n814), .A2(new_n689), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n813), .A2(new_n815), .A3(KEYINPUT122), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n780), .A3(new_n597), .A4(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n784), .A2(new_n735), .A3(new_n814), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n700), .A2(new_n451), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n824), .B1(new_n659), .B2(new_n660), .ZN(new_n825));
  AND2_X1   g639(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n826));
  OR3_X1    g640(.A1(new_n805), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n828));
  OAI211_X1 g642(.A(KEYINPUT120), .B(KEYINPUT50), .C1(new_n805), .C2(new_n825), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n828), .B1(new_n827), .B2(new_n829), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n822), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT51), .B1(new_n812), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n818), .A2(new_n612), .A3(new_n819), .ZN(new_n834));
  OAI211_X1 g648(.A(G952), .B(new_n220), .C1(new_n805), .C2(new_n744), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n784), .A2(new_n814), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n642), .A2(new_n689), .ZN(new_n837));
  OR3_X1    g651(.A1(new_n836), .A2(KEYINPUT48), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT48), .B1(new_n836), .B2(new_n837), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n806), .A2(new_n791), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n797), .A2(new_n799), .ZN(new_n842));
  INV_X1    g656(.A(new_n811), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n827), .A2(new_n829), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(KEYINPUT51), .A3(new_n821), .A4(new_n820), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n834), .B(new_n840), .C1(new_n844), .C2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n833), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n383), .A2(new_n393), .A3(new_n439), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n599), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n448), .B1(new_n533), .B2(new_n534), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n851), .A2(new_n619), .A3(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n587), .A2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n637), .A2(new_n718), .A3(new_n725), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n713), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n738), .B1(new_n730), .B2(new_n734), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n644), .A2(new_n675), .A3(new_n648), .ZN(new_n858));
  AOI211_X1 g672(.A(new_n677), .B(new_n858), .C1(new_n318), .C2(new_n329), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n753), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n760), .A2(new_n860), .A3(new_n762), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n705), .A2(new_n856), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n586), .A2(new_n677), .A3(new_n648), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n611), .A2(new_n676), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n864), .A2(new_n865), .A3(new_n666), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT103), .B1(new_n643), .B2(new_n682), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n685), .A2(new_n681), .A3(new_n684), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n735), .A2(new_n745), .A3(new_n748), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n748), .B1(new_n735), .B2(new_n745), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n655), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n863), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n866), .B1(new_n683), .B2(new_n686), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(new_n750), .A3(KEYINPUT52), .A4(new_n655), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT117), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n750), .A3(new_n655), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n878), .B1(new_n879), .B2(new_n863), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n849), .B(new_n862), .C1(new_n877), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n874), .A2(new_n876), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n862), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT53), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n881), .A2(KEYINPUT54), .A3(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT118), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n881), .A2(new_n884), .A3(KEYINPUT118), .A4(KEYINPUT54), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n862), .B1(new_n877), .B2(new_n880), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT53), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n882), .A2(new_n849), .A3(new_n862), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n893), .B1(new_n891), .B2(KEYINPUT53), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n898), .A2(KEYINPUT119), .A3(KEYINPUT54), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n848), .B(new_n889), .C1(new_n897), .C2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(G952), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n220), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n810), .A2(KEYINPUT49), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(KEYINPUT116), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(KEYINPUT116), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n689), .A2(new_n584), .A3(new_n451), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n908), .B1(KEYINPUT49), .B2(new_n810), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  OR4_X1    g724(.A1(new_n670), .A2(new_n910), .A3(new_n661), .A4(new_n781), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n903), .A2(new_n911), .ZN(G75));
  NOR2_X1   g726(.A1(new_n220), .A2(G952), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n895), .A2(new_n226), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT56), .B1(new_n915), .B2(G210), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n515), .A2(new_n522), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT123), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT55), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(new_n519), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n914), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  AOI211_X1 g736(.A(KEYINPUT56), .B(new_n920), .C1(new_n915), .C2(G210), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(G51));
  XOR2_X1   g738(.A(new_n582), .B(KEYINPUT57), .Z(new_n925));
  NOR2_X1   g739(.A1(new_n895), .A2(new_n896), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n898), .A2(KEYINPUT54), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n579), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n771), .A2(new_n772), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n915), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n913), .B1(new_n929), .B2(new_n931), .ZN(G54));
  NAND3_X1  g746(.A1(new_n915), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n376), .ZN(new_n934));
  INV_X1    g748(.A(new_n376), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n915), .A2(KEYINPUT58), .A3(G475), .A4(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n934), .A2(new_n914), .A3(new_n936), .ZN(G60));
  INV_X1    g751(.A(new_n595), .ZN(new_n938));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  NOR2_X1   g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n941), .B1(new_n926), .B2(new_n927), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n914), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n889), .B1(new_n897), .B2(new_n899), .ZN(new_n944));
  INV_X1    g758(.A(new_n940), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n943), .B1(new_n946), .B2(new_n938), .ZN(G63));
  NAND2_X1  g761(.A1(G217), .A2(G902), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT60), .Z(new_n949));
  NAND3_X1  g763(.A1(new_n898), .A2(new_n634), .A3(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n898), .A2(new_n949), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n914), .B(new_n950), .C1(new_n951), .C2(new_n225), .ZN(new_n952));
  XNOR2_X1  g766(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n952), .B(new_n954), .ZN(G66));
  AOI21_X1  g769(.A(new_n220), .B1(new_n444), .B2(G224), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n705), .A2(new_n856), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT125), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n958), .B2(new_n220), .ZN(new_n959));
  INV_X1    g773(.A(G898), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n918), .B1(new_n960), .B2(G953), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n959), .B(new_n961), .ZN(G69));
  NAND2_X1  g776(.A1(new_n270), .A2(new_n284), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(new_n365), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n778), .A2(new_n837), .A3(new_n865), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n760), .A2(new_n762), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n778), .B2(new_n792), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n873), .B1(new_n686), .B2(new_n683), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n965), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(G953), .B1(new_n970), .B2(new_n802), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n220), .A2(G900), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n964), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n968), .A2(new_n679), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n974), .A2(KEYINPUT62), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n330), .A2(new_n851), .A3(new_n671), .A4(new_n753), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n778), .B2(new_n792), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n974), .A2(KEYINPUT62), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n975), .A2(new_n978), .A3(new_n802), .A4(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT126), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n977), .B1(new_n809), .B2(new_n801), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n983), .A2(KEYINPUT126), .A3(new_n975), .A4(new_n979), .ZN(new_n984));
  AOI21_X1  g798(.A(G953), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n973), .B1(new_n985), .B2(new_n964), .ZN(new_n986));
  INV_X1    g800(.A(G227), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n972), .B1(new_n987), .B2(G953), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT127), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n989), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n973), .B(new_n991), .C1(new_n985), .C2(new_n964), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(G72));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  NAND2_X1  g809(.A1(new_n970), .A2(new_n802), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n996), .B2(new_n958), .ZN(new_n997));
  INV_X1    g811(.A(new_n322), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n663), .A2(new_n322), .A3(new_n995), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n881), .A2(new_n884), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n999), .A2(new_n914), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n663), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n982), .A2(new_n984), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n995), .B1(new_n1004), .B2(new_n958), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1002), .B1(new_n1003), .B2(new_n1005), .ZN(G57));
endmodule


