

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U560 ( .A1(n534), .A2(G2104), .ZN(n882) );
  NOR2_X1 U561 ( .A1(n702), .A2(n701), .ZN(n700) );
  NOR2_X1 U562 ( .A1(G651), .A2(G543), .ZN(n649) );
  AND2_X1 U563 ( .A1(n818), .A2(n833), .ZN(n526) );
  NOR2_X1 U564 ( .A1(n783), .A2(n765), .ZN(n527) );
  NOR2_X1 U565 ( .A1(n747), .A2(n934), .ZN(n703) );
  NOR2_X1 U566 ( .A1(n986), .A2(n706), .ZN(n707) );
  XNOR2_X1 U567 ( .A(n695), .B(n747), .ZN(n723) );
  XNOR2_X1 U568 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n738) );
  XNOR2_X1 U569 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U570 ( .A1(G2084), .A2(n747), .ZN(n694) );
  INV_X1 U571 ( .A(KEYINPUT101), .ZN(n776) );
  NAND2_X1 U572 ( .A1(n693), .A2(n799), .ZN(n747) );
  NOR2_X1 U573 ( .A1(n819), .A2(n526), .ZN(n820) );
  NOR2_X1 U574 ( .A1(G651), .A2(n636), .ZN(n647) );
  XNOR2_X1 U575 ( .A(KEYINPUT72), .B(n590), .ZN(n711) );
  XOR2_X1 U576 ( .A(KEYINPUT1), .B(n554), .Z(n650) );
  NAND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XNOR2_X2 U578 ( .A(n528), .B(KEYINPUT65), .ZN(n886) );
  NAND2_X1 U579 ( .A1(G113), .A2(n886), .ZN(n529) );
  XNOR2_X1 U580 ( .A(n529), .B(KEYINPUT66), .ZN(n532) );
  INV_X1 U581 ( .A(G2105), .ZN(n534) );
  NAND2_X1 U582 ( .A1(G101), .A2(n882), .ZN(n530) );
  XOR2_X1 U583 ( .A(KEYINPUT23), .B(n530), .Z(n531) );
  NAND2_X1 U584 ( .A1(n532), .A2(n531), .ZN(n538) );
  NOR2_X1 U585 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  XOR2_X2 U586 ( .A(KEYINPUT17), .B(n533), .Z(n881) );
  NAND2_X1 U587 ( .A1(G137), .A2(n881), .ZN(n536) );
  NOR2_X1 U588 ( .A1(G2104), .A2(n534), .ZN(n887) );
  NAND2_X1 U589 ( .A1(G125), .A2(n887), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X2 U591 ( .A1(n538), .A2(n537), .ZN(G160) );
  XOR2_X1 U592 ( .A(G2446), .B(KEYINPUT104), .Z(n540) );
  XNOR2_X1 U593 ( .A(G2451), .B(G2430), .ZN(n539) );
  XNOR2_X1 U594 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U595 ( .A(n541), .B(G2427), .Z(n543) );
  XNOR2_X1 U596 ( .A(G1348), .B(G1341), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n543), .B(n542), .ZN(n547) );
  XOR2_X1 U598 ( .A(G2443), .B(G2435), .Z(n545) );
  XNOR2_X1 U599 ( .A(G2438), .B(G2454), .ZN(n544) );
  XNOR2_X1 U600 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U601 ( .A(n547), .B(n546), .Z(n548) );
  AND2_X1 U602 ( .A1(G14), .A2(n548), .ZN(G401) );
  AND2_X1 U603 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U604 ( .A(G57), .ZN(G237) );
  NAND2_X1 U605 ( .A1(G90), .A2(n649), .ZN(n550) );
  XOR2_X1 U606 ( .A(KEYINPUT0), .B(G543), .Z(n636) );
  INV_X1 U607 ( .A(G651), .ZN(n553) );
  NOR2_X1 U608 ( .A1(n636), .A2(n553), .ZN(n653) );
  NAND2_X1 U609 ( .A1(G77), .A2(n653), .ZN(n549) );
  NAND2_X1 U610 ( .A1(n550), .A2(n549), .ZN(n552) );
  XOR2_X1 U611 ( .A(KEYINPUT9), .B(KEYINPUT69), .Z(n551) );
  XNOR2_X1 U612 ( .A(n552), .B(n551), .ZN(n558) );
  NOR2_X1 U613 ( .A1(G543), .A2(n553), .ZN(n554) );
  NAND2_X1 U614 ( .A1(G64), .A2(n650), .ZN(n556) );
  NAND2_X1 U615 ( .A1(G52), .A2(n647), .ZN(n555) );
  AND2_X1 U616 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(G301) );
  NAND2_X1 U618 ( .A1(n649), .A2(G89), .ZN(n559) );
  XNOR2_X1 U619 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G76), .A2(n653), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U622 ( .A(n562), .B(KEYINPUT5), .ZN(n568) );
  NAND2_X1 U623 ( .A1(n650), .A2(G63), .ZN(n563) );
  XNOR2_X1 U624 ( .A(n563), .B(KEYINPUT74), .ZN(n565) );
  NAND2_X1 U625 ( .A1(G51), .A2(n647), .ZN(n564) );
  NAND2_X1 U626 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U627 ( .A(KEYINPUT6), .B(n566), .Z(n567) );
  NAND2_X1 U628 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U629 ( .A(n569), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U632 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U633 ( .A(KEYINPUT70), .B(KEYINPUT11), .Z(n572) );
  INV_X1 U634 ( .A(G223), .ZN(n838) );
  NAND2_X1 U635 ( .A1(G567), .A2(n838), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n572), .B(n571), .ZN(G234) );
  NAND2_X1 U637 ( .A1(G56), .A2(n650), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT14), .B(n573), .Z(n579) );
  NAND2_X1 U639 ( .A1(n649), .A2(G81), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(KEYINPUT12), .ZN(n576) );
  NAND2_X1 U641 ( .A1(G68), .A2(n653), .ZN(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U643 ( .A(KEYINPUT13), .B(n577), .Z(n578) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U645 ( .A1(n647), .A2(G43), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n986) );
  INV_X1 U647 ( .A(G860), .ZN(n603) );
  OR2_X1 U648 ( .A1(n986), .A2(n603), .ZN(G153) );
  NAND2_X1 U649 ( .A1(G54), .A2(n647), .ZN(n588) );
  NAND2_X1 U650 ( .A1(G92), .A2(n649), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G79), .A2(n653), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U653 ( .A1(G66), .A2(n650), .ZN(n584) );
  XNOR2_X1 U654 ( .A(KEYINPUT71), .B(n584), .ZN(n585) );
  NOR2_X1 U655 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U657 ( .A(n589), .B(KEYINPUT15), .ZN(n590) );
  NOR2_X1 U658 ( .A1(G868), .A2(n711), .ZN(n591) );
  XNOR2_X1 U659 ( .A(n591), .B(KEYINPUT73), .ZN(n593) );
  NAND2_X1 U660 ( .A1(G868), .A2(G301), .ZN(n592) );
  NAND2_X1 U661 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U662 ( .A1(G91), .A2(n649), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G65), .A2(n650), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U665 ( .A1(G78), .A2(n653), .ZN(n597) );
  NAND2_X1 U666 ( .A1(G53), .A2(n647), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U668 ( .A1(n599), .A2(n598), .ZN(n701) );
  INV_X1 U669 ( .A(G868), .ZN(n659) );
  NAND2_X1 U670 ( .A1(n701), .A2(n659), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT75), .ZN(n602) );
  NOR2_X1 U672 ( .A1(n659), .A2(G286), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(G297) );
  INV_X1 U674 ( .A(n701), .ZN(G299) );
  NAND2_X1 U675 ( .A1(n603), .A2(G559), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n604), .A2(n711), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U678 ( .A1(G868), .A2(n986), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n711), .A2(G868), .ZN(n606) );
  NOR2_X1 U680 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U682 ( .A(KEYINPUT76), .B(n609), .ZN(G282) );
  NAND2_X1 U683 ( .A1(G135), .A2(n881), .ZN(n611) );
  NAND2_X1 U684 ( .A1(G111), .A2(n886), .ZN(n610) );
  NAND2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n887), .A2(G123), .ZN(n612) );
  XOR2_X1 U687 ( .A(KEYINPUT18), .B(n612), .Z(n613) );
  NOR2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n882), .A2(G99), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n948) );
  XNOR2_X1 U691 ( .A(G2096), .B(n948), .ZN(n617) );
  NOR2_X1 U692 ( .A1(n617), .A2(G2100), .ZN(n618) );
  XNOR2_X1 U693 ( .A(n618), .B(KEYINPUT77), .ZN(G156) );
  NAND2_X1 U694 ( .A1(n711), .A2(G559), .ZN(n619) );
  XNOR2_X1 U695 ( .A(n619), .B(n986), .ZN(n667) );
  NOR2_X1 U696 ( .A1(n667), .A2(G860), .ZN(n626) );
  NAND2_X1 U697 ( .A1(G67), .A2(n650), .ZN(n621) );
  NAND2_X1 U698 ( .A1(G55), .A2(n647), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G93), .A2(n649), .ZN(n623) );
  NAND2_X1 U701 ( .A1(G80), .A2(n653), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n664) );
  XNOR2_X1 U704 ( .A(n626), .B(n664), .ZN(G145) );
  NAND2_X1 U705 ( .A1(G88), .A2(n649), .ZN(n628) );
  NAND2_X1 U706 ( .A1(G75), .A2(n653), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n632) );
  NAND2_X1 U708 ( .A1(G62), .A2(n650), .ZN(n630) );
  NAND2_X1 U709 ( .A1(G50), .A2(n647), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U711 ( .A1(n632), .A2(n631), .ZN(G166) );
  NAND2_X1 U712 ( .A1(G49), .A2(n647), .ZN(n634) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U715 ( .A1(n650), .A2(n635), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n636), .A2(G87), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(G288) );
  NAND2_X1 U718 ( .A1(n647), .A2(G47), .ZN(n639) );
  XOR2_X1 U719 ( .A(KEYINPUT67), .B(n639), .Z(n641) );
  NAND2_X1 U720 ( .A1(n650), .A2(G60), .ZN(n640) );
  NAND2_X1 U721 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U722 ( .A(KEYINPUT68), .B(n642), .Z(n646) );
  NAND2_X1 U723 ( .A1(G85), .A2(n649), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G72), .A2(n653), .ZN(n643) );
  AND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(G290) );
  NAND2_X1 U727 ( .A1(G48), .A2(n647), .ZN(n648) );
  XNOR2_X1 U728 ( .A(n648), .B(KEYINPUT78), .ZN(n658) );
  NAND2_X1 U729 ( .A1(G86), .A2(n649), .ZN(n652) );
  NAND2_X1 U730 ( .A1(G61), .A2(n650), .ZN(n651) );
  NAND2_X1 U731 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U732 ( .A1(n653), .A2(G73), .ZN(n654) );
  XOR2_X1 U733 ( .A(KEYINPUT2), .B(n654), .Z(n655) );
  NOR2_X1 U734 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n658), .A2(n657), .ZN(G305) );
  NAND2_X1 U736 ( .A1(n659), .A2(n664), .ZN(n671) );
  XNOR2_X1 U737 ( .A(G166), .B(KEYINPUT79), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n660), .B(KEYINPUT19), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n701), .B(G288), .ZN(n661) );
  XNOR2_X1 U740 ( .A(n661), .B(G290), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n663), .B(n662), .ZN(n666) );
  XNOR2_X1 U742 ( .A(G305), .B(n664), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n666), .B(n665), .ZN(n908) );
  XNOR2_X1 U744 ( .A(n667), .B(n908), .ZN(n668) );
  XNOR2_X1 U745 ( .A(n668), .B(KEYINPUT80), .ZN(n669) );
  NAND2_X1 U746 ( .A1(n669), .A2(G868), .ZN(n670) );
  NAND2_X1 U747 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U748 ( .A(n672), .B(KEYINPUT81), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2084), .A2(G2078), .ZN(n673) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n673), .Z(n674) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U753 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U755 ( .A1(G132), .A2(G82), .ZN(n677) );
  XNOR2_X1 U756 ( .A(n677), .B(KEYINPUT82), .ZN(n678) );
  XNOR2_X1 U757 ( .A(n678), .B(KEYINPUT22), .ZN(n679) );
  NOR2_X1 U758 ( .A1(G218), .A2(n679), .ZN(n680) );
  NAND2_X1 U759 ( .A1(G96), .A2(n680), .ZN(n842) );
  NAND2_X1 U760 ( .A1(G2106), .A2(n842), .ZN(n684) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n681) );
  NOR2_X1 U762 ( .A1(G237), .A2(n681), .ZN(n682) );
  NAND2_X1 U763 ( .A1(G108), .A2(n682), .ZN(n843) );
  NAND2_X1 U764 ( .A1(G567), .A2(n843), .ZN(n683) );
  NAND2_X1 U765 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U766 ( .A(KEYINPUT83), .B(n685), .ZN(G319) );
  INV_X1 U767 ( .A(G319), .ZN(n914) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n686) );
  NOR2_X1 U769 ( .A1(n914), .A2(n686), .ZN(n841) );
  NAND2_X1 U770 ( .A1(n841), .A2(G36), .ZN(G176) );
  NAND2_X1 U771 ( .A1(G138), .A2(n881), .ZN(n688) );
  NAND2_X1 U772 ( .A1(G102), .A2(n882), .ZN(n687) );
  NAND2_X1 U773 ( .A1(n688), .A2(n687), .ZN(n692) );
  NAND2_X1 U774 ( .A1(G114), .A2(n886), .ZN(n690) );
  NAND2_X1 U775 ( .A1(G126), .A2(n887), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U777 ( .A1(n692), .A2(n691), .ZN(G164) );
  INV_X1 U778 ( .A(G166), .ZN(G303) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n800) );
  XNOR2_X1 U780 ( .A(n800), .B(KEYINPUT89), .ZN(n693) );
  NOR2_X1 U781 ( .A1(G164), .A2(G1384), .ZN(n799) );
  XNOR2_X1 U782 ( .A(KEYINPUT90), .B(n694), .ZN(n728) );
  NAND2_X1 U783 ( .A1(n728), .A2(G8), .ZN(n745) );
  NAND2_X1 U784 ( .A1(G8), .A2(n747), .ZN(n783) );
  NOR2_X1 U785 ( .A1(G1966), .A2(n783), .ZN(n729) );
  INV_X1 U786 ( .A(KEYINPUT93), .ZN(n695) );
  INV_X1 U787 ( .A(G2072), .ZN(n965) );
  NOR2_X1 U788 ( .A1(n723), .A2(n965), .ZN(n697) );
  XNOR2_X1 U789 ( .A(KEYINPUT94), .B(KEYINPUT27), .ZN(n696) );
  XNOR2_X1 U790 ( .A(n697), .B(n696), .ZN(n699) );
  NAND2_X1 U791 ( .A1(n723), .A2(G1956), .ZN(n698) );
  AND2_X1 U792 ( .A1(n699), .A2(n698), .ZN(n702) );
  XOR2_X1 U793 ( .A(n700), .B(KEYINPUT28), .Z(n720) );
  NAND2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n718) );
  XNOR2_X1 U795 ( .A(G1996), .B(KEYINPUT95), .ZN(n934) );
  XOR2_X1 U796 ( .A(n703), .B(KEYINPUT26), .Z(n705) );
  NAND2_X1 U797 ( .A1(n747), .A2(G1341), .ZN(n704) );
  NAND2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U799 ( .A(KEYINPUT64), .B(n707), .Z(n713) );
  NAND2_X1 U800 ( .A1(n747), .A2(G1348), .ZN(n710) );
  INV_X1 U801 ( .A(n723), .ZN(n708) );
  NAND2_X1 U802 ( .A1(G2067), .A2(n708), .ZN(n709) );
  NAND2_X1 U803 ( .A1(n710), .A2(n709), .ZN(n714) );
  INV_X1 U804 ( .A(n711), .ZN(n977) );
  AND2_X1 U805 ( .A1(n714), .A2(n977), .ZN(n712) );
  NOR2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n716) );
  NOR2_X1 U807 ( .A1(n977), .A2(n714), .ZN(n715) );
  NOR2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U810 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U811 ( .A(n721), .B(KEYINPUT29), .ZN(n727) );
  XNOR2_X1 U812 ( .A(G1961), .B(KEYINPUT91), .ZN(n1001) );
  NAND2_X1 U813 ( .A1(n747), .A2(n1001), .ZN(n722) );
  XOR2_X1 U814 ( .A(KEYINPUT92), .B(n722), .Z(n725) );
  XOR2_X1 U815 ( .A(G2078), .B(KEYINPUT25), .Z(n929) );
  NOR2_X1 U816 ( .A1(n929), .A2(n723), .ZN(n724) );
  NOR2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n734) );
  NOR2_X1 U818 ( .A1(G301), .A2(n734), .ZN(n726) );
  NOR2_X1 U819 ( .A1(n727), .A2(n726), .ZN(n741) );
  NOR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U821 ( .A(n730), .B(KEYINPUT96), .ZN(n731) );
  NAND2_X1 U822 ( .A1(n731), .A2(G8), .ZN(n732) );
  XNOR2_X1 U823 ( .A(n732), .B(KEYINPUT30), .ZN(n733) );
  NOR2_X1 U824 ( .A1(n733), .A2(G168), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n734), .A2(G301), .ZN(n735) );
  XNOR2_X1 U826 ( .A(n735), .B(KEYINPUT97), .ZN(n736) );
  NOR2_X1 U827 ( .A1(n737), .A2(n736), .ZN(n739) );
  NOR2_X1 U828 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U829 ( .A(n742), .B(KEYINPUT99), .ZN(n746) );
  INV_X1 U830 ( .A(n746), .ZN(n743) );
  NOR2_X1 U831 ( .A1(n729), .A2(n743), .ZN(n744) );
  NAND2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n757) );
  NAND2_X1 U833 ( .A1(n746), .A2(G286), .ZN(n754) );
  INV_X1 U834 ( .A(G8), .ZN(n752) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n747), .ZN(n749) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n783), .ZN(n748) );
  NOR2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n750), .A2(G303), .ZN(n751) );
  OR2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n753) );
  AND2_X1 U840 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U841 ( .A(n755), .B(KEYINPUT32), .ZN(n756) );
  NAND2_X1 U842 ( .A1(n757), .A2(n756), .ZN(n775) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n758) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n987) );
  NOR2_X1 U845 ( .A1(n758), .A2(n987), .ZN(n760) );
  INV_X1 U846 ( .A(KEYINPUT33), .ZN(n759) );
  AND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n775), .A2(n761), .ZN(n764) );
  INV_X1 U849 ( .A(KEYINPUT100), .ZN(n765) );
  NAND2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n989) );
  AND2_X1 U851 ( .A1(n527), .A2(n989), .ZN(n762) );
  OR2_X1 U852 ( .A1(KEYINPUT33), .A2(n762), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n771) );
  NAND2_X1 U854 ( .A1(n765), .A2(n987), .ZN(n768) );
  NAND2_X1 U855 ( .A1(n987), .A2(KEYINPUT33), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n766), .A2(KEYINPUT100), .ZN(n767) );
  NAND2_X1 U857 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U858 ( .A1(n783), .A2(n769), .ZN(n770) );
  NOR2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U860 ( .A(G1981), .B(G305), .Z(n982) );
  NAND2_X1 U861 ( .A1(n772), .A2(n982), .ZN(n780) );
  NOR2_X1 U862 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U863 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n777) );
  XNOR2_X1 U865 ( .A(n777), .B(n776), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n778), .A2(n783), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n785) );
  NOR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n781) );
  XOR2_X1 U869 ( .A(n781), .B(KEYINPUT24), .Z(n782) );
  NOR2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n786) );
  INV_X1 U872 ( .A(n786), .ZN(n821) );
  XNOR2_X1 U873 ( .A(G2067), .B(KEYINPUT37), .ZN(n831) );
  NAND2_X1 U874 ( .A1(n882), .A2(G104), .ZN(n787) );
  XOR2_X1 U875 ( .A(KEYINPUT85), .B(n787), .Z(n789) );
  NAND2_X1 U876 ( .A1(n881), .A2(G140), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U878 ( .A(KEYINPUT34), .B(n790), .ZN(n796) );
  NAND2_X1 U879 ( .A1(G116), .A2(n886), .ZN(n792) );
  NAND2_X1 U880 ( .A1(G128), .A2(n887), .ZN(n791) );
  NAND2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U882 ( .A(KEYINPUT35), .B(n793), .Z(n794) );
  XNOR2_X1 U883 ( .A(KEYINPUT86), .B(n794), .ZN(n795) );
  NOR2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U885 ( .A(n797), .B(KEYINPUT36), .Z(n798) );
  XNOR2_X1 U886 ( .A(KEYINPUT87), .B(n798), .ZN(n905) );
  NOR2_X1 U887 ( .A1(n831), .A2(n905), .ZN(n954) );
  NOR2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U889 ( .A(n801), .B(KEYINPUT84), .ZN(n833) );
  NAND2_X1 U890 ( .A1(n954), .A2(n833), .ZN(n829) );
  INV_X1 U891 ( .A(n829), .ZN(n819) );
  NAND2_X1 U892 ( .A1(G141), .A2(n881), .ZN(n803) );
  NAND2_X1 U893 ( .A1(G117), .A2(n886), .ZN(n802) );
  NAND2_X1 U894 ( .A1(n803), .A2(n802), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n882), .A2(G105), .ZN(n804) );
  XOR2_X1 U896 ( .A(KEYINPUT38), .B(n804), .Z(n805) );
  NOR2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n808) );
  NAND2_X1 U898 ( .A1(n887), .A2(G129), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n808), .A2(n807), .ZN(n880) );
  NAND2_X1 U900 ( .A1(n880), .A2(G1996), .ZN(n817) );
  NAND2_X1 U901 ( .A1(G95), .A2(n882), .ZN(n810) );
  NAND2_X1 U902 ( .A1(G119), .A2(n887), .ZN(n809) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n813) );
  NAND2_X1 U904 ( .A1(n886), .A2(G107), .ZN(n811) );
  XOR2_X1 U905 ( .A(KEYINPUT88), .B(n811), .Z(n812) );
  NOR2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n815) );
  NAND2_X1 U907 ( .A1(n881), .A2(G131), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n897) );
  NAND2_X1 U909 ( .A1(G1991), .A2(n897), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n824) );
  INV_X1 U911 ( .A(n824), .ZN(n951) );
  XOR2_X1 U912 ( .A(G1986), .B(G290), .Z(n998) );
  NAND2_X1 U913 ( .A1(n951), .A2(n998), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n836) );
  XOR2_X1 U915 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n828) );
  NOR2_X1 U916 ( .A1(G1996), .A2(n880), .ZN(n959) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n822) );
  NOR2_X1 U918 ( .A1(G1991), .A2(n897), .ZN(n947) );
  NOR2_X1 U919 ( .A1(n822), .A2(n947), .ZN(n823) );
  NOR2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n825), .B(KEYINPUT102), .ZN(n826) );
  NOR2_X1 U922 ( .A1(n959), .A2(n826), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n828), .B(n827), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(n832) );
  NAND2_X1 U925 ( .A1(n831), .A2(n905), .ZN(n956) );
  NAND2_X1 U926 ( .A1(n832), .A2(n956), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U929 ( .A(KEYINPUT40), .B(n837), .ZN(G329) );
  INV_X1 U930 ( .A(G301), .ZN(G171) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n838), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U933 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(G188) );
  INV_X1 U937 ( .A(G132), .ZN(G219) );
  INV_X1 U938 ( .A(G120), .ZN(G236) );
  INV_X1 U939 ( .A(G82), .ZN(G220) );
  INV_X1 U940 ( .A(G69), .ZN(G235) );
  NOR2_X1 U941 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  XOR2_X1 U943 ( .A(G2100), .B(G2096), .Z(n845) );
  XNOR2_X1 U944 ( .A(KEYINPUT42), .B(G2678), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U946 ( .A(KEYINPUT43), .B(G2090), .Z(n847) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2072), .ZN(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U949 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U950 ( .A(G2084), .B(G2078), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(G227) );
  XOR2_X1 U952 ( .A(KEYINPUT41), .B(G1976), .Z(n853) );
  XNOR2_X1 U953 ( .A(G1956), .B(G1971), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U955 ( .A(n854), .B(KEYINPUT106), .Z(n856) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U958 ( .A(G1986), .B(G1981), .Z(n858) );
  XNOR2_X1 U959 ( .A(G1966), .B(G1961), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U961 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U962 ( .A(KEYINPUT105), .B(G2474), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U964 ( .A1(G124), .A2(n887), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n886), .A2(G112), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G136), .A2(n881), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G100), .A2(n882), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U971 ( .A1(n869), .A2(n868), .ZN(G162) );
  NAND2_X1 U972 ( .A1(n886), .A2(G115), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n870), .B(KEYINPUT110), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G127), .A2(n887), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U976 ( .A(n873), .B(KEYINPUT47), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G103), .A2(n882), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G139), .A2(n881), .ZN(n876) );
  XNOR2_X1 U980 ( .A(KEYINPUT109), .B(n876), .ZN(n877) );
  NOR2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U982 ( .A(KEYINPUT111), .B(n879), .Z(n964) );
  XNOR2_X1 U983 ( .A(n964), .B(n880), .ZN(n895) );
  NAND2_X1 U984 ( .A1(G142), .A2(n881), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G106), .A2(n882), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U987 ( .A(n885), .B(KEYINPUT45), .ZN(n892) );
  NAND2_X1 U988 ( .A1(G118), .A2(n886), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G130), .A2(n887), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U991 ( .A(KEYINPUT107), .B(n890), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n893), .B(n948), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n899) );
  XOR2_X1 U995 ( .A(G160), .B(G162), .Z(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U997 ( .A(n899), .B(n898), .Z(n904) );
  XOR2_X1 U998 ( .A(KEYINPUT108), .B(KEYINPUT48), .Z(n901) );
  XNOR2_X1 U999 ( .A(KEYINPUT112), .B(KEYINPUT46), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(G164), .B(n902), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1003 ( .A(n906), .B(n905), .Z(n907) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n907), .ZN(G395) );
  XOR2_X1 U1005 ( .A(KEYINPUT113), .B(n908), .Z(n910) );
  XNOR2_X1 U1006 ( .A(G171), .B(G286), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n912) );
  XOR2_X1 U1008 ( .A(n986), .B(n977), .Z(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n913), .ZN(G397) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n914), .ZN(n915) );
  XOR2_X1 U1012 ( .A(KEYINPUT114), .B(n915), .Z(n919) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n916) );
  XOR2_X1 U1014 ( .A(KEYINPUT115), .B(n916), .Z(n917) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(KEYINPUT116), .B(n920), .ZN(n922) );
  NOR2_X1 U1018 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1020 ( .A(G225), .ZN(G308) );
  INV_X1 U1021 ( .A(G108), .ZN(G238) );
  INV_X1 U1022 ( .A(G96), .ZN(G221) );
  XNOR2_X1 U1023 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(n923), .B(G34), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(G2084), .B(n924), .ZN(n942) );
  XNOR2_X1 U1026 ( .A(G2090), .B(G35), .ZN(n925) );
  XNOR2_X1 U1027 ( .A(n925), .B(KEYINPUT120), .ZN(n939) );
  XNOR2_X1 U1028 ( .A(G2067), .B(G26), .ZN(n927) );
  XNOR2_X1 U1029 ( .A(G1991), .B(G25), .ZN(n926) );
  NOR2_X1 U1030 ( .A1(n927), .A2(n926), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(G33), .B(n965), .ZN(n928) );
  NAND2_X1 U1032 ( .A1(n928), .A2(G28), .ZN(n931) );
  XNOR2_X1 U1033 ( .A(G27), .B(n929), .ZN(n930) );
  NOR2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n936) );
  XOR2_X1 U1036 ( .A(G32), .B(n934), .Z(n935) );
  NOR2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(n937), .B(KEYINPUT53), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT121), .B(n940), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1042 ( .A(KEYINPUT123), .B(n943), .Z(n944) );
  NOR2_X1 U1043 ( .A1(G29), .A2(n944), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(n945), .B(KEYINPUT55), .ZN(n974) );
  XOR2_X1 U1045 ( .A(G2084), .B(G160), .Z(n946) );
  NOR2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n949) );
  NAND2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(KEYINPUT117), .B(n950), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(n955), .B(KEYINPUT118), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n962) );
  XOR2_X1 U1053 ( .A(G2090), .B(G162), .Z(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n960), .B(KEYINPUT51), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1057 ( .A(KEYINPUT119), .B(n963), .Z(n970) );
  XOR2_X1 U1058 ( .A(G164), .B(G2078), .Z(n967) );
  XNOR2_X1 U1059 ( .A(n965), .B(n964), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT50), .B(n968), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(KEYINPUT52), .B(n971), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(G29), .A2(n972), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n974), .A2(n973), .ZN(n1029) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n1000) );
  XNOR2_X1 U1067 ( .A(G299), .B(G1956), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(G303), .B(G1971), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G301), .B(G1961), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n977), .B(G1348), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n996) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G168), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(n984), .B(KEYINPUT57), .ZN(n994) );
  XOR2_X1 U1077 ( .A(G1341), .B(KEYINPUT125), .Z(n985) );
  XNOR2_X1 U1078 ( .A(n986), .B(n985), .ZN(n992) );
  INV_X1 U1079 ( .A(n987), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(KEYINPUT124), .B(n990), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1083 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1086 ( .A1(n1000), .A2(n999), .ZN(n1026) );
  INV_X1 U1087 ( .A(G16), .ZN(n1024) );
  XNOR2_X1 U1088 ( .A(G5), .B(n1001), .ZN(n1021) );
  XOR2_X1 U1089 ( .A(G1966), .B(G21), .Z(n1012) );
  XOR2_X1 U1090 ( .A(G1956), .B(G20), .Z(n1005) );
  XNOR2_X1 U1091 ( .A(G1341), .B(G19), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G1981), .B(G6), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(KEYINPUT126), .B(n1006), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(KEYINPUT59), .B(G1348), .Z(n1007) );
  XNOR2_X1 U1097 ( .A(G4), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(KEYINPUT60), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(G1986), .B(G24), .Z(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1022), .Z(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT127), .B(n1027), .Z(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(G11), .ZN(n1031) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

