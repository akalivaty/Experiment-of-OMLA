//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G952), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(G234), .A2(G237), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT21), .B(G898), .Z(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(G902), .A3(G953), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(G214), .B1(G237), .B2(G902), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G101), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G104), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(new_n197), .A3(G104), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n199), .A2(new_n197), .A3(KEYINPUT79), .A4(G104), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n198), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(new_n205), .B2(G107), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT78), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n197), .A2(G104), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n196), .B1(new_n204), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT4), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n202), .A2(new_n203), .ZN(new_n215));
  INV_X1    g029(.A(new_n198), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n211), .A2(new_n215), .A3(new_n196), .A4(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT80), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT80), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n204), .A2(new_n219), .A3(new_n196), .A4(new_n211), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n214), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n213), .B1(new_n221), .B2(new_n212), .ZN(new_n222));
  XOR2_X1   g036(.A(KEYINPUT2), .B(G113), .Z(new_n223));
  XNOR2_X1  g037(.A(G116), .B(G119), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n216), .A2(new_n209), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G101), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n224), .A2(KEYINPUT5), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT5), .ZN(new_n231));
  INV_X1    g045(.A(G119), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(G116), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n230), .A2(G113), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n223), .A2(new_n224), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI211_X1 g050(.A(new_n229), .B(new_n236), .C1(new_n218), .C2(new_n220), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n226), .A2(new_n238), .ZN(new_n239));
  XOR2_X1   g053(.A(G110), .B(G122), .Z(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n240), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n226), .A2(new_n238), .A3(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n241), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n242), .B1(new_n226), .B2(new_n238), .ZN(new_n245));
  AOI211_X1 g059(.A(new_n240), .B(new_n237), .C1(new_n222), .C2(new_n225), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT6), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n239), .A2(new_n247), .A3(new_n240), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT85), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n244), .B1(new_n248), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G143), .ZN(new_n255));
  INV_X1    g069(.A(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G146), .ZN(new_n257));
  AND4_X1   g071(.A1(new_n253), .A2(new_n255), .A3(new_n257), .A4(G128), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n255), .A2(new_n257), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n254), .A2(G143), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n260), .A2(new_n261), .B1(KEYINPUT1), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(KEYINPUT69), .ZN(new_n264));
  AOI21_X1  g078(.A(G128), .B1(new_n255), .B2(new_n257), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n257), .A2(new_n253), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n259), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G125), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n272));
  NAND2_X1  g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n272), .B1(new_n260), .B2(new_n273), .ZN(new_n274));
  OR2_X1    g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n260), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n274), .B(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G125), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n271), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G224), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(G953), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n280), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n252), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n286));
  OR3_X1    g100(.A1(new_n280), .A2(new_n286), .A3(new_n282), .ZN(new_n287));
  XOR2_X1   g101(.A(new_n240), .B(KEYINPUT8), .Z(new_n288));
  AOI21_X1  g102(.A(new_n229), .B1(new_n218), .B2(new_n220), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n289), .B1(new_n235), .B2(new_n234), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n288), .B1(new_n290), .B2(new_n237), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n280), .B1(new_n286), .B2(new_n282), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n287), .A2(new_n291), .A3(new_n292), .A4(new_n243), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n284), .A2(new_n285), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G210), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT86), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n284), .A2(new_n285), .A3(new_n297), .A4(new_n293), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n195), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G469), .ZN(new_n302));
  XOR2_X1   g116(.A(G110), .B(G140), .Z(new_n303));
  XNOR2_X1  g117(.A(new_n303), .B(KEYINPUT77), .ZN(new_n304));
  INV_X1    g118(.A(G227), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(G953), .ZN(new_n306));
  XOR2_X1   g120(.A(new_n304), .B(new_n306), .Z(new_n307));
  INV_X1    g121(.A(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n218), .A2(new_n220), .ZN(new_n309));
  XNOR2_X1  g123(.A(G143), .B(G146), .ZN(new_n310));
  OAI22_X1  g124(.A1(new_n310), .A2(G128), .B1(new_n253), .B2(new_n257), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n228), .B1(new_n311), .B2(new_n258), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT81), .B1(new_n309), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n315));
  AOI211_X1 g129(.A(new_n315), .B(new_n312), .C1(new_n218), .C2(new_n220), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n308), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT82), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n277), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n270), .A2(new_n308), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n222), .A2(new_n320), .B1(new_n289), .B2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(KEYINPUT82), .B(new_n308), .C1(new_n314), .C2(new_n316), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n319), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G131), .ZN(new_n325));
  OR2_X1    g139(.A1(KEYINPUT65), .A2(G134), .ZN(new_n326));
  INV_X1    g140(.A(G137), .ZN(new_n327));
  NAND2_X1  g141(.A1(KEYINPUT65), .A2(G134), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT11), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n329), .A2(KEYINPUT66), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT66), .B1(new_n329), .B2(new_n330), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(KEYINPUT67), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT67), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G137), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n330), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n326), .A2(new_n328), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n337), .A2(G134), .B1(new_n338), .B2(G137), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n325), .B1(new_n333), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT66), .ZN(new_n341));
  AND2_X1   g155(.A1(KEYINPUT65), .A2(G134), .ZN(new_n342));
  NOR2_X1   g156(.A1(KEYINPUT65), .A2(G134), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n342), .A2(new_n343), .A3(G137), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n341), .B1(new_n344), .B2(KEYINPUT11), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n329), .A2(KEYINPUT66), .A3(new_n330), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n339), .A2(new_n345), .A3(new_n325), .A4(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n340), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n324), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT83), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n324), .A2(KEYINPUT83), .A3(new_n350), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n319), .A2(new_n349), .A3(new_n322), .A4(new_n323), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n307), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n356), .A2(KEYINPUT84), .A3(new_n307), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT12), .ZN(new_n359));
  OAI22_X1  g173(.A1(new_n314), .A2(new_n316), .B1(new_n289), .B2(new_n269), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n359), .B1(new_n361), .B2(new_n349), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n360), .A2(KEYINPUT12), .A3(new_n350), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT84), .B1(new_n356), .B2(new_n307), .ZN(new_n366));
  NOR3_X1   g180(.A1(new_n358), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n302), .B(new_n285), .C1(new_n357), .C2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n302), .A2(new_n285), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n307), .B1(new_n364), .B2(new_n356), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n356), .A2(new_n307), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n370), .B1(new_n355), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n369), .B1(new_n373), .B2(G469), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT9), .B(G234), .Z(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(G221), .B1(new_n377), .B2(G902), .ZN(new_n378));
  XNOR2_X1  g192(.A(G125), .B(G140), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(new_n254), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT87), .ZN(new_n381));
  NOR2_X1   g195(.A1(G237), .A2(G953), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(G143), .A3(G214), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(G143), .B1(new_n382), .B2(G214), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n381), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(KEYINPUT18), .A2(G131), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G237), .ZN(new_n389));
  INV_X1    g203(.A(G953), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(G214), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n256), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(KEYINPUT87), .A3(new_n383), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n386), .A2(new_n388), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT88), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n384), .A2(new_n385), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n395), .B1(new_n396), .B2(new_n387), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n392), .A2(new_n383), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n398), .A2(KEYINPUT88), .A3(new_n388), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n380), .B(new_n394), .C1(new_n397), .C2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G131), .B1(new_n384), .B2(new_n385), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT17), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n392), .A2(new_n325), .A3(new_n383), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n379), .A2(KEYINPUT16), .ZN(new_n405));
  OR3_X1    g219(.A1(new_n278), .A2(KEYINPUT16), .A3(G140), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n254), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n398), .A2(KEYINPUT17), .A3(G131), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(G146), .A3(new_n406), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n404), .A2(new_n408), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G113), .B(G122), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n412), .B(new_n205), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n400), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT89), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n400), .A2(new_n411), .A3(KEYINPUT89), .A4(new_n413), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n400), .A2(new_n411), .ZN(new_n419));
  INV_X1    g233(.A(new_n413), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT90), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n285), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n416), .A2(new_n417), .B1(new_n420), .B2(new_n419), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT90), .B1(new_n425), .B2(G902), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n426), .A3(G475), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n401), .A2(new_n403), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n379), .B(KEYINPUT19), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n254), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n410), .A2(KEYINPUT74), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n410), .A2(KEYINPUT74), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n429), .B(new_n431), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n400), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n416), .A2(new_n417), .B1(new_n420), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(G475), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n428), .B1(new_n437), .B2(new_n285), .ZN(new_n438));
  NOR4_X1   g252(.A1(new_n436), .A2(KEYINPUT20), .A3(G475), .A4(G902), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n427), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n261), .A2(G143), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT91), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n256), .A2(G128), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT13), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n256), .A2(KEYINPUT13), .A3(G128), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G134), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n444), .A2(new_n338), .A3(new_n445), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(G116), .B(G122), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(new_n197), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n444), .A2(KEYINPUT92), .A3(new_n338), .A4(new_n445), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n450), .A2(new_n453), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT14), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G122), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n460), .A2(G116), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n197), .B1(new_n461), .B2(KEYINPUT14), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n459), .A2(new_n462), .B1(new_n197), .B2(new_n454), .ZN(new_n463));
  INV_X1    g277(.A(new_n451), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n338), .B1(new_n444), .B2(new_n445), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n457), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G217), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n377), .A2(new_n468), .A3(G953), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n457), .A2(new_n466), .A3(new_n469), .ZN(new_n472));
  AOI21_X1  g286(.A(G902), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G478), .ZN(new_n474));
  OR3_X1    g288(.A1(new_n473), .A2(KEYINPUT15), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n473), .B1(KEYINPUT15), .B2(new_n474), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n441), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n301), .A2(new_n375), .A3(new_n378), .A4(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT93), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n468), .B1(G234), .B2(new_n285), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT23), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n232), .B2(G128), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n232), .A2(G128), .ZN(new_n488));
  MUX2_X1   g302(.A(new_n487), .B(new_n486), .S(new_n488), .Z(new_n489));
  INV_X1    g303(.A(G110), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  XOR2_X1   g305(.A(G119), .B(G128), .Z(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT24), .B(G110), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n491), .A2(new_n494), .B1(new_n254), .B2(new_n379), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n495), .B1(new_n432), .B2(new_n433), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n408), .A2(new_n410), .ZN(new_n497));
  OAI221_X1 g311(.A(new_n497), .B1(new_n490), .B2(new_n489), .C1(new_n492), .C2(new_n493), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n390), .A2(G221), .A3(G234), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(G137), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT75), .B(KEYINPUT22), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n501), .B(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n499), .B(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(G902), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n505), .A2(KEYINPUT25), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(KEYINPUT25), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n485), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n485), .A2(new_n285), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT76), .ZN(new_n510));
  INV_X1    g324(.A(new_n504), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G472), .ZN(new_n514));
  INV_X1    g328(.A(G134), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n334), .A2(new_n336), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n325), .B1(new_n329), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT68), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n518), .A2(new_n269), .A3(new_n347), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n339), .A2(new_n345), .A3(new_n346), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(G131), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n277), .B1(new_n521), .B2(new_n347), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n519), .A2(new_n522), .A3(KEYINPUT30), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n320), .B1(new_n340), .B2(new_n348), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n518), .A2(new_n269), .A3(new_n347), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n225), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT70), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n382), .A2(G210), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(new_n196), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n532));
  XOR2_X1   g346(.A(new_n531), .B(new_n532), .Z(new_n533));
  XNOR2_X1  g347(.A(new_n225), .B(KEYINPUT71), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n535), .A2(new_n525), .A3(new_n526), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT30), .B1(new_n519), .B2(new_n522), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n525), .A2(new_n524), .A3(new_n526), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT70), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n540), .A3(new_n225), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n529), .A2(new_n533), .A3(new_n536), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT31), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n519), .A2(new_n522), .A3(new_n534), .ZN(new_n545));
  INV_X1    g359(.A(new_n225), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n525), .B2(new_n526), .ZN(new_n547));
  OAI21_X1  g361(.A(KEYINPUT28), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT72), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n545), .B2(KEYINPUT28), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT28), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n536), .A2(KEYINPUT72), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n548), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n533), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n542), .B2(KEYINPUT31), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n514), .B(new_n285), .C1(new_n544), .C2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT32), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT73), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT73), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n557), .A2(new_n561), .A3(new_n558), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n540), .B1(new_n539), .B2(new_n225), .ZN(new_n564));
  AOI211_X1 g378(.A(KEYINPUT70), .B(new_n546), .C1(new_n537), .C2(new_n538), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT31), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n533), .A4(new_n536), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(new_n543), .A3(new_n555), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n569), .A2(KEYINPUT32), .A3(new_n514), .A4(new_n285), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n533), .B1(new_n553), .B2(KEYINPUT29), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n534), .B1(new_n519), .B2(new_n522), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n536), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT28), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n550), .A3(new_n552), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n285), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n529), .A2(new_n554), .A3(new_n536), .A4(new_n541), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT29), .B1(new_n571), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(G472), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n570), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n513), .B1(new_n563), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n378), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n368), .B2(new_n374), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n583), .A2(KEYINPUT93), .A3(new_n301), .A4(new_n480), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n483), .A2(new_n581), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  XNOR2_X1  g400(.A(new_n294), .B(new_n296), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n193), .A3(new_n194), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT33), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n457), .A2(new_n466), .A3(new_n469), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n469), .B1(new_n457), .B2(new_n466), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n471), .A2(KEYINPUT33), .A3(new_n472), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n592), .A2(new_n593), .A3(new_n285), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT94), .B1(new_n473), .B2(G478), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n285), .B1(new_n590), .B2(new_n591), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT94), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n474), .ZN(new_n598));
  AOI22_X1  g412(.A1(G478), .A2(new_n594), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n435), .A2(new_n420), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n418), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(G475), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n601), .A2(new_n602), .A3(new_n285), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT20), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n437), .A2(new_n428), .A3(new_n285), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n599), .B1(new_n606), .B2(new_n427), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n588), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n569), .A2(new_n285), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(G472), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n557), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n375), .A2(new_n378), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n513), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n609), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  NOR3_X1   g432(.A1(new_n588), .A2(new_n478), .A3(new_n440), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n613), .A3(new_n615), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT35), .B(G107), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  INV_X1    g436(.A(new_n508), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n503), .A2(KEYINPUT36), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n499), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n510), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n483), .A2(new_n584), .A3(new_n613), .A4(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT37), .B(G110), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G12));
  AOI22_X1  g444(.A1(new_n563), .A2(new_n580), .B1(new_n623), .B2(new_n626), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n587), .A2(new_n194), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n614), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n190), .B1(G900), .B2(new_n192), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n441), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n478), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n631), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT95), .B(G128), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G30));
  XOR2_X1   g453(.A(new_n634), .B(KEYINPUT39), .Z(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n583), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(KEYINPUT40), .Z(new_n643));
  INV_X1    g457(.A(new_n194), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n440), .A2(new_n477), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n627), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT96), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n566), .A2(new_n536), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n533), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n285), .B1(new_n573), .B2(new_n533), .ZN(new_n651));
  OAI21_X1  g465(.A(G472), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n563), .A2(new_n570), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n299), .A2(new_n300), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT38), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n643), .A2(new_n647), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G143), .ZN(G45));
  INV_X1    g471(.A(KEYINPUT97), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n607), .B2(new_n634), .ZN(new_n659));
  INV_X1    g473(.A(new_n599), .ZN(new_n660));
  AND4_X1   g474(.A1(new_n658), .A2(new_n440), .A3(new_n660), .A4(new_n634), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n631), .A2(new_n633), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G146), .ZN(G48));
  NAND2_X1  g478(.A1(new_n368), .A2(KEYINPUT98), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n324), .A2(KEYINPUT83), .A3(new_n350), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT83), .B1(new_n324), .B2(new_n350), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n356), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n307), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n358), .A2(new_n366), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n364), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n302), .B1(new_n673), .B2(new_n285), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n665), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT98), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n668), .A2(new_n669), .B1(new_n671), .B2(new_n364), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n676), .B(G469), .C1(new_n677), .C2(G902), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n378), .B1(new_n675), .B2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT99), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(G469), .B1(new_n677), .B2(G902), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(KEYINPUT98), .A3(new_n368), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n678), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(KEYINPUT99), .A3(new_n378), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n682), .A2(new_n581), .A3(new_n609), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G15));
  NAND4_X1  g503(.A1(new_n682), .A2(new_n581), .A3(new_n619), .A4(new_n686), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G116), .ZN(G18));
  AOI21_X1  g505(.A(KEYINPUT99), .B1(new_n685), .B2(new_n378), .ZN(new_n692));
  AOI211_X1 g506(.A(new_n681), .B(new_n582), .C1(new_n684), .C2(new_n678), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n632), .ZN(new_n695));
  AND2_X1   g509(.A1(new_n631), .A2(new_n193), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n694), .A2(new_n480), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G119), .ZN(G21));
  INV_X1    g512(.A(new_n645), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n575), .A2(new_n554), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n568), .A2(new_n543), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n514), .A3(new_n285), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n611), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n512), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n588), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n682), .A2(new_n699), .A3(new_n686), .A4(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT100), .B(G122), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G24));
  AND4_X1   g522(.A1(new_n611), .A2(new_n662), .A3(new_n627), .A4(new_n702), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n682), .A2(new_n695), .A3(new_n686), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  OAI211_X1 g525(.A(new_n570), .B(new_n579), .C1(new_n559), .C2(KEYINPUT101), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n557), .B2(new_n558), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n512), .B(new_n662), .C1(new_n712), .C2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n299), .A2(new_n300), .A3(new_n194), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n583), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(KEYINPUT42), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n717), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n659), .A2(new_n661), .A3(KEYINPUT42), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n581), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G131), .ZN(G33));
  NAND3_X1  g537(.A1(new_n581), .A2(new_n719), .A3(new_n636), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G134), .ZN(G36));
  INV_X1    g539(.A(KEYINPUT103), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT43), .B1(new_n441), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n441), .A2(new_n660), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n612), .A3(new_n627), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n729), .A2(KEYINPUT44), .A3(new_n612), .A4(new_n627), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n716), .A3(new_n733), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n734), .A2(KEYINPUT104), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n373), .A2(KEYINPUT45), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n371), .B1(new_n353), .B2(new_n354), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n737), .B1(new_n738), .B2(new_n370), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(G469), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT102), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n736), .A2(KEYINPUT102), .A3(G469), .A4(new_n739), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n369), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(KEYINPUT46), .ZN(new_n745));
  INV_X1    g559(.A(new_n368), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(new_n744), .B2(KEYINPUT46), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n582), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n734), .A2(KEYINPUT104), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n735), .A2(new_n641), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G137), .ZN(G39));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n557), .A2(new_n561), .A3(new_n558), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n561), .B1(new_n557), .B2(new_n558), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n580), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n299), .A2(new_n300), .A3(new_n194), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n757), .A2(new_n512), .A3(new_n758), .ZN(new_n759));
  AOI211_X1 g573(.A(KEYINPUT47), .B(new_n582), .C1(new_n745), .C2(new_n747), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n754), .A2(new_n662), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT105), .B(G140), .Z(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G42));
  NOR2_X1   g578(.A1(new_n758), .A2(new_n190), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n694), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n653), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n512), .A3(new_n607), .A4(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n655), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n729), .A2(new_n189), .A3(new_n188), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n512), .A3(new_n703), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n694), .A2(new_n644), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(KEYINPUT50), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n441), .A2(new_n599), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n766), .A2(new_n512), .A3(new_n767), .A4(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n694), .A2(new_n729), .A3(new_n765), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n703), .A2(new_n627), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n773), .A2(KEYINPUT50), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n774), .A2(new_n777), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT113), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n685), .A2(new_n582), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n753), .B2(new_n760), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n771), .A2(new_n758), .ZN(new_n788));
  OAI211_X1 g602(.A(KEYINPUT114), .B(new_n784), .C1(new_n753), .C2(new_n760), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AND2_X1   g604(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n783), .B(new_n790), .C1(new_n782), .C2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n785), .A2(new_n788), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n793), .B1(new_n794), .B2(new_n782), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n512), .B1(new_n712), .B2(new_n714), .ZN(new_n796));
  INV_X1    g610(.A(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n778), .A2(new_n797), .B1(new_n798), .B2(KEYINPUT48), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n798), .B2(KEYINPUT48), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n778), .A2(new_n798), .A3(KEYINPUT48), .A4(new_n797), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n800), .A2(new_n188), .A3(new_n801), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n768), .A2(new_n792), .A3(new_n795), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n631), .B(new_n633), .C1(new_n636), .C2(new_n662), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n646), .A2(new_n587), .A3(new_n634), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n653), .A2(new_n806), .A3(new_n583), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n710), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n808), .A2(KEYINPUT112), .A3(KEYINPUT52), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT52), .B1(new_n808), .B2(KEYINPUT112), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n697), .A2(new_n687), .A3(new_n690), .A4(new_n706), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n477), .B(KEYINPUT109), .Z(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n441), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n615), .A2(new_n301), .A3(new_n613), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n628), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT108), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n607), .B(KEYINPUT107), .Z(new_n820));
  NAND4_X1  g634(.A1(new_n615), .A2(new_n301), .A3(new_n613), .A4(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n585), .A2(new_n819), .A3(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n819), .B1(new_n585), .B2(new_n821), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n818), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n757), .A2(new_n583), .A3(new_n627), .A4(new_n716), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n813), .A2(new_n635), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n825), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n631), .A2(new_n719), .A3(KEYINPUT110), .A4(new_n827), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n662), .A2(new_n611), .A3(new_n627), .A4(new_n702), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n832), .B1(new_n717), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n709), .A2(KEYINPUT111), .A3(new_n583), .A4(new_n716), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n722), .A2(new_n831), .A3(new_n724), .A4(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n812), .A2(new_n824), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n811), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n585), .A2(new_n821), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT108), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n585), .A2(new_n819), .A3(new_n821), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n817), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n687), .A2(new_n690), .A3(new_n706), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n829), .A2(new_n830), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n836), .A2(new_n718), .A3(new_n721), .A4(new_n724), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n845), .A2(new_n846), .A3(new_n849), .A4(new_n697), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n808), .A2(KEYINPUT52), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n710), .A2(new_n852), .A3(new_n805), .A4(new_n807), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n850), .A2(new_n854), .A3(new_n840), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n804), .B1(new_n841), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n811), .A2(KEYINPUT53), .A3(new_n838), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n840), .B1(new_n850), .B2(new_n854), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n858), .A2(new_n804), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n694), .A2(new_n695), .A3(new_n772), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n803), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n811), .B2(new_n838), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT54), .B1(new_n865), .B2(new_n855), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n858), .A2(new_n804), .A3(new_n859), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n863), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n792), .A2(new_n795), .A3(new_n768), .A4(new_n802), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT116), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n187), .A2(new_n390), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n864), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n685), .ZN(new_n873));
  AOI211_X1 g687(.A(new_n644), .B(new_n728), .C1(new_n873), .C2(KEYINPUT49), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n767), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n769), .B(new_n512), .C1(KEYINPUT49), .C2(new_n873), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n875), .A2(new_n876), .A3(new_n582), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT106), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n872), .A2(new_n878), .ZN(G75));
  AOI21_X1  g693(.A(new_n285), .B1(new_n858), .B2(new_n859), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT56), .B1(new_n880), .B2(G210), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n252), .B(new_n283), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT55), .Z(new_n883));
  AND2_X1   g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n881), .A2(new_n883), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n390), .A2(G952), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G51));
  NAND2_X1  g701(.A1(new_n742), .A2(new_n743), .ZN(new_n888));
  AOI211_X1 g702(.A(new_n285), .B(new_n888), .C1(new_n858), .C2(new_n859), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n369), .B(KEYINPUT57), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n804), .B1(new_n858), .B2(new_n859), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n890), .B1(new_n860), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n889), .B1(new_n892), .B2(new_n673), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT117), .B1(new_n893), .B2(new_n886), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n895));
  INV_X1    g709(.A(new_n886), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n858), .A2(new_n859), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n867), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n677), .B1(new_n899), .B2(new_n890), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n895), .B(new_n896), .C1(new_n900), .C2(new_n889), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n894), .A2(new_n901), .ZN(G54));
  NAND3_X1  g716(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n903), .A2(new_n436), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n436), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n904), .A2(new_n905), .A3(new_n886), .ZN(G60));
  NAND2_X1  g720(.A1(new_n592), .A2(new_n593), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT59), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n899), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT118), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n910), .B1(new_n857), .B2(new_n860), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n886), .B1(new_n913), .B2(new_n907), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT118), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n899), .A2(new_n915), .A3(new_n908), .A4(new_n910), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n912), .A2(new_n914), .A3(new_n916), .ZN(G63));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT119), .Z(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT60), .Z(new_n920));
  AOI21_X1  g734(.A(KEYINPUT120), .B1(new_n897), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n922));
  INV_X1    g736(.A(new_n920), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n922), .B(new_n923), .C1(new_n858), .C2(new_n859), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n625), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NOR4_X1   g739(.A1(new_n850), .A2(new_n809), .A3(new_n810), .A4(new_n840), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n851), .A2(new_n853), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT53), .B1(new_n838), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n920), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n922), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n897), .A2(KEYINPUT120), .A3(new_n920), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n504), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n925), .A2(new_n932), .A3(new_n896), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n925), .A2(new_n932), .A3(KEYINPUT61), .A4(new_n896), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(G66));
  INV_X1    g751(.A(new_n191), .ZN(new_n938));
  OAI21_X1  g752(.A(G953), .B1(new_n938), .B2(new_n281), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n812), .A2(new_n824), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(G953), .ZN(new_n941));
  INV_X1    g755(.A(new_n252), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(G898), .B2(new_n390), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(G69));
  INV_X1    g758(.A(G900), .ZN(new_n945));
  OAI21_X1  g759(.A(G953), .B1(new_n305), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(KEYINPUT124), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n710), .A2(new_n805), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n750), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT123), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n722), .A2(new_n724), .ZN(new_n952));
  INV_X1    g766(.A(new_n748), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(new_n640), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n796), .A2(new_n632), .A3(new_n645), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n951), .A2(new_n390), .A3(new_n762), .A4(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n539), .B(new_n430), .ZN(new_n958));
  NAND2_X1  g772(.A1(G900), .A2(G953), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n820), .A2(new_n815), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n581), .A2(new_n719), .A3(new_n641), .A4(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n750), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n949), .B(new_n656), .C1(KEYINPUT121), .C2(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(KEYINPUT121), .B(KEYINPUT62), .Z(new_n966));
  INV_X1    g780(.A(new_n656), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(new_n948), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n963), .A2(new_n762), .A3(new_n965), .A4(new_n968), .ZN(new_n969));
  OR2_X1    g783(.A1(new_n969), .A2(KEYINPUT122), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(KEYINPUT122), .ZN(new_n971));
  AOI21_X1  g785(.A(G953), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n947), .B(new_n960), .C1(new_n972), .C2(new_n958), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n946), .A2(KEYINPUT124), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(G72));
  NAND2_X1  g789(.A1(new_n841), .A2(new_n856), .ZN(new_n976));
  NAND2_X1  g790(.A1(G472), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT63), .Z(new_n978));
  NAND2_X1  g792(.A1(new_n648), .A2(new_n554), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(KEYINPUT127), .A3(new_n542), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n979), .A2(KEYINPUT127), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n976), .A2(new_n978), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n970), .A2(new_n940), .A3(new_n971), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n978), .B(KEYINPUT125), .Z(new_n984));
  AOI21_X1  g798(.A(new_n649), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT126), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n951), .A2(new_n762), .A3(new_n940), .A4(new_n956), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n987), .A2(new_n984), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n986), .B(new_n896), .C1(new_n988), .C2(new_n577), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n577), .B1(new_n987), .B2(new_n984), .ZN(new_n990));
  OAI21_X1  g804(.A(KEYINPUT126), .B1(new_n990), .B2(new_n886), .ZN(new_n991));
  AOI211_X1 g805(.A(new_n982), .B(new_n985), .C1(new_n989), .C2(new_n991), .ZN(G57));
endmodule


