//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT32), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT25), .ZN(new_n204));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT24), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G183gat), .B2(G190gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n206), .B(new_n209), .C1(G183gat), .C2(G190gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(G169gat), .B2(G176gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n208), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(KEYINPUT23), .ZN(new_n215));
  XOR2_X1   g014(.A(new_n215), .B(KEYINPUT65), .Z(new_n216));
  OAI21_X1  g015(.A(new_n204), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(KEYINPUT67), .A2(G190gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n223), .A2(KEYINPUT68), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n224), .A2(new_n225), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(new_n222), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n206), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n231), .A2(KEYINPUT25), .A3(new_n213), .A4(new_n215), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(KEYINPUT27), .B(G183gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n229), .A2(new_n234), .A3(KEYINPUT28), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n220), .A2(KEYINPUT27), .A3(new_n221), .ZN(new_n236));
  OR2_X1    g035(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n226), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  XOR2_X1   g037(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n239));
  OAI21_X1  g038(.A(new_n235), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(KEYINPUT70), .B(new_n235), .C1(new_n238), .C2(new_n239), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n245));
  INV_X1    g044(.A(G169gat), .ZN(new_n246));
  INV_X1    g045(.A(G176gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NOR3_X1   g047(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n205), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT71), .B1(new_n244), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT71), .ZN(new_n253));
  AOI211_X1 g052(.A(new_n253), .B(new_n250), .C1(new_n242), .C2(new_n243), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n233), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G113gat), .ZN(new_n256));
  INV_X1    g055(.A(G120gat), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT1), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n258), .B1(new_n256), .B2(new_n257), .ZN(new_n259));
  OR2_X1    g058(.A1(G127gat), .A2(G134gat), .ZN(new_n260));
  INV_X1    g059(.A(G127gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT72), .B(G134gat), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n259), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264));
  XOR2_X1   g063(.A(KEYINPUT73), .B(G120gat), .Z(new_n265));
  OAI211_X1 g064(.A(new_n258), .B(new_n264), .C1(new_n265), .C2(new_n256), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n255), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G227gat), .ZN(new_n270));
  INV_X1    g069(.A(G233gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n233), .B(new_n267), .C1(new_n252), .C2(new_n254), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT74), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT74), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n269), .A2(new_n276), .A3(new_n272), .A4(new_n273), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n203), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT33), .ZN(new_n279));
  XNOR2_X1  g078(.A(G15gat), .B(G43gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(G71gat), .ZN(new_n281));
  INV_X1    g080(.A(G99gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n278), .B1(new_n279), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n275), .A2(new_n277), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n279), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT75), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT33), .B1(new_n275), .B2(new_n277), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT75), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n283), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n286), .A2(KEYINPUT32), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT76), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT76), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n285), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n269), .A2(new_n273), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(new_n270), .B2(new_n271), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT77), .B(KEYINPUT34), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n300), .B(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n298), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n304), .A2(new_n291), .A3(new_n294), .A4(new_n296), .ZN(new_n305));
  INV_X1    g104(.A(new_n302), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n285), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  XOR2_X1   g107(.A(G141gat), .B(G148gat), .Z(new_n309));
  INV_X1    g108(.A(KEYINPUT81), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(KEYINPUT82), .B2(KEYINPUT2), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n309), .B(new_n311), .C1(new_n310), .C2(KEYINPUT2), .ZN(new_n312));
  NAND2_X1  g111(.A1(G155gat), .A2(G162gat), .ZN(new_n313));
  INV_X1    g112(.A(G155gat), .ZN(new_n314));
  INV_X1    g113(.A(G162gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n313), .B1(new_n316), .B2(KEYINPUT2), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT82), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n309), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G197gat), .B(G204gat), .ZN(new_n322));
  INV_X1    g121(.A(G211gat), .ZN(new_n323));
  INV_X1    g122(.A(G218gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n322), .B1(KEYINPUT22), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G211gat), .B(G218gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(KEYINPUT29), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n321), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT83), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n330), .A2(new_n331), .B1(G228gat), .B2(G233gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n328), .B1(new_n333), .B2(KEYINPUT29), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n330), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n332), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(G22gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G78gat), .B(G106gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT31), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(G50gat), .ZN(new_n340));
  OR3_X1    g139(.A1(new_n337), .A2(KEYINPUT84), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n336), .A2(KEYINPUT84), .A3(G22gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(new_n340), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT30), .ZN(new_n346));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(KEYINPUT78), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n255), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n328), .ZN(new_n350));
  INV_X1    g149(.A(new_n348), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n217), .A2(new_n232), .B1(new_n244), .B2(new_n251), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(KEYINPUT29), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT79), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n348), .B1(new_n255), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n352), .A2(new_n351), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n328), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n349), .A2(new_n353), .A3(new_n360), .A4(new_n350), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n355), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G8gat), .B(G36gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT80), .ZN(new_n364));
  INV_X1    g163(.A(G64gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G92gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n346), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n362), .B2(new_n368), .ZN(new_n370));
  OR3_X1    g169(.A1(new_n362), .A2(KEYINPUT30), .A3(new_n368), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n333), .A2(new_n268), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OR3_X1    g175(.A1(new_n321), .A2(KEYINPUT4), .A3(new_n267), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n268), .A2(new_n317), .A3(new_n320), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT4), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n376), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n321), .B(new_n268), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(new_n381), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT5), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT5), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G1gat), .B(G29gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT0), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n392), .B(G57gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(G85gat), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT6), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n374), .A2(new_n375), .B1(new_n377), .B2(new_n379), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n384), .B1(new_n397), .B2(new_n381), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n389), .B(new_n394), .C1(new_n398), .C2(new_n388), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n396), .B(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n373), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n308), .A2(new_n345), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT35), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n344), .B1(new_n303), .B2(new_n307), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT35), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n399), .A2(KEYINPUT86), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n387), .A2(new_n408), .A3(new_n394), .A4(new_n389), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n410), .A2(new_n396), .B1(KEYINPUT6), .B2(new_n400), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n405), .A2(new_n406), .A3(new_n412), .A4(new_n372), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT36), .ZN(new_n414));
  INV_X1    g213(.A(new_n285), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n283), .B1(new_n290), .B2(KEYINPUT75), .ZN(new_n416));
  AOI211_X1 g215(.A(new_n288), .B(KEYINPUT33), .C1(new_n275), .C2(new_n277), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n278), .B(KEYINPUT76), .ZN(new_n419));
  AOI211_X1 g218(.A(new_n415), .B(new_n302), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n306), .B1(new_n305), .B2(new_n285), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n303), .A2(KEYINPUT36), .A3(new_n307), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n401), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n425), .A2(new_n344), .A3(new_n372), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n383), .A2(new_n381), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT39), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n428), .B(KEYINPUT85), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n397), .A2(new_n381), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n430), .A2(KEYINPUT39), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n395), .A3(new_n432), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n433), .A2(KEYINPUT40), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(KEYINPUT40), .ZN(new_n435));
  AOI22_X1  g234(.A1(new_n434), .A2(new_n435), .B1(new_n407), .B2(new_n409), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT37), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n355), .A2(new_n359), .A3(new_n437), .A4(new_n361), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT87), .B(KEYINPUT38), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n350), .B1(new_n357), .B2(new_n358), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n349), .A2(new_n328), .A3(new_n353), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(KEYINPUT37), .A3(new_n442), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n438), .A2(new_n368), .A3(new_n440), .A4(new_n443), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n411), .A2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n362), .A2(new_n368), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n362), .A2(KEYINPUT37), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n447), .A2(new_n438), .A3(new_n368), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n446), .B1(new_n448), .B2(new_n439), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n373), .A2(new_n436), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n426), .B1(new_n450), .B2(new_n344), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n404), .A2(new_n413), .B1(new_n424), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(G29gat), .A2(G36gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n453), .B(KEYINPUT14), .Z(new_n454));
  XNOR2_X1  g253(.A(G43gat), .B(G50gat), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n455), .A2(KEYINPUT15), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(KEYINPUT15), .ZN(new_n457));
  NAND2_X1  g256(.A1(G29gat), .A2(G36gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT91), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n454), .A2(new_n456), .A3(new_n457), .A4(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT92), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n453), .B(KEYINPUT14), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n463), .A2(KEYINPUT90), .B1(G29gat), .B2(G36gat), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(KEYINPUT90), .B2(new_n463), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(KEYINPUT15), .A3(new_n455), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(KEYINPUT17), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT16), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n469), .B1(new_n470), .B2(G1gat), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n471), .B1(G1gat), .B2(new_n469), .ZN(new_n472));
  INV_X1    g271(.A(G8gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(KEYINPUT93), .ZN(new_n476));
  INV_X1    g275(.A(new_n467), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G229gat), .A2(G233gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT18), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT95), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(KEYINPUT95), .A3(new_n483), .ZN(new_n487));
  XNOR2_X1  g286(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT89), .ZN(new_n489));
  XNOR2_X1  g288(.A(G113gat), .B(G141gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  XOR2_X1   g290(.A(G169gat), .B(G197gat), .Z(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n493), .B(KEYINPUT12), .Z(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n479), .B1(G229gat), .B2(G233gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n476), .B(new_n467), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n481), .B(KEYINPUT13), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n496), .A2(KEYINPUT18), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n486), .A2(new_n487), .A3(new_n495), .A4(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT96), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n503), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n484), .B(KEYINPUT94), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(new_n501), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n494), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n202), .B1(new_n452), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n451), .A2(new_n423), .A3(new_n422), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n345), .B(new_n372), .C1(new_n420), .C2(new_n421), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n514), .A2(KEYINPUT35), .A3(new_n411), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n406), .B1(new_n405), .B2(new_n402), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT97), .A3(new_n510), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT102), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g320(.A1(G85gat), .A2(G92gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n521), .A2(new_n522), .B1(KEYINPUT8), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT102), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n525), .A2(new_n527), .A3(G85gat), .A4(G92gat), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n524), .B(new_n528), .C1(G85gat), .C2(G92gat), .ZN(new_n529));
  XOR2_X1   g328(.A(G99gat), .B(G106gat), .Z(new_n530));
  OR2_X1    g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n468), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n533), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n467), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G190gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(new_n324), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT103), .ZN(new_n542));
  XOR2_X1   g341(.A(G134gat), .B(G162gat), .Z(new_n543));
  AOI21_X1  g342(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n540), .B(G218gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT103), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n542), .A2(new_n549), .A3(new_n545), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G57gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n552), .A2(G64gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n365), .A2(G57gat), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT9), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  INV_X1    g355(.A(G71gat), .ZN(new_n557));
  INV_X1    g356(.A(G78gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n556), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT98), .B1(new_n365), .B2(G57gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(new_n552), .A3(G64gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n562), .B1(new_n566), .B2(new_n553), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT99), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(KEYINPUT100), .B(KEYINPUT21), .Z(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n569), .A2(KEYINPUT21), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n476), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n476), .B2(new_n572), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n575), .B(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(new_n261), .ZN(new_n581));
  XNOR2_X1  g380(.A(KEYINPUT101), .B(G155gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n579), .B(new_n583), .Z(new_n584));
  NAND2_X1  g383(.A1(new_n551), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g384(.A1(new_n531), .A2(new_n568), .A3(new_n532), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n586), .B1(new_n570), .B2(new_n533), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT10), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n569), .A2(KEYINPUT10), .A3(new_n535), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT104), .ZN(new_n592));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT105), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G176gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G204gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n587), .A2(new_n593), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n594), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n598), .B(KEYINPUT106), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n591), .A2(new_n593), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n602), .B1(new_n603), .B2(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n585), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n519), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n401), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g408(.A1(new_n519), .A2(new_n606), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(new_n372), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n470), .A2(new_n473), .ZN(new_n612));
  NAND2_X1  g411(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n611), .B2(new_n473), .ZN(new_n615));
  MUX2_X1   g414(.A(new_n614), .B(new_n615), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g415(.A(KEYINPUT107), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n422), .A2(new_n617), .A3(new_n423), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n617), .B1(new_n422), .B2(new_n423), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n607), .A2(G15gat), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(G15gat), .B1(new_n607), .B2(new_n308), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(G1326gat));
  NAND3_X1  g422(.A1(new_n607), .A2(KEYINPUT108), .A3(new_n344), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT108), .B1(new_n607), .B2(new_n344), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT43), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n607), .A2(new_n344), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT108), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n624), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n627), .A2(G22gat), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g432(.A(G22gat), .B1(new_n627), .B2(new_n632), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(G1327gat));
  INV_X1    g434(.A(new_n551), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n584), .A2(new_n605), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT109), .Z(new_n639));
  AND2_X1   g438(.A1(new_n519), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(G29gat), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n640), .A2(new_n641), .A3(new_n401), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  AND2_X1   g443(.A1(new_n510), .A2(new_n637), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n517), .A2(KEYINPUT44), .A3(new_n636), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n451), .B1(new_n618), .B2(new_n619), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n404), .A2(new_n413), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n551), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n645), .B(new_n646), .C1(new_n649), .C2(KEYINPUT44), .ZN(new_n650));
  OAI21_X1  g449(.A(G29gat), .B1(new_n650), .B2(new_n425), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n644), .A2(new_n651), .ZN(G1328gat));
  INV_X1    g451(.A(G36gat), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n640), .A2(new_n653), .A3(new_n373), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(KEYINPUT46), .Z(new_n655));
  OAI21_X1  g454(.A(G36gat), .B1(new_n650), .B2(new_n372), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(G1329gat));
  AND2_X1   g456(.A1(new_n640), .A2(new_n308), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n620), .A2(G43gat), .ZN(new_n659));
  OAI22_X1  g458(.A1(new_n658), .A2(G43gat), .B1(new_n650), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g460(.A(G50gat), .B1(new_n650), .B2(new_n345), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT111), .ZN(new_n663));
  INV_X1    g462(.A(G50gat), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n519), .A2(new_n664), .A3(new_n639), .A4(new_n344), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT111), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n666), .B(G50gat), .C1(new_n650), .C2(new_n345), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT48), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n662), .A2(KEYINPUT48), .A3(new_n665), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT112), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n662), .A2(KEYINPUT112), .A3(KEYINPUT48), .A4(new_n665), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT113), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT113), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n670), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(G1331gat));
  AOI21_X1  g479(.A(new_n585), .B1(new_n647), .B2(new_n648), .ZN(new_n681));
  INV_X1    g480(.A(new_n605), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n510), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n425), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(new_n552), .ZN(G1332gat));
  INV_X1    g485(.A(new_n684), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n372), .B(KEYINPUT114), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT49), .B(G64gat), .Z(new_n692));
  OAI21_X1  g491(.A(new_n691), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT115), .ZN(G1333gat));
  AOI21_X1  g493(.A(G71gat), .B1(new_n687), .B2(new_n308), .ZN(new_n695));
  INV_X1    g494(.A(new_n620), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n684), .A2(new_n557), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n345), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(new_n558), .ZN(G1335gat));
  OR2_X1    g500(.A1(new_n649), .A2(KEYINPUT44), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n510), .A2(new_n584), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n702), .A2(new_n646), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n682), .A2(new_n425), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G85gat), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n649), .A2(new_n703), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT51), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n706), .A2(G85gat), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(G1336gat));
  NAND4_X1  g510(.A1(new_n702), .A2(new_n605), .A3(new_n646), .A4(new_n703), .ZN(new_n712));
  OAI21_X1  g511(.A(G92gat), .B1(new_n712), .B2(new_n688), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT52), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n689), .A2(new_n367), .A3(new_n605), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n713), .B(new_n714), .C1(new_n709), .C2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n712), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n367), .B1(new_n717), .B2(new_n373), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n708), .A2(KEYINPUT117), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n709), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT51), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n708), .A2(KEYINPUT117), .A3(new_n721), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n715), .B(KEYINPUT116), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n718), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n716), .B1(new_n725), .B2(new_n714), .ZN(G1337gat));
  OAI21_X1  g525(.A(G99gat), .B1(new_n712), .B2(new_n696), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n308), .A2(new_n282), .A3(new_n605), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n709), .B2(new_n728), .ZN(G1338gat));
  OR3_X1    g528(.A1(new_n712), .A2(KEYINPUT119), .A3(new_n345), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT119), .B1(new_n712), .B2(new_n345), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(G106gat), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT53), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n345), .A2(new_n682), .A3(G106gat), .ZN(new_n734));
  INV_X1    g533(.A(new_n734), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n732), .B(new_n733), .C1(new_n709), .C2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n722), .A3(new_n734), .ZN(new_n737));
  OAI21_X1  g536(.A(G106gat), .B1(new_n712), .B2(new_n345), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT118), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g539(.A(KEYINPUT118), .B(G106gat), .C1(new_n712), .C2(new_n345), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n737), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT53), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n736), .A2(new_n743), .ZN(G1339gat));
  XNOR2_X1  g543(.A(KEYINPUT120), .B(G113gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(KEYINPUT120), .A2(G113gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n480), .A2(new_n481), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n498), .A2(new_n500), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n493), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n750), .B1(new_n504), .B2(new_n505), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n751), .A2(new_n605), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n594), .B(KEYINPUT54), .C1(new_n593), .C2(new_n591), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT54), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n598), .B1(new_n603), .B2(new_n755), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n753), .B2(new_n756), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n601), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n506), .B2(new_n509), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n551), .B1(new_n752), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n759), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n636), .A2(new_n751), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n584), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n585), .A2(new_n510), .A3(new_n605), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n405), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n401), .A3(new_n688), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n511), .ZN(new_n770));
  MUX2_X1   g569(.A(new_n745), .B(new_n746), .S(new_n770), .Z(G1340gat));
  NOR2_X1   g570(.A1(new_n769), .A2(new_n682), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n265), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n257), .B2(new_n772), .ZN(G1341gat));
  INV_X1    g573(.A(new_n584), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n769), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT121), .A2(G127gat), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1342gat));
  INV_X1    g577(.A(new_n766), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n779), .A2(new_n401), .A3(new_n372), .A4(new_n636), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n781), .A2(new_n262), .A3(new_n405), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT56), .Z(new_n783));
  OAI21_X1  g582(.A(G134gat), .B1(new_n769), .B2(new_n551), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1343gat));
  NOR3_X1   g584(.A1(new_n620), .A2(new_n425), .A3(new_n689), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n761), .A2(KEYINPUT122), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT122), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n788), .B(new_n551), .C1(new_n752), .C2(new_n760), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(new_n763), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n765), .B1(new_n790), .B2(new_n775), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n791), .A2(new_n792), .A3(new_n345), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n766), .B2(new_n345), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n510), .B(new_n786), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G141gat), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n766), .A2(new_n345), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n798), .A2(new_n786), .ZN(new_n799));
  INV_X1    g598(.A(G141gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n800), .A3(new_n510), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n801), .B2(KEYINPUT123), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n797), .B(new_n801), .C1(KEYINPUT123), .C2(new_n803), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1344gat));
  INV_X1    g606(.A(G148gat), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n799), .A2(new_n808), .A3(new_n605), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810));
  OAI211_X1 g609(.A(KEYINPUT57), .B(new_n344), .C1(new_n764), .C2(new_n765), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n682), .B1(new_n794), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n786), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT124), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n808), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(KEYINPUT124), .A3(new_n786), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n810), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n605), .B(new_n786), .C1(new_n793), .C2(new_n795), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n818), .A2(new_n810), .A3(G148gat), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n809), .B1(new_n817), .B2(new_n819), .ZN(G1345gat));
  OAI21_X1  g619(.A(new_n786), .B1(new_n793), .B2(new_n795), .ZN(new_n821));
  OAI21_X1  g620(.A(G155gat), .B1(new_n821), .B2(new_n775), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n799), .A2(new_n314), .A3(new_n584), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1346gat));
  OAI211_X1 g623(.A(new_n636), .B(new_n786), .C1(new_n793), .C2(new_n795), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(G162gat), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n620), .A2(new_n345), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n781), .A2(new_n315), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT125), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT125), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n826), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1347gat));
  NAND3_X1  g632(.A1(new_n779), .A2(new_n425), .A3(new_n689), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n767), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n246), .A3(new_n510), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n372), .A2(new_n401), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n768), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(G169gat), .B1(new_n838), .B2(new_n511), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n839), .ZN(G1348gat));
  NOR3_X1   g639(.A1(new_n838), .A2(new_n247), .A3(new_n682), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n835), .A2(new_n605), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n247), .ZN(G1349gat));
  NAND3_X1  g642(.A1(new_n835), .A2(new_n234), .A3(new_n584), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n223), .B1(new_n838), .B2(new_n775), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g646(.A1(new_n835), .A2(new_n229), .A3(new_n636), .ZN(new_n848));
  OAI21_X1  g647(.A(G190gat), .B1(new_n838), .B2(new_n551), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n849), .A2(KEYINPUT61), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(KEYINPUT61), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(G1351gat));
  NAND2_X1  g651(.A1(new_n794), .A2(new_n811), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n696), .A2(new_n837), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT126), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n510), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G197gat), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n834), .A2(new_n345), .A3(new_n620), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n511), .A2(G197gat), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(G1352gat));
  INV_X1    g661(.A(G204gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n859), .A2(new_n863), .A3(new_n605), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT62), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(KEYINPUT62), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n812), .A2(new_n855), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n865), .B(new_n866), .C1(new_n863), .C2(new_n867), .ZN(G1353gat));
  NAND3_X1  g667(.A1(new_n853), .A2(new_n584), .A3(new_n855), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT63), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT127), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(G211gat), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n870), .A2(KEYINPUT127), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n859), .A2(new_n323), .A3(new_n584), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n872), .A2(new_n873), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(G1354gat));
  AOI21_X1  g676(.A(G218gat), .B1(new_n859), .B2(new_n636), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n551), .A2(new_n324), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n856), .B2(new_n879), .ZN(G1355gat));
endmodule


