//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n445, new_n446, new_n451, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n565, new_n567, new_n568, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1162, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  INV_X1    g018(.A(G2072), .ZN(new_n444));
  INV_X1    g019(.A(G2078), .ZN(new_n445));
  NOR2_X1   g020(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g021(.A1(new_n446), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g027(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G325));
  XOR2_X1   g033(.A(G325), .B(KEYINPUT66), .Z(G261));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT67), .Z(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G125), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n467), .A2(new_n468), .B1(G113), .B2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(KEYINPUT68), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n471), .A2(G2105), .ZN(new_n479));
  AOI22_X1  g054(.A1(new_n478), .A2(G137), .B1(G101), .B2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n477), .A2(new_n480), .ZN(G160));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n482), .B1(new_n472), .B2(new_n473), .ZN(new_n483));
  AOI22_X1  g058(.A1(G124), .A2(new_n483), .B1(new_n478), .B2(G136), .ZN(new_n484));
  INV_X1    g059(.A(G100), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n485), .A2(new_n482), .A3(KEYINPUT69), .ZN(new_n486));
  AOI21_X1  g061(.A(KEYINPUT69), .B1(new_n485), .B2(new_n482), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G112), .B2(new_n482), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n465), .B2(new_n466), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n474), .A2(KEYINPUT71), .A3(new_n492), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n493), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT70), .B1(new_n482), .B2(G114), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(G126), .A2(new_n483), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n497), .A2(new_n499), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n514), .A2(KEYINPUT72), .A3(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n510), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n513), .A2(new_n515), .B1(KEYINPUT5), .B2(new_n512), .ZN(new_n523));
  INV_X1    g098(.A(new_n521), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(KEYINPUT73), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT74), .B(G88), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(G75), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G62), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n518), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n521), .A2(new_n512), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n531), .A2(G651), .B1(G50), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n528), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  XNOR2_X1  g110(.A(KEYINPUT75), .B(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n526), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(G76), .A2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G651), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n524), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G51), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G63), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n518), .A2(new_n545), .B1(new_n538), .B2(new_n539), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n544), .B1(G651), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n537), .A2(new_n547), .ZN(G168));
  AOI22_X1  g123(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n549), .B2(KEYINPUT76), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(KEYINPUT76), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n532), .A2(G52), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n522), .A2(new_n525), .ZN(new_n553));
  INV_X1    g128(.A(G90), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n551), .A2(new_n555), .ZN(G171));
  NAND2_X1  g131(.A1(new_n526), .A2(G81), .ZN(new_n557));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n518), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n560), .A2(G651), .B1(G43), .B2(new_n532), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  INV_X1    g144(.A(KEYINPUT78), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G53), .ZN(new_n571));
  OR3_X1    g146(.A1(new_n542), .A2(KEYINPUT9), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(KEYINPUT9), .B1(new_n542), .B2(new_n571), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G65), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n518), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n572), .A2(new_n573), .B1(G651), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n526), .A2(G91), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G299));
  OR2_X1    g154(.A1(new_n551), .A2(new_n555), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT79), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  NAND2_X1  g157(.A1(G171), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G301));
  INV_X1    g160(.A(G168), .ZN(G286));
  NAND2_X1  g161(.A1(new_n526), .A2(G87), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n523), .A2(G74), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(G49), .B2(new_n532), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n587), .A2(new_n589), .ZN(G288));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n518), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n593), .A2(G651), .B1(G48), .B2(new_n532), .ZN(new_n594));
  INV_X1    g169(.A(G86), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(new_n553), .ZN(G305));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n518), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G47), .B2(new_n532), .ZN(new_n600));
  INV_X1    g175(.A(G85), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n553), .ZN(G290));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(KEYINPUT81), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n603), .A2(KEYINPUT81), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n604), .B(new_n605), .C1(new_n518), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G651), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n532), .A2(G54), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n553), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n610), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT80), .B1(new_n615), .B2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n584), .A2(new_n617), .ZN(new_n618));
  MUX2_X1   g193(.A(new_n616), .B(KEYINPUT80), .S(new_n618), .Z(G321));
  XNOR2_X1  g194(.A(G321), .B(KEYINPUT82), .ZN(G284));
  NOR2_X1   g195(.A1(G286), .A2(new_n617), .ZN(new_n621));
  XOR2_X1   g196(.A(G299), .B(KEYINPUT83), .Z(new_n622));
  AOI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n617), .ZN(G297));
  AOI21_X1  g198(.A(new_n621), .B1(new_n622), .B2(new_n617), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n615), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND3_X1  g201(.A1(new_n615), .A2(KEYINPUT84), .A3(new_n625), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(KEYINPUT84), .B1(new_n615), .B2(new_n625), .ZN(new_n629));
  NOR3_X1   g204(.A1(new_n628), .A2(new_n617), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(new_n617), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n474), .A2(new_n479), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT85), .B(KEYINPUT12), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(G2100), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  AOI22_X1  g214(.A1(G123), .A2(new_n483), .B1(new_n478), .B2(G135), .ZN(new_n640));
  NOR3_X1   g215(.A1(new_n482), .A2(KEYINPUT86), .A3(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(KEYINPUT86), .B1(new_n482), .B2(G111), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n642), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n640), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n638), .A2(new_n639), .A3(new_n645), .ZN(G156));
  INV_X1    g221(.A(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2430), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT87), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n659), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n660), .A2(new_n661), .A3(G14), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT88), .ZN(new_n665));
  NOR2_X1   g240(.A1(G2072), .A2(G2078), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n446), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n663), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(KEYINPUT17), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n668), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n663), .B(new_n664), .C1(new_n446), .C2(new_n666), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n671), .B(KEYINPUT18), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n665), .A3(new_n663), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT20), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NOR3_X1   g259(.A1(new_n678), .A2(new_n681), .A3(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(new_n678), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT89), .Z(new_n688));
  XOR2_X1   g263(.A(G1981), .B(G1986), .Z(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n688), .B(new_n693), .ZN(G229));
  XOR2_X1   g269(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n695));
  NAND3_X1  g270(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n478), .A2(G139), .ZN(new_n698));
  AOI22_X1  g273(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n697), .B(new_n698), .C1(new_n482), .C2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT93), .Z(new_n701));
  MUX2_X1   g276(.A(G33), .B(new_n701), .S(G29), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(new_n444), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT95), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G29), .B2(G32), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n478), .A2(G141), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT94), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n483), .A2(G129), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT26), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n479), .A2(G105), .ZN(new_n711));
  AND4_X1   g286(.A1(new_n707), .A2(new_n708), .A3(new_n710), .A4(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G29), .ZN(new_n713));
  MUX2_X1   g288(.A(new_n704), .B(new_n705), .S(new_n713), .Z(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT24), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(G34), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n717), .B2(G34), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G160), .B2(G29), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n714), .A2(new_n715), .B1(G2084), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n703), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT96), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NOR2_X1   g299(.A1(G168), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n724), .B2(G21), .ZN(new_n726));
  INV_X1    g301(.A(G1966), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n563), .A2(new_n724), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n724), .B2(G19), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n728), .B1(G1341), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G1341), .B2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n716), .A2(G35), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G162), .B2(new_n716), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT29), .ZN(new_n736));
  INV_X1    g311(.A(G2090), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  OAI221_X1 g313(.A(new_n738), .B1(G2084), .B2(new_n720), .C1(new_n715), .C2(new_n714), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n726), .A2(new_n727), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n478), .A2(G140), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n483), .A2(G128), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n482), .A2(G116), .ZN(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n716), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(G2067), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT30), .B(G28), .ZN(new_n752));
  OR2_X1    g327(.A1(KEYINPUT31), .A2(G11), .ZN(new_n753));
  NAND2_X1  g328(.A1(KEYINPUT31), .A2(G11), .ZN(new_n754));
  AOI22_X1  g329(.A1(new_n752), .A2(new_n716), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n644), .B2(new_n716), .ZN(new_n756));
  NOR2_X1   g331(.A1(G164), .A2(new_n716), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G27), .B2(new_n716), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n756), .B1(new_n758), .B2(new_n445), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n445), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n740), .A2(new_n751), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n733), .A2(new_n739), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n724), .A2(G4), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n615), .B2(new_n724), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1348), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n724), .A2(G20), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT23), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G299), .B2(G16), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G1956), .Z(new_n769));
  NAND2_X1  g344(.A1(new_n724), .A2(G5), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G171), .B2(new_n724), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1961), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n765), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n723), .A2(new_n762), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n724), .A2(G23), .ZN(new_n775));
  INV_X1    g350(.A(G288), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(new_n724), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT33), .B(G1976), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n724), .A2(G22), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G166), .B2(new_n724), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT91), .Z(new_n782));
  AOI21_X1  g357(.A(new_n779), .B1(new_n782), .B2(G1971), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G1971), .B2(new_n782), .ZN(new_n784));
  MUX2_X1   g359(.A(G6), .B(G305), .S(G16), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT32), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1981), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT34), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(KEYINPUT34), .B1(new_n784), .B2(new_n787), .ZN(new_n791));
  INV_X1    g366(.A(G290), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(new_n724), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n724), .B2(G24), .ZN(new_n794));
  INV_X1    g369(.A(G1986), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n478), .A2(G131), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n483), .A2(G119), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n482), .A2(G107), .ZN(new_n800));
  OAI21_X1  g375(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n798), .B(new_n799), .C1(new_n800), .C2(new_n801), .ZN(new_n802));
  MUX2_X1   g377(.A(G25), .B(new_n802), .S(G29), .Z(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT35), .B(G1991), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT90), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n803), .B(new_n805), .Z(new_n806));
  NAND3_X1  g381(.A1(new_n796), .A2(new_n797), .A3(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n790), .A2(new_n791), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT36), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n807), .B1(new_n788), .B2(new_n789), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT36), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n811), .A2(new_n812), .A3(new_n791), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n774), .B1(new_n810), .B2(new_n813), .ZN(G311));
  INV_X1    g389(.A(new_n774), .ZN(new_n815));
  AND3_X1   g390(.A1(new_n811), .A2(new_n812), .A3(new_n791), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n812), .B1(new_n811), .B2(new_n791), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n815), .B1(new_n816), .B2(new_n817), .ZN(G150));
  AOI22_X1  g393(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  OAI21_X1  g394(.A(G651), .B1(new_n819), .B2(KEYINPUT97), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(KEYINPUT97), .B2(new_n819), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n532), .A2(G55), .ZN(new_n822));
  INV_X1    g397(.A(G93), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n553), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(G860), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n615), .A2(G559), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT98), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n825), .B(new_n562), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n833), .A2(KEYINPUT39), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n826), .B1(new_n833), .B2(KEYINPUT39), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n828), .B1(new_n834), .B2(new_n835), .ZN(G145));
  XNOR2_X1  g411(.A(G160), .B(KEYINPUT99), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G162), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n644), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n508), .B(new_n745), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n712), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(new_n700), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n701), .B2(new_n841), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n635), .B(new_n802), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n483), .A2(G130), .ZN(new_n845));
  OR2_X1    g420(.A1(G106), .A2(G2105), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(G2104), .C1(G118), .C2(new_n482), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G142), .B2(new_n478), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n844), .B(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n850), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n842), .B(new_n852), .C1(new_n701), .C2(new_n841), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n839), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT100), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n839), .B1(new_n851), .B2(new_n853), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(G37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g434(.A(new_n615), .ZN(new_n860));
  INV_X1    g435(.A(G299), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n615), .A2(G299), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(KEYINPUT101), .A3(new_n863), .ZN(new_n864));
  OR3_X1    g439(.A1(new_n860), .A2(KEYINPUT101), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n563), .B(new_n825), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n628), .B2(new_n629), .ZN(new_n868));
  INV_X1    g443(.A(new_n629), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n832), .A2(new_n869), .A3(new_n627), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n866), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n866), .A2(KEYINPUT41), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n862), .A2(new_n874), .A3(new_n863), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n860), .A2(new_n861), .A3(KEYINPUT102), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n868), .A2(new_n870), .ZN(new_n880));
  OAI211_X1 g455(.A(KEYINPUT103), .B(new_n872), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT103), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n873), .B2(new_n878), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(new_n871), .ZN(new_n884));
  XOR2_X1   g459(.A(G288), .B(G305), .Z(new_n885));
  XNOR2_X1  g460(.A(new_n792), .B(G303), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT42), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n881), .A2(new_n884), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n883), .A2(new_n871), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n889), .B(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n894), .A3(KEYINPUT103), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(G868), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n897));
  INV_X1    g472(.A(new_n825), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n898), .B2(new_n617), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n891), .A2(new_n897), .A3(G868), .A4(new_n895), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(G295));
  AND2_X1   g477(.A1(new_n900), .A2(new_n901), .ZN(G331));
  NAND2_X1  g478(.A1(new_n584), .A2(G168), .ZN(new_n904));
  NOR2_X1   g479(.A1(G171), .A2(G168), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n867), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G286), .B1(new_n581), .B2(new_n583), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n832), .B1(new_n908), .B2(new_n905), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n866), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n873), .A2(new_n878), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n907), .A2(new_n909), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(G37), .B1(new_n913), .B2(new_n889), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n907), .A2(new_n909), .ZN(new_n915));
  INV_X1    g490(.A(new_n866), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n917), .B1(new_n879), .B2(new_n915), .ZN(new_n918));
  INV_X1    g493(.A(new_n889), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT43), .B1(new_n914), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n866), .B1(new_n915), .B2(new_n876), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n875), .A2(new_n877), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n907), .A2(new_n923), .A3(new_n909), .A4(KEYINPUT41), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n919), .A3(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n889), .B(new_n917), .C1(new_n879), .C2(new_n915), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  AND4_X1   g502(.A1(KEYINPUT43), .A2(new_n925), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT44), .B1(new_n921), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(new_n914), .B2(new_n920), .ZN(new_n932));
  AND4_X1   g507(.A1(new_n931), .A2(new_n925), .A3(new_n926), .A4(new_n927), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n934), .ZN(G397));
  INV_X1    g510(.A(G1384), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n495), .A2(KEYINPUT4), .A3(new_n496), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n504), .A2(new_n506), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n483), .A2(G126), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n499), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n936), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n942), .A2(KEYINPUT45), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n477), .A2(G40), .A3(new_n480), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n945), .B(KEYINPUT107), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n745), .B(new_n750), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT108), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(new_n712), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1996), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n950), .B1(new_n951), .B2(new_n948), .ZN(new_n952));
  INV_X1    g527(.A(new_n945), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(new_n951), .A3(new_n712), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT106), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n802), .B(new_n805), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT109), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n946), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n792), .A2(new_n795), .ZN(new_n960));
  NAND2_X1  g535(.A1(G290), .A2(G1986), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n961), .A3(KEYINPUT105), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n962), .B(new_n953), .C1(KEYINPUT105), .C2(new_n961), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n956), .A2(new_n959), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT111), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n965), .B(new_n936), .C1(new_n937), .C2(new_n940), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n965), .B1(new_n508), .B2(new_n936), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT50), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n970), .B(new_n936), .C1(new_n937), .C2(new_n940), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT115), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n508), .A2(KEYINPUT115), .A3(new_n970), .A4(new_n936), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n969), .A2(new_n944), .A3(new_n975), .ZN(new_n976));
  XOR2_X1   g551(.A(KEYINPUT120), .B(G1956), .Z(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(G299), .A2(KEYINPUT57), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT57), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n577), .B2(new_n578), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT110), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n508), .A2(new_n985), .A3(KEYINPUT45), .A4(new_n936), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n477), .A2(G40), .A3(new_n480), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n988), .B1(new_n989), .B2(new_n941), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(new_n444), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n987), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n978), .A2(new_n982), .A3(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n967), .A2(new_n968), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT122), .B1(new_n995), .B2(new_n944), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n941), .A2(KEYINPUT111), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n997), .A2(new_n944), .A3(KEYINPUT122), .A4(new_n966), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n750), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n970), .A3(new_n966), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n941), .A2(KEYINPUT50), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1001), .A2(new_n1002), .A3(new_n944), .ZN(new_n1003));
  INV_X1    g578(.A(G1348), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n860), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n982), .B1(new_n978), .B2(new_n993), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n994), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT61), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n978), .A2(new_n982), .A3(new_n993), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(new_n1007), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT60), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n997), .A2(new_n944), .A3(new_n966), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT122), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(G2067), .B1(new_n1016), .B2(new_n998), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1012), .B1(new_n1013), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1000), .A2(KEYINPUT60), .A3(new_n1005), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n615), .ZN(new_n1020));
  INV_X1    g595(.A(new_n977), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n997), .A2(new_n966), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n988), .B1(new_n1022), .B2(KEYINPUT50), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1023), .B2(new_n975), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n990), .A2(new_n984), .A3(new_n986), .ZN(new_n1025));
  INV_X1    g600(.A(new_n992), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI22_X1  g602(.A1(new_n1024), .A2(new_n1027), .B1(new_n981), .B2(new_n979), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(KEYINPUT61), .A3(new_n994), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1011), .A2(new_n1020), .A3(new_n1029), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT58), .B(G1341), .Z(new_n1031));
  NAND3_X1  g606(.A1(new_n1016), .A2(new_n998), .A3(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT123), .B(G1996), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n987), .A2(new_n990), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n562), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT124), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(KEYINPUT59), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1000), .A2(KEYINPUT60), .A3(new_n860), .A4(new_n1005), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n1039));
  OAI211_X1 g614(.A(new_n1037), .B(new_n1038), .C1(new_n1035), .C2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1008), .B1(new_n1030), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(G303), .A2(G8), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1042), .B(KEYINPUT55), .ZN(new_n1043));
  INV_X1    g618(.A(G1971), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1025), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n969), .A2(new_n975), .A3(new_n737), .A4(new_n944), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  OAI211_X1 g623(.A(KEYINPUT116), .B(new_n1043), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1051));
  XOR2_X1   g626(.A(new_n1042), .B(KEYINPUT55), .Z(new_n1052));
  OAI21_X1  g627(.A(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G305), .A2(G1981), .ZN(new_n1055));
  INV_X1    g630(.A(G1981), .ZN(new_n1056));
  OAI211_X1 g631(.A(new_n594), .B(new_n1056), .C1(new_n595), .C2(new_n553), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT49), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1055), .A2(new_n1057), .A3(KEYINPUT49), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1060), .A2(G8), .A3(new_n1014), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G1976), .ZN(new_n1063));
  NOR2_X1   g638(.A1(G288), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT113), .B(G1976), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT52), .B1(G288), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1065), .A2(new_n1067), .A3(G8), .A4(new_n1014), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1014), .A2(G8), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT52), .B1(new_n1069), .B2(new_n1064), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1062), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1001), .A2(new_n737), .A3(new_n1002), .A4(new_n944), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1072), .A2(KEYINPUT112), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1072), .A2(KEYINPUT112), .B1(new_n1025), .B2(new_n1044), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1048), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1071), .B1(new_n1075), .B2(new_n1052), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1054), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT125), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n944), .A2(new_n983), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n989), .B1(new_n967), .B2(new_n968), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1966), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT117), .B(G2084), .Z(new_n1083));
  NOR2_X1   g658(.A1(new_n988), .A2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1001), .A2(new_n1002), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1078), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(G168), .A2(new_n1048), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT45), .B1(new_n997), .B2(new_n966), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n727), .B1(new_n1088), .B2(new_n1079), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1001), .A2(new_n1002), .A3(new_n1084), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(KEYINPUT125), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1086), .A2(new_n1087), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(G168), .ZN(new_n1095));
  OAI21_X1  g670(.A(G8), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1087), .A2(KEYINPUT51), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(KEYINPUT126), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT126), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1048), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1087), .A2(KEYINPUT51), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1092), .B1(new_n1095), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1025), .B2(G2078), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(G2078), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1080), .A2(new_n1081), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(G1961), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1003), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n584), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT127), .B1(new_n943), .B2(new_n988), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT127), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n990), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1113), .A2(new_n1115), .A3(new_n987), .A4(new_n1107), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(new_n1106), .A3(new_n1110), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1112), .B1(new_n584), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1111), .A2(new_n584), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1119), .B1(new_n1117), .B2(G171), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1118), .A2(new_n1119), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1041), .A2(new_n1077), .A3(new_n1104), .A4(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1104), .A2(KEYINPUT62), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1092), .B(new_n1125), .C1(new_n1095), .C2(new_n1103), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1112), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1054), .A2(new_n1076), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1075), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1130), .A2(new_n1043), .A3(new_n1071), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1062), .A2(new_n1063), .A3(new_n776), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1057), .B(KEYINPUT114), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1069), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1123), .A2(new_n1129), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1130), .A2(new_n1043), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT118), .B1(new_n1096), .B2(G286), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT118), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1100), .A2(new_n1139), .A3(G168), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  AND4_X1   g716(.A1(KEYINPUT63), .A2(new_n1137), .A3(new_n1076), .A4(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1054), .A2(new_n1076), .A3(new_n1141), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1143), .A2(KEYINPUT119), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT63), .B1(new_n1143), .B2(KEYINPUT119), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1142), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n964), .B1(new_n1136), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n953), .A2(new_n951), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT46), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n950), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT47), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n956), .A2(new_n959), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n945), .A2(new_n960), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT48), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1151), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n802), .A2(new_n805), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n956), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(G2067), .B2(new_n745), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1155), .B1(new_n946), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1147), .A2(new_n1159), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g735(.A1(new_n463), .A2(G227), .ZN(new_n1162));
  NOR3_X1   g736(.A1(G401), .A2(G229), .A3(new_n1162), .ZN(new_n1163));
  OAI211_X1 g737(.A(new_n1163), .B(new_n858), .C1(new_n932), .C2(new_n933), .ZN(G225));
  INV_X1    g738(.A(G225), .ZN(G308));
endmodule


