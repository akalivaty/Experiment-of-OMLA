//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004;
  AND2_X1   g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT82), .ZN(new_n204));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  INV_X1    g004(.A(G155gat), .ZN(new_n206));
  INV_X1    g005(.A(G162gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G141gat), .B(G148gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n205), .B(new_n208), .C1(new_n209), .C2(KEYINPUT2), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n211));
  INV_X1    g010(.A(G141gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G148gat), .ZN(new_n213));
  INV_X1    g012(.A(G148gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G155gat), .B(G162gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n205), .A2(KEYINPUT2), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n210), .A2(new_n211), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G211gat), .B(G218gat), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G211gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT72), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT72), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(G211gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT22), .B1(new_n230), .B2(G218gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(G197gat), .B(G204gat), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n225), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(G218gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n235), .B1(new_n227), .B2(new_n229), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n232), .B(new_n224), .C1(new_n236), .C2(KEYINPUT22), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n204), .B1(new_n223), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n237), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT22), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT72), .B(G211gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(new_n235), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n224), .B1(new_n243), .B2(new_n232), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n240), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n220), .A2(new_n222), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(KEYINPUT82), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT74), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n217), .B1(new_n218), .B2(new_n216), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n210), .A2(KEYINPUT74), .A3(new_n219), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n222), .B1(new_n240), .B2(new_n244), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n253), .B1(new_n254), .B2(new_n211), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n239), .B(new_n247), .C1(new_n255), .C2(KEYINPUT81), .ZN(new_n256));
  INV_X1    g055(.A(new_n253), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n221), .B1(new_n234), .B2(new_n237), .ZN(new_n258));
  OAI211_X1 g057(.A(new_n257), .B(KEYINPUT81), .C1(KEYINPUT3), .C2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  OAI211_X1 g059(.A(KEYINPUT83), .B(new_n203), .C1(new_n256), .C2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT85), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(new_n223), .B2(new_n238), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n245), .A2(KEYINPUT85), .A3(new_n246), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n203), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n210), .A2(new_n219), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT29), .B1(new_n234), .B2(new_n237), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT84), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n211), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AOI211_X1 g068(.A(KEYINPUT84), .B(KEYINPUT29), .C1(new_n234), .C2(new_n237), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n265), .A2(new_n271), .A3(KEYINPUT86), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT86), .B1(new_n265), .B2(new_n271), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n261), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT81), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n275), .B1(new_n276), .B2(new_n253), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n277), .A2(new_n259), .A3(new_n239), .A4(new_n247), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT83), .B1(new_n278), .B2(new_n203), .ZN(new_n279));
  OAI21_X1  g078(.A(G22gat), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n203), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT83), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n271), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT86), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n265), .A2(new_n271), .A3(KEYINPUT86), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(G22gat), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n283), .A2(new_n288), .A3(new_n289), .A4(new_n261), .ZN(new_n290));
  XNOR2_X1  g089(.A(G78gat), .B(G106gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT31), .B(G50gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n280), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n294), .A2(KEYINPUT88), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT88), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n280), .A2(new_n290), .A3(new_n296), .A4(new_n293), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n290), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n293), .B(KEYINPUT80), .Z(new_n300));
  AOI21_X1  g099(.A(KEYINPUT87), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT87), .ZN(new_n302));
  INV_X1    g101(.A(new_n300), .ZN(new_n303));
  AOI211_X1 g102(.A(new_n302), .B(new_n303), .C1(new_n280), .C2(new_n290), .ZN(new_n304));
  OAI22_X1  g103(.A1(new_n295), .A2(new_n298), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(KEYINPUT26), .ZN(new_n307));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n306), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT68), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT27), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(G183gat), .ZN(new_n317));
  INV_X1    g116(.A(G190gat), .ZN(new_n318));
  INV_X1    g117(.A(G183gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n317), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(G183gat), .B1(KEYINPUT67), .B2(KEYINPUT27), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n322), .B1(KEYINPUT67), .B2(KEYINPUT27), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n314), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT28), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n319), .A2(KEYINPUT27), .ZN(new_n326));
  AOI21_X1  g125(.A(G190gat), .B1(new_n326), .B2(new_n315), .ZN(new_n327));
  OR2_X1    g126(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n328));
  NAND2_X1  g127(.A1(KEYINPUT67), .A2(KEYINPUT27), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(G183gat), .A3(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n327), .A2(new_n330), .A3(KEYINPUT68), .A4(new_n320), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n324), .A2(new_n325), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n316), .A2(G183gat), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n326), .A2(new_n333), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n334), .A2(KEYINPUT28), .A3(new_n318), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n313), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n306), .A2(KEYINPUT23), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT23), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(G169gat), .B2(G176gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n308), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT65), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT24), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n319), .A2(G190gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n318), .A2(G183gat), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(G183gat), .A3(G190gat), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n343), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n349), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n347), .A2(KEYINPUT65), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n342), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(G183gat), .B(G190gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n349), .B1(new_n354), .B2(new_n344), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n341), .B1(new_n355), .B2(new_n340), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT64), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT64), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n358), .B(new_n341), .C1(new_n355), .C2(new_n340), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n353), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n336), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G226gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n363), .B1(new_n361), .B2(new_n222), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n245), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT29), .B1(new_n336), .B2(new_n360), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n364), .B(new_n238), .C1(new_n363), .C2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G8gat), .B(G36gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n371), .B(new_n372), .Z(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n367), .A2(new_n369), .A3(new_n373), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(KEYINPUT30), .A3(new_n376), .ZN(new_n377));
  OR3_X1    g176(.A1(new_n370), .A2(KEYINPUT30), .A3(new_n374), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G113gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G120gat), .ZN(new_n384));
  INV_X1    g183(.A(G120gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G113gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT1), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G127gat), .B(G134gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n385), .A2(KEYINPUT70), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT70), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(G120gat), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT71), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n393), .A2(new_n395), .A3(new_n396), .A4(G113gat), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(new_n388), .A3(new_n390), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n384), .A2(KEYINPUT71), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT70), .B(G120gat), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n399), .B1(new_n400), .B2(G113gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n392), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n402), .B(new_n266), .Z(new_n403));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n382), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n266), .A2(KEYINPUT3), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n406), .A2(new_n402), .A3(new_n220), .ZN(new_n407));
  INV_X1    g206(.A(new_n404), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n402), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n253), .A2(new_n410), .A3(KEYINPUT4), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n412), .B1(new_n402), .B2(new_n266), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n409), .A2(KEYINPUT75), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n415));
  INV_X1    g214(.A(new_n411), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n406), .A2(new_n402), .A3(new_n220), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(new_n413), .A3(new_n404), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n415), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n405), .B1(new_n414), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G1gat), .B(G29gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT0), .ZN(new_n422));
  XNOR2_X1  g221(.A(G57gat), .B(G85gat), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n422), .B(new_n423), .Z(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n253), .A2(new_n410), .A3(new_n412), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT4), .B1(new_n402), .B2(new_n266), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n409), .A2(new_n428), .A3(new_n381), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n420), .A2(new_n425), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT78), .ZN(new_n432));
  XOR2_X1   g231(.A(KEYINPUT77), .B(KEYINPUT6), .Z(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n425), .B1(new_n420), .B2(new_n429), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT79), .ZN(new_n437));
  INV_X1    g236(.A(new_n433), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT78), .B1(new_n430), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT79), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n434), .A2(new_n437), .A3(new_n439), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n436), .A2(new_n438), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n380), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n361), .A2(new_n410), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n336), .A2(new_n360), .A3(new_n402), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT34), .ZN(new_n448));
  INV_X1    g247(.A(G227gat), .ZN(new_n449));
  INV_X1    g248(.A(G233gat), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n447), .A2(new_n448), .A3(new_n452), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n336), .A2(new_n360), .A3(new_n402), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n402), .B1(new_n336), .B2(new_n360), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT34), .B1(new_n456), .B2(new_n451), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT33), .B1(new_n456), .B2(new_n451), .ZN(new_n458));
  XNOR2_X1  g257(.A(G15gat), .B(G43gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(G71gat), .B(G99gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n453), .B(new_n457), .C1(new_n458), .C2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n451), .A3(new_n446), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT32), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n461), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n448), .B1(new_n447), .B2(new_n452), .ZN(new_n468));
  AOI211_X1 g267(.A(KEYINPUT34), .B(new_n451), .C1(new_n445), .C2(new_n446), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n462), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n465), .B1(new_n462), .B2(new_n470), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n305), .A2(new_n444), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT35), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT91), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n435), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g276(.A(KEYINPUT91), .B(new_n425), .C1(new_n420), .C2(new_n429), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(new_n431), .A3(new_n433), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n443), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT94), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n471), .B2(new_n472), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n462), .A2(new_n470), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n464), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n462), .A2(new_n470), .A3(new_n465), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(KEYINPUT94), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT35), .B1(new_n377), .B2(new_n378), .ZN(new_n487));
  AND4_X1   g286(.A1(new_n480), .A2(new_n482), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n305), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n475), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n477), .A2(new_n478), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n428), .A2(new_n417), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(KEYINPUT89), .A3(new_n408), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n407), .B1(new_n426), .B2(new_n427), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(new_n404), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT39), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n403), .B2(new_n404), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n494), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n500), .A2(KEYINPUT40), .A3(new_n424), .A4(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n492), .A2(new_n378), .A3(new_n377), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n500), .A2(new_n424), .A3(new_n502), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT40), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n505), .A2(KEYINPUT90), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT90), .B1(new_n505), .B2(new_n506), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n491), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n479), .A2(new_n443), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n374), .B1(new_n370), .B2(KEYINPUT37), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT37), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(new_n367), .B2(new_n369), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT38), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT93), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n517), .B(KEYINPUT38), .C1(new_n512), .C2(new_n514), .ZN(new_n518));
  INV_X1    g317(.A(new_n512), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n368), .A2(new_n363), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n365), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n513), .B1(new_n521), .B2(new_n245), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n238), .B1(new_n365), .B2(new_n366), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT38), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n370), .ZN(new_n525));
  AOI22_X1  g324(.A1(new_n519), .A2(new_n524), .B1(new_n525), .B2(new_n373), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n511), .A2(new_n516), .A3(new_n518), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n503), .A2(new_n477), .A3(new_n478), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n379), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n508), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n505), .A2(KEYINPUT90), .A3(new_n506), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n532), .A3(KEYINPUT92), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n305), .A2(new_n510), .A3(new_n527), .A4(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n471), .B2(new_n472), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n484), .A2(KEYINPUT36), .A3(new_n485), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n299), .A2(new_n300), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n302), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n299), .A2(KEYINPUT87), .A3(new_n300), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n294), .A2(KEYINPUT88), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n540), .A2(new_n541), .B1(new_n542), .B2(new_n297), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n442), .A2(new_n443), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n379), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n538), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n534), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n490), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G57gat), .B(G64gat), .Z(new_n549));
  INV_X1    g348(.A(KEYINPUT9), .ZN(new_n550));
  INV_X1    g349(.A(G71gat), .ZN(new_n551));
  INV_X1    g350(.A(G78gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G71gat), .B(G78gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n549), .A2(new_n555), .A3(new_n553), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT21), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XOR2_X1   g363(.A(G127gat), .B(G155gat), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT20), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n564), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G183gat), .B(G211gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G15gat), .B(G22gat), .ZN(new_n570));
  INV_X1    g369(.A(G1gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(KEYINPUT16), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n571), .B2(new_n570), .ZN(new_n573));
  INV_X1    g372(.A(G8gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT98), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(KEYINPUT98), .A3(new_n574), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n570), .A2(new_n571), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n579), .A2(G8gat), .A3(new_n572), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(KEYINPUT97), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT97), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n579), .A2(new_n582), .A3(G8gat), .A4(new_n572), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n577), .A2(new_n578), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n561), .B2(new_n560), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT101), .B(KEYINPUT19), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n569), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n587), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  INV_X1    g391(.A(G92gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(new_n592), .B2(new_n593), .ZN(new_n596));
  NAND3_X1  g395(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G99gat), .B(G106gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n598), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT95), .B(G36gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(G29gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(G29gat), .A2(G36gat), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n604), .A2(KEYINPUT14), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(KEYINPUT14), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n603), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G43gat), .B(G50gat), .Z(new_n608));
  INV_X1    g407(.A(KEYINPUT15), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n607), .B(new_n610), .C1(KEYINPUT96), .C2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n610), .A2(new_n603), .A3(new_n605), .A4(new_n606), .ZN(new_n613));
  INV_X1    g412(.A(new_n611), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n603), .A2(KEYINPUT96), .A3(new_n605), .A4(new_n606), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n612), .A2(KEYINPUT17), .A3(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT17), .B1(new_n612), .B2(new_n616), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n601), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT103), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n598), .B(new_n599), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n612), .A2(new_n616), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(KEYINPUT102), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT102), .B1(new_n624), .B2(new_n625), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n620), .B(new_n622), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n621), .A2(KEYINPUT103), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n626), .ZN(new_n633));
  INV_X1    g432(.A(new_n630), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n622), .A4(new_n620), .ZN(new_n635));
  XNOR2_X1  g434(.A(G134gat), .B(G162gat), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n631), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n638), .B1(new_n631), .B2(new_n635), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n590), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n612), .A2(new_n616), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT17), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(new_n617), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n581), .A2(new_n583), .ZN(new_n648));
  INV_X1    g447(.A(new_n578), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT98), .B1(new_n573), .B2(new_n574), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n584), .A2(KEYINPUT99), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n647), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(G229gat), .A2(G233gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n644), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n655), .A2(KEYINPUT18), .A3(new_n656), .A4(new_n658), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT100), .B1(new_n584), .B2(new_n644), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(new_n658), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n656), .B(KEYINPUT13), .Z(new_n665));
  NAND3_X1  g464(.A1(new_n651), .A2(new_n657), .A3(KEYINPUT100), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n661), .A2(new_n662), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G113gat), .B(G141gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G197gat), .ZN(new_n670));
  XOR2_X1   g469(.A(KEYINPUT11), .B(G169gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT12), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n668), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n661), .A2(new_n675), .A3(new_n662), .A4(new_n667), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G230gat), .A2(G233gat), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n600), .A2(KEYINPUT104), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n559), .A2(new_n623), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT10), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n557), .A2(new_n558), .A3(new_n681), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n601), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n559), .A2(new_n623), .A3(KEYINPUT10), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n680), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n679), .B1(new_n682), .B2(new_n685), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(G120gat), .B(G148gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(G176gat), .B(G204gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n691), .B(new_n692), .Z(new_n693));
  AOI21_X1  g492(.A(KEYINPUT105), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695));
  INV_X1    g494(.A(new_n693), .ZN(new_n696));
  NOR4_X1   g495(.A1(new_n688), .A2(new_n695), .A3(new_n689), .A4(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n690), .A2(new_n693), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n643), .A2(new_n678), .A3(new_n702), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n548), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n544), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n380), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G8gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT106), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT16), .B(G8gat), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n708), .A2(KEYINPUT42), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT42), .B1(new_n708), .B2(new_n711), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n710), .A2(new_n714), .ZN(G1325gat));
  INV_X1    g514(.A(new_n704), .ZN(new_n716));
  INV_X1    g515(.A(new_n538), .ZN(new_n717));
  OAI21_X1  g516(.A(G15gat), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n482), .A2(new_n486), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OR2_X1    g519(.A1(new_n720), .A2(G15gat), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n718), .B1(new_n716), .B2(new_n721), .ZN(G1326gat));
  NAND2_X1  g521(.A1(new_n704), .A2(new_n543), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT43), .B(G22gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1327gat));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n475), .A2(new_n489), .B1(new_n534), .B2(new_n546), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(new_n642), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n534), .A2(new_n546), .ZN(new_n729));
  AOI22_X1  g528(.A1(new_n474), .A2(KEYINPUT35), .B1(new_n305), .B2(new_n488), .ZN(new_n730));
  OAI211_X1 g529(.A(KEYINPUT44), .B(new_n641), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n590), .A2(new_n678), .A3(new_n702), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n728), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G29gat), .B1(new_n733), .B2(new_n544), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n548), .A2(new_n641), .A3(new_n732), .ZN(new_n736));
  INV_X1    g535(.A(G29gat), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n705), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n736), .A2(new_n735), .A3(new_n738), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n734), .A2(new_n739), .A3(new_n740), .ZN(G1328gat));
  OAI21_X1  g540(.A(new_n602), .B1(new_n733), .B2(new_n379), .ZN(new_n742));
  INV_X1    g541(.A(new_n602), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n380), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT46), .B1(new_n736), .B2(new_n744), .ZN(new_n745));
  OR3_X1    g544(.A1(new_n736), .A2(KEYINPUT46), .A3(new_n744), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n742), .A2(new_n745), .A3(new_n746), .ZN(G1329gat));
  OAI21_X1  g546(.A(G43gat), .B1(new_n733), .B2(new_n717), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n720), .A2(G43gat), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(KEYINPUT107), .B1(new_n736), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n727), .A2(new_n642), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n752), .A2(new_n753), .A3(new_n732), .A4(new_n749), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n748), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n748), .A2(new_n755), .A3(KEYINPUT47), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(G1330gat));
  NAND4_X1  g559(.A1(new_n728), .A2(new_n543), .A3(new_n731), .A4(new_n732), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT108), .B1(new_n761), .B2(G50gat), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n305), .A2(G50gat), .ZN(new_n763));
  AND4_X1   g562(.A1(new_n548), .A2(new_n641), .A3(new_n732), .A4(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n761), .B2(G50gat), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT48), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n762), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI221_X4 g566(.A(new_n764), .B1(KEYINPUT108), .B2(KEYINPUT48), .C1(new_n761), .C2(G50gat), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n767), .A2(new_n768), .ZN(G1331gat));
  INV_X1    g568(.A(new_n702), .ZN(new_n770));
  NOR4_X1   g569(.A1(new_n727), .A2(new_n677), .A3(new_n643), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n705), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g572(.A(new_n379), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT109), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n771), .A2(new_n777), .A3(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1333gat));
  NAND2_X1  g580(.A1(new_n771), .A2(new_n538), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G71gat), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n771), .A2(new_n551), .A3(new_n719), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n785), .B(new_n786), .ZN(G1334gat));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n543), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(G78gat), .ZN(G1335gat));
  INV_X1    g588(.A(new_n590), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n678), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT110), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n792), .A2(new_n702), .ZN(new_n793));
  AND4_X1   g592(.A1(new_n705), .A2(new_n728), .A3(new_n731), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n548), .A2(new_n641), .A3(new_n792), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT51), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n548), .A2(new_n797), .A3(new_n641), .A4(new_n792), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n705), .A2(new_n592), .A3(new_n702), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n794), .A2(new_n592), .B1(new_n799), .B2(new_n800), .ZN(G1336gat));
  NAND4_X1  g600(.A1(new_n728), .A2(new_n793), .A3(new_n731), .A4(new_n380), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G92gat), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n770), .A2(new_n379), .A3(G92gat), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n796), .A2(new_n798), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n795), .A2(new_n808), .A3(new_n797), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n797), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n752), .A2(new_n792), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n812), .A2(new_n804), .B1(G92gat), .B2(new_n802), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n807), .B1(new_n813), .B2(new_n806), .ZN(G1337gat));
  NOR2_X1   g613(.A1(new_n720), .A2(G99gat), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n796), .A2(new_n702), .A3(new_n798), .A4(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n728), .A2(new_n793), .A3(new_n731), .A4(new_n538), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT112), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G99gat), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n817), .A2(KEYINPUT112), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n816), .B1(new_n819), .B2(new_n820), .ZN(G1338gat));
  NOR2_X1   g620(.A1(new_n305), .A2(G106gat), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n796), .A2(new_n702), .A3(new_n798), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT113), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n728), .A2(new_n793), .A3(new_n731), .A4(new_n543), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT53), .B1(new_n825), .B2(G106gat), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n823), .A2(KEYINPUT113), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n305), .A2(G106gat), .A3(new_n770), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n812), .A2(new_n830), .B1(G106gat), .B2(new_n825), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n827), .A2(new_n828), .B1(new_n829), .B2(new_n831), .ZN(G1339gat));
  NAND2_X1  g631(.A1(new_n686), .A2(new_n687), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n679), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n686), .A2(new_n680), .A3(new_n687), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(KEYINPUT54), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n693), .B1(new_n688), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(KEYINPUT55), .A3(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n840));
  OAI211_X1 g639(.A(new_n839), .B(new_n840), .C1(new_n694), .C2(new_n697), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n839), .B1(new_n694), .B2(new_n697), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT114), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n836), .A2(new_n838), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n677), .A2(new_n841), .A3(new_n843), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n664), .A2(new_n666), .ZN(new_n848));
  INV_X1    g647(.A(new_n665), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n656), .B1(new_n655), .B2(new_n658), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n672), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n702), .A2(new_n855), .A3(new_n676), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n641), .B1(new_n847), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n641), .A2(new_n855), .A3(new_n676), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n843), .A2(new_n841), .A3(new_n846), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n790), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n590), .A2(new_n678), .A3(new_n642), .A4(new_n770), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n861), .A2(KEYINPUT116), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT116), .B1(new_n861), .B2(new_n862), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n305), .A2(new_n379), .A3(new_n473), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n865), .A2(new_n705), .A3(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(G113gat), .B1(new_n868), .B2(new_n677), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n544), .A2(new_n380), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n865), .A2(new_n305), .A3(new_n719), .A4(new_n870), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n871), .A2(new_n383), .A3(new_n678), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n869), .A2(new_n872), .ZN(G1340gat));
  OAI21_X1  g672(.A(G120gat), .B1(new_n871), .B2(new_n770), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n702), .A2(new_n400), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT117), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n874), .B1(new_n867), .B2(new_n876), .ZN(G1341gat));
  OAI21_X1  g676(.A(G127gat), .B1(new_n871), .B2(new_n790), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n790), .A2(G127gat), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n878), .B1(new_n867), .B2(new_n879), .ZN(G1342gat));
  OAI21_X1  g679(.A(G134gat), .B1(new_n871), .B2(new_n642), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT56), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n642), .A2(G134gat), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n867), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n884), .A2(KEYINPUT118), .A3(new_n882), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT118), .B1(new_n884), .B2(new_n882), .ZN(new_n886));
  OAI221_X1 g685(.A(new_n881), .B1(new_n882), .B2(new_n884), .C1(new_n885), .C2(new_n886), .ZN(G1343gat));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT55), .B1(new_n844), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n888), .B2(new_n844), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n677), .A2(new_n699), .A3(new_n839), .A4(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n641), .B1(new_n891), .B2(new_n856), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n790), .B1(new_n892), .B2(new_n860), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n862), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n305), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n856), .B1(new_n678), .B2(new_n859), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n860), .B1(new_n899), .B2(new_n642), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n862), .B1(new_n900), .B2(new_n590), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n861), .A2(KEYINPUT116), .A3(new_n862), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n543), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n898), .B1(new_n905), .B2(new_n895), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n717), .A2(new_n870), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n906), .A2(new_n678), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(new_n212), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n903), .A2(new_n904), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n544), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n717), .A2(new_n543), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(new_n380), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n677), .A2(new_n212), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT58), .B1(new_n909), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  OAI221_X1 g717(.A(new_n918), .B1(new_n914), .B2(new_n915), .C1(new_n908), .C2(new_n212), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1344gat));
  NOR3_X1   g719(.A1(new_n906), .A2(new_n770), .A3(new_n907), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n214), .A2(KEYINPUT59), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT121), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n907), .ZN(new_n925));
  AOI21_X1  g724(.A(KEYINPUT57), .B1(new_n865), .B2(new_n543), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n702), .B(new_n925), .C1(new_n926), .C2(new_n898), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n928), .A3(new_n922), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT57), .B1(new_n894), .B2(new_n543), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n903), .A2(new_n904), .A3(new_n896), .ZN(new_n932));
  AOI211_X1 g731(.A(new_n770), .B(new_n907), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT59), .B1(new_n933), .B2(new_n214), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n924), .A2(new_n929), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n770), .A2(G148gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n911), .A2(new_n913), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT120), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n935), .A2(new_n938), .ZN(G1345gat));
  NOR3_X1   g738(.A1(new_n906), .A2(new_n790), .A3(new_n907), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n590), .A2(new_n206), .ZN(new_n941));
  OAI22_X1  g740(.A1(new_n940), .A2(new_n206), .B1(new_n914), .B2(new_n941), .ZN(G1346gat));
  NOR2_X1   g741(.A1(new_n906), .A2(new_n907), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n642), .A2(new_n207), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n911), .A2(new_n641), .A3(new_n913), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n943), .A2(new_n944), .B1(new_n945), .B2(new_n207), .ZN(G1347gat));
  NAND2_X1  g745(.A1(new_n544), .A2(new_n380), .ZN(new_n947));
  XOR2_X1   g746(.A(new_n947), .B(KEYINPUT123), .Z(new_n948));
  NAND4_X1  g747(.A1(new_n865), .A2(new_n305), .A3(new_n719), .A4(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(G169gat), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n949), .A2(new_n950), .A3(new_n678), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n910), .A2(new_n705), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n305), .A2(new_n380), .A3(new_n473), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT122), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n952), .A2(new_n677), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n951), .B1(new_n950), .B2(new_n955), .ZN(G1348gat));
  OAI21_X1  g755(.A(G176gat), .B1(new_n949), .B2(new_n770), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n952), .A2(new_n954), .ZN(new_n958));
  OR2_X1    g757(.A1(new_n770), .A2(G176gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT124), .ZN(G1349gat));
  OAI21_X1  g760(.A(G183gat), .B1(new_n949), .B2(new_n790), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT60), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n952), .A2(new_n334), .A3(new_n590), .A4(new_n954), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n962), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OR2_X1    g765(.A1(new_n963), .A2(KEYINPUT60), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n966), .B(new_n967), .ZN(G1350gat));
  OAI21_X1  g767(.A(G190gat), .B1(new_n949), .B2(new_n642), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT61), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n641), .A2(new_n318), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n958), .B2(new_n971), .ZN(G1351gat));
  NAND2_X1  g771(.A1(new_n948), .A2(new_n717), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n931), .A2(new_n932), .ZN(new_n976));
  NAND4_X1  g775(.A1(new_n975), .A2(G197gat), .A3(new_n677), .A4(new_n976), .ZN(new_n977));
  INV_X1    g776(.A(G197gat), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n912), .A2(new_n379), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n952), .A2(new_n979), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n978), .B1(new_n980), .B2(new_n678), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(KEYINPUT127), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n977), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n983), .A2(new_n985), .ZN(G1352gat));
  INV_X1    g785(.A(G204gat), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n702), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g787(.A(KEYINPUT62), .B1(new_n980), .B2(new_n988), .ZN(new_n989));
  OR3_X1    g788(.A1(new_n980), .A2(KEYINPUT62), .A3(new_n988), .ZN(new_n990));
  INV_X1    g789(.A(new_n975), .ZN(new_n991));
  INV_X1    g790(.A(new_n976), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n991), .A2(new_n770), .A3(new_n992), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n989), .B(new_n990), .C1(new_n993), .C2(new_n987), .ZN(G1353gat));
  AOI211_X1 g793(.A(new_n790), .B(new_n973), .C1(new_n931), .C2(new_n932), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n995), .A2(new_n226), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n996), .A2(KEYINPUT63), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT63), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n995), .A2(new_n998), .A3(new_n226), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n590), .A2(new_n242), .ZN(new_n1000));
  OAI22_X1  g799(.A1(new_n997), .A2(new_n999), .B1(new_n980), .B2(new_n1000), .ZN(G1354gat));
  NOR2_X1   g800(.A1(new_n991), .A2(new_n992), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n642), .A2(new_n235), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n952), .A2(new_n641), .A3(new_n979), .ZN(new_n1004));
  AOI22_X1  g803(.A1(new_n1002), .A2(new_n1003), .B1(new_n235), .B2(new_n1004), .ZN(G1355gat));
endmodule


