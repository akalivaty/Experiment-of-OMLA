//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G141gat), .B(G148gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT78), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT2), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n205), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(new_n206), .B2(new_n209), .ZN(new_n211));
  XNOR2_X1  g010(.A(G155gat), .B(G162gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT77), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n205), .B(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT80), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n218), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n217), .A2(new_n209), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n215), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT29), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(G211gat), .A2(G218gat), .ZN(new_n226));
  AND2_X1   g025(.A1(G197gat), .A2(G204gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(G197gat), .A2(G204gat), .ZN(new_n228));
  OAI22_X1  g027(.A1(KEYINPUT22), .A2(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(G211gat), .B(G218gat), .Z(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(KEYINPUT74), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n229), .A2(new_n230), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(new_n231), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT74), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n225), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n215), .A2(new_n221), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT29), .B1(new_n234), .B2(new_n231), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(KEYINPUT3), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n204), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n204), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n244), .B1(new_n225), .B2(new_n237), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT83), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n222), .B1(new_n237), .B2(KEYINPUT29), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n239), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n245), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n246), .B1(new_n245), .B2(new_n248), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n243), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(G22gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(G78gat), .B(G106gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT31), .B(G50gat), .ZN(new_n254));
  XOR2_X1   g053(.A(new_n253), .B(new_n254), .Z(new_n255));
  NOR2_X1   g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n245), .A2(new_n248), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT83), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n245), .A2(new_n246), .A3(new_n248), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n242), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(G22gat), .B1(new_n260), .B2(KEYINPUT84), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT84), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n251), .A2(new_n262), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n261), .A2(new_n263), .A3(KEYINPUT85), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT85), .ZN(new_n265));
  INV_X1    g064(.A(G22gat), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n266), .B1(new_n251), .B2(new_n262), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n260), .A2(KEYINPUT84), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n265), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n256), .B1(new_n264), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n251), .B(new_n266), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n255), .B(KEYINPUT82), .Z(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT27), .B(G183gat), .ZN(new_n276));
  INV_X1    g075(.A(G190gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT28), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT26), .ZN(new_n283));
  NOR2_X1   g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n284), .A2(KEYINPUT67), .A3(new_n283), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT67), .B1(new_n284), .B2(new_n283), .ZN(new_n286));
  OAI221_X1 g085(.A(new_n282), .B1(new_n283), .B2(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n280), .A2(new_n281), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT68), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n280), .A2(KEYINPUT68), .A3(new_n281), .A4(new_n287), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(G183gat), .B2(G190gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT65), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT24), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n296), .A2(new_n297), .B1(G183gat), .B2(G190gat), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n294), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n282), .A2(KEYINPUT23), .ZN(new_n300));
  INV_X1    g099(.A(G169gat), .ZN(new_n301));
  INV_X1    g100(.A(G176gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n284), .A2(KEYINPUT23), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(KEYINPUT25), .A3(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n305), .B(KEYINPUT64), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n304), .B1(new_n294), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n310), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n309), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n292), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G113gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(G120gat), .ZN(new_n318));
  OR2_X1    g117(.A1(new_n318), .A2(KEYINPUT70), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(KEYINPUT70), .ZN(new_n320));
  INV_X1    g119(.A(G120gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n319), .B(new_n320), .C1(G113gat), .C2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323));
  XNOR2_X1  g122(.A(G127gat), .B(G134gat), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT69), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n324), .B(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n321), .A2(G113gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n323), .B1(new_n318), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n331), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n290), .A2(new_n291), .B1(new_n309), .B2(new_n314), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n325), .A2(new_n330), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G227gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n332), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT32), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n338), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n342));
  XNOR2_X1  g141(.A(G15gat), .B(G43gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(G71gat), .B(G99gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT33), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n345), .B1(new_n338), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n342), .A3(new_n347), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n338), .B(KEYINPUT32), .C1(new_n346), .C2(new_n345), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT72), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT34), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n332), .A2(new_n335), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(new_n336), .ZN(new_n354));
  AOI211_X1 g153(.A(KEYINPUT34), .B(new_n337), .C1(new_n332), .C2(new_n335), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n356), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n350), .A2(KEYINPUT72), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n275), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n239), .A2(new_n334), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n239), .A2(new_n334), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT5), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n239), .A2(KEYINPUT3), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n366), .A2(new_n223), .A3(new_n334), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(KEYINPUT4), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n239), .B2(new_n334), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n367), .A2(new_n368), .A3(new_n364), .A4(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n368), .A2(new_n370), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n373), .A2(KEYINPUT5), .A3(new_n364), .A4(new_n367), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(KEYINPUT0), .ZN(new_n377));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n377), .B(new_n378), .Z(new_n379));
  NAND2_X1  g178(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT6), .ZN(new_n381));
  INV_X1    g180(.A(new_n379), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n372), .A2(new_n374), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT81), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n380), .A2(new_n386), .A3(new_n381), .A4(new_n383), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n383), .A2(new_n381), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(new_n333), .B2(KEYINPUT29), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT75), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT75), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n393), .B(new_n390), .C1(new_n333), .C2(KEYINPUT29), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n315), .A2(new_n288), .ZN(new_n395));
  INV_X1    g194(.A(new_n390), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n392), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(new_n237), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n224), .A3(new_n390), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n333), .A2(new_n396), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n237), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G8gat), .B(G36gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(G64gat), .B(G92gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n405), .B(new_n406), .Z(new_n407));
  NAND3_X1  g206(.A1(new_n399), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(KEYINPUT76), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n407), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n391), .A2(KEYINPUT75), .B1(new_n396), .B2(new_n395), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n403), .B1(new_n412), .B2(new_n394), .ZN(new_n413));
  INV_X1    g212(.A(new_n404), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n413), .A2(new_n414), .A3(new_n411), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT76), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT30), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n389), .A2(new_n410), .A3(new_n415), .A4(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT35), .B1(new_n360), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT73), .B1(new_n350), .B2(new_n358), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n350), .A2(new_n358), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT73), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n348), .A2(new_n356), .A3(new_n349), .A4(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT85), .B1(new_n261), .B2(new_n263), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n267), .A2(new_n265), .A3(new_n268), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n273), .B1(new_n428), .B2(new_n256), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n418), .A2(new_n410), .A3(new_n415), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT35), .B1(new_n384), .B2(new_n388), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n420), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n373), .A2(new_n367), .ZN(new_n436));
  INV_X1    g235(.A(new_n364), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n363), .A2(new_n364), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(KEYINPUT39), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT39), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n436), .A2(new_n441), .A3(new_n437), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n379), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT40), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n440), .A2(KEYINPUT40), .A3(new_n379), .A4(new_n442), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n445), .A2(new_n383), .A3(new_n446), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n431), .A2(new_n447), .B1(new_n270), .B2(new_n274), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n411), .A2(KEYINPUT37), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n399), .A2(new_n404), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n415), .A2(new_n450), .B1(new_n451), .B2(KEYINPUT37), .ZN(new_n452));
  XOR2_X1   g251(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n453));
  OAI21_X1  g252(.A(new_n449), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n384), .A2(new_n408), .A3(new_n388), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n415), .A2(new_n450), .ZN(new_n456));
  INV_X1    g255(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n398), .A2(new_n403), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT37), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n402), .B2(new_n237), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n457), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n455), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n411), .B1(new_n451), .B2(KEYINPUT37), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n459), .B1(new_n399), .B2(new_n404), .ZN(new_n464));
  OAI211_X1 g263(.A(KEYINPUT87), .B(new_n457), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n454), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n425), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n357), .A2(KEYINPUT36), .A3(new_n359), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n419), .A2(new_n429), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n467), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n435), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT88), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT88), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n435), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G29gat), .ZN(new_n478));
  OR2_X1    g277(.A1(KEYINPUT89), .A2(G36gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(KEYINPUT89), .A2(G36gat), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(G50gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G43gat), .ZN(new_n483));
  INV_X1    g282(.A(G43gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G50gat), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT90), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(G36gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n478), .A2(new_n487), .A3(KEYINPUT14), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT14), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(G29gat), .B2(G36gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n481), .A2(new_n486), .A3(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n484), .A2(G50gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n482), .A2(G43gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n488), .A2(new_n490), .ZN(new_n496));
  INV_X1    g295(.A(new_n480), .ZN(new_n497));
  NOR2_X1   g296(.A1(KEYINPUT89), .A2(G36gat), .ZN(new_n498));
  OAI21_X1  g297(.A(G29gat), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n495), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT15), .B1(new_n492), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT90), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(new_n493), .B2(new_n494), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n496), .A2(new_n504), .A3(new_n499), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT15), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n501), .A2(new_n502), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n483), .A2(new_n485), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(new_n481), .B2(new_n491), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n506), .B1(new_n505), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n481), .A2(new_n491), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT15), .B1(new_n512), .B2(new_n504), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT17), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT91), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G8gat), .ZN(new_n517));
  INV_X1    g316(.A(G8gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(KEYINPUT91), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  AOI21_X1  g320(.A(G1gat), .B1(new_n515), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n517), .A2(new_n522), .A3(new_n519), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n514), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n528), .B(KEYINPUT92), .Z(new_n529));
  NOR2_X1   g328(.A1(new_n511), .A2(new_n513), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(new_n525), .A3(new_n524), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT18), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT94), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n532), .A2(KEYINPUT94), .A3(new_n533), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n527), .A2(KEYINPUT18), .A3(new_n529), .A4(new_n531), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT93), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n529), .B(KEYINPUT13), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n526), .B1(new_n511), .B2(new_n513), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(new_n531), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(new_n539), .B2(new_n540), .ZN(new_n545));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(G197gat), .ZN(new_n547));
  XOR2_X1   g346(.A(KEYINPUT11), .B(G169gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT12), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n538), .A2(new_n541), .A3(new_n545), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n541), .A2(new_n545), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n552), .B1(new_n533), .B2(new_n532), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n551), .B1(new_n553), .B2(new_n550), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n475), .A2(new_n477), .A3(new_n554), .ZN(new_n555));
  AND2_X1   g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G57gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(G64gat), .ZN(new_n563));
  INV_X1    g362(.A(G64gat), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(G57gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G71gat), .B(G78gat), .ZN(new_n567));
  INV_X1    g366(.A(new_n560), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(G231gat), .A2(G233gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(G127gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n526), .B1(new_n571), .B2(new_n570), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(new_n207), .ZN(new_n579));
  XOR2_X1   g378(.A(G183gat), .B(G211gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n577), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n577), .A2(new_n582), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT8), .ZN(new_n590));
  OR2_X1    g389(.A1(G85gat), .A2(G92gat), .ZN(new_n591));
  NAND4_X1  g390(.A1(KEYINPUT95), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n588), .A2(new_n590), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT96), .ZN(new_n594));
  OR2_X1    g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n589), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n594), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n588), .A2(new_n592), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n590), .A2(new_n591), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n595), .A2(KEYINPUT96), .A3(new_n589), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n508), .A2(new_n514), .A3(new_n597), .A4(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n597), .ZN(new_n604));
  AND2_X1   g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n530), .A2(new_n604), .B1(KEYINPUT41), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G190gat), .B(G218gat), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n607), .B(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n611));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n610), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n585), .A2(new_n614), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n561), .A2(new_n569), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n593), .A2(KEYINPUT97), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n596), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n593), .A2(KEYINPUT97), .A3(new_n589), .A4(new_n595), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT10), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n602), .A2(new_n570), .A3(new_n597), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n616), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(new_n620), .B2(new_n622), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n628), .A2(KEYINPUT98), .ZN(new_n629));
  XNOR2_X1  g428(.A(G120gat), .B(G148gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(G176gat), .B(G204gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n630), .B(new_n631), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(KEYINPUT98), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n627), .A2(new_n629), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n626), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n623), .B2(new_n624), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(new_n628), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n632), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT99), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT99), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n634), .B(new_n641), .C1(new_n638), .C2(new_n632), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n615), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n555), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n389), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g446(.A1(new_n645), .A2(new_n432), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT16), .B(G8gat), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n650), .B1(new_n518), .B2(new_n648), .ZN(new_n651));
  MUX2_X1   g450(.A(new_n650), .B(new_n651), .S(KEYINPUT42), .Z(G1325gat));
  AND2_X1   g451(.A1(new_n422), .A2(new_n424), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT36), .B1(new_n653), .B2(new_n421), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n357), .A2(KEYINPUT36), .A3(new_n359), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT100), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n469), .A2(new_n657), .A3(new_n470), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(G15gat), .B1(new_n645), .B2(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n425), .A2(G15gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n645), .B2(new_n661), .ZN(G1326gat));
  OR3_X1    g461(.A1(new_n645), .A2(KEYINPUT101), .A3(new_n275), .ZN(new_n663));
  OAI21_X1  g462(.A(KEYINPUT101), .B1(new_n645), .B2(new_n275), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT43), .B(G22gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1327gat));
  NOR3_X1   g466(.A1(new_n585), .A2(new_n614), .A3(new_n643), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n555), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n389), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(new_n478), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT45), .ZN(new_n673));
  INV_X1    g472(.A(new_n614), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n475), .A2(KEYINPUT44), .A3(new_n477), .A4(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676));
  AOI22_X1  g475(.A1(new_n448), .A2(new_n466), .B1(new_n419), .B2(new_n429), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n659), .A2(new_n677), .B1(new_n420), .B2(new_n434), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n678), .B2(new_n614), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n585), .ZN(new_n681));
  INV_X1    g480(.A(new_n643), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n680), .A2(new_n554), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(G29gat), .B1(new_n683), .B2(new_n389), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n673), .A2(new_n684), .ZN(G1328gat));
  NAND2_X1  g484(.A1(new_n479), .A2(new_n480), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n669), .A2(new_n432), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT46), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n686), .B1(new_n683), .B2(new_n432), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1329gat));
  OAI21_X1  g489(.A(new_n484), .B1(new_n669), .B2(new_n425), .ZN(new_n691));
  INV_X1    g490(.A(new_n659), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G43gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n683), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g494(.A1(new_n669), .A2(G50gat), .A3(new_n275), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT48), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(KEYINPUT102), .B2(new_n697), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n697), .A2(KEYINPUT102), .ZN(new_n699));
  OAI21_X1  g498(.A(G50gat), .B1(new_n683), .B2(new_n275), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(G1331gat));
  AND3_X1   g502(.A1(new_n469), .A2(new_n657), .A3(new_n470), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n657), .B1(new_n469), .B2(new_n470), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n677), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n435), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n615), .A2(new_n554), .A3(new_n682), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n389), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(new_n562), .ZN(G1332gat));
  XOR2_X1   g510(.A(new_n709), .B(KEYINPUT103), .Z(new_n712));
  OAI22_X1  g511(.A1(new_n712), .A2(new_n432), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  OR2_X1    g512(.A1(new_n712), .A2(new_n432), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT49), .B(G64gat), .Z(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT104), .ZN(G1333gat));
  NAND2_X1  g516(.A1(new_n692), .A2(G71gat), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n709), .A2(new_n425), .ZN(new_n719));
  OAI22_X1  g518(.A1(new_n712), .A2(new_n718), .B1(G71gat), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1334gat));
  NOR2_X1   g521(.A1(new_n712), .A2(new_n275), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT106), .B(G78gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1335gat));
  NOR2_X1   g524(.A1(new_n554), .A2(new_n585), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n707), .A2(new_n674), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT51), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g528(.A1(new_n707), .A2(KEYINPUT51), .A3(new_n674), .A4(new_n726), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n729), .A2(KEYINPUT107), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n727), .A2(new_n732), .A3(new_n728), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR4_X1   g533(.A1(new_n734), .A2(G85gat), .A3(new_n389), .A4(new_n682), .ZN(new_n735));
  INV_X1    g534(.A(G85gat), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n554), .A2(new_n585), .A3(new_n682), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n680), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(new_n671), .ZN(new_n739));
  OR2_X1    g538(.A1(new_n735), .A2(new_n739), .ZN(G1336gat));
  NAND4_X1  g539(.A1(new_n675), .A2(new_n679), .A3(new_n431), .A4(new_n737), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n741), .A2(G92gat), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n432), .A2(G92gat), .A3(new_n682), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT108), .Z(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n729), .B2(new_n730), .ZN(new_n745));
  OAI21_X1  g544(.A(KEYINPUT52), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT52), .B1(new_n741), .B2(G92gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n733), .A3(new_n743), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n749), .B1(new_n747), .B2(new_n748), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n746), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI211_X1 g553(.A(KEYINPUT110), .B(new_n746), .C1(new_n750), .C2(new_n751), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(G1337gat));
  NOR4_X1   g555(.A1(new_n734), .A2(G99gat), .A3(new_n425), .A4(new_n682), .ZN(new_n757));
  INV_X1    g556(.A(G99gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n738), .B2(new_n692), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n757), .A2(new_n759), .ZN(G1338gat));
  NAND2_X1  g559(.A1(new_n738), .A2(new_n429), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G106gat), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n275), .A2(G106gat), .A3(new_n682), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n731), .A2(new_n733), .A3(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n729), .A2(new_n730), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n761), .A2(G106gat), .B1(new_n767), .B2(new_n765), .ZN(new_n768));
  OAI22_X1  g567(.A1(new_n764), .A2(new_n766), .B1(new_n768), .B2(new_n763), .ZN(G1339gat));
  NAND3_X1  g568(.A1(new_n623), .A2(new_n636), .A3(new_n624), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n623), .A2(KEYINPUT111), .A3(new_n636), .A4(new_n624), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n772), .A2(new_n627), .A3(KEYINPUT54), .A4(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n632), .B1(new_n637), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(KEYINPUT55), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n614), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n774), .A2(KEYINPUT55), .A3(new_n776), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n774), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(new_n776), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT113), .B1(new_n784), .B2(new_n634), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  AOI211_X1 g585(.A(new_n786), .B(new_n635), .C1(new_n782), .C2(new_n783), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n779), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n543), .A2(new_n531), .A3(new_n542), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n529), .B1(new_n527), .B2(new_n531), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n549), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n551), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n532), .A2(KEYINPUT94), .A3(new_n533), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT94), .B1(new_n532), .B2(new_n533), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n550), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(KEYINPUT114), .B(new_n791), .C1(new_n797), .C2(new_n552), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT115), .B1(new_n788), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n634), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n786), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n635), .B1(new_n782), .B2(new_n783), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT113), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n806));
  AOI21_X1  g605(.A(KEYINPUT114), .B1(new_n551), .B2(new_n791), .ZN(new_n807));
  INV_X1    g606(.A(new_n798), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n805), .A2(new_n806), .A3(new_n779), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n800), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n643), .A2(new_n551), .A3(new_n791), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n785), .A2(new_n787), .ZN(new_n813));
  INV_X1    g612(.A(new_n778), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n554), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n614), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n585), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n554), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n644), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT116), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n800), .A2(new_n810), .B1(new_n816), .B2(new_n614), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n823), .B(new_n820), .C1(new_n824), .C2(new_n585), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(new_n671), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n827), .A2(new_n432), .A3(new_n430), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(new_n317), .A3(new_n819), .ZN(new_n829));
  INV_X1    g628(.A(new_n360), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n432), .A3(new_n830), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n831), .A2(new_n819), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n829), .B1(new_n317), .B2(new_n832), .ZN(G1340gat));
  OAI21_X1  g632(.A(G120gat), .B1(new_n828), .B2(new_n682), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n643), .A2(new_n321), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT117), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n834), .B1(new_n831), .B2(new_n836), .ZN(G1341gat));
  OAI21_X1  g636(.A(G127gat), .B1(new_n828), .B2(new_n681), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n681), .A2(G127gat), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n831), .B2(new_n839), .ZN(G1342gat));
  NOR3_X1   g639(.A1(new_n831), .A2(G134gat), .A3(new_n614), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT56), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT118), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n828), .B2(new_n614), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n844), .B(new_n845), .C1(new_n842), .C2(new_n841), .ZN(G1343gat));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n822), .A2(new_n429), .A3(new_n825), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n848), .A2(KEYINPUT119), .A3(new_n849), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n778), .B(KEYINPUT120), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n554), .A3(new_n803), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n812), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n614), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n811), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n681), .ZN(new_n859));
  AOI211_X1 g658(.A(new_n849), .B(new_n275), .C1(new_n859), .C2(new_n820), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n852), .A2(new_n853), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n659), .A2(new_n671), .A3(new_n432), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n862), .A2(new_n554), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(G141gat), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n847), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(G141gat), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n860), .B1(new_n850), .B2(new_n851), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n863), .B1(new_n870), .B2(new_n853), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n869), .B1(new_n871), .B2(new_n554), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n848), .A2(new_n863), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n819), .A2(G141gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT122), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n866), .A2(new_n878), .A3(new_n875), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n868), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  AOI211_X1 g679(.A(new_n819), .B(new_n863), .C1(new_n870), .C2(new_n853), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n867), .B1(new_n881), .B2(new_n869), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n877), .A2(new_n879), .B1(KEYINPUT58), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n880), .A2(new_n883), .ZN(G1344gat));
  INV_X1    g683(.A(G148gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n873), .A2(new_n885), .A3(new_n643), .ZN(new_n886));
  AOI211_X1 g685(.A(KEYINPUT59), .B(new_n885), .C1(new_n871), .C2(new_n643), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888));
  INV_X1    g687(.A(new_n788), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n799), .B1(new_n889), .B2(KEYINPUT123), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n890), .B1(KEYINPUT123), .B2(new_n889), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n585), .B1(new_n891), .B2(new_n857), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n821), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(KEYINPUT57), .A3(new_n275), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(KEYINPUT57), .B2(new_n848), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n895), .A2(new_n643), .A3(new_n864), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n888), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n886), .B1(new_n887), .B2(new_n897), .ZN(G1345gat));
  AOI21_X1  g697(.A(G155gat), .B1(new_n873), .B2(new_n585), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n585), .A2(G155gat), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n900), .B(KEYINPUT124), .Z(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n871), .B2(new_n901), .ZN(G1346gat));
  NAND3_X1  g701(.A1(new_n873), .A2(new_n208), .A3(new_n674), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n871), .A2(new_n674), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n208), .ZN(G1347gat));
  AND2_X1   g704(.A1(new_n826), .A2(new_n389), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n906), .A2(new_n431), .A3(new_n830), .ZN(new_n907));
  AOI21_X1  g706(.A(G169gat), .B1(new_n907), .B2(new_n554), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n431), .A3(new_n430), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(new_n301), .A3(new_n819), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n908), .A2(new_n910), .ZN(G1348gat));
  NAND3_X1  g710(.A1(new_n907), .A2(new_n302), .A3(new_n643), .ZN(new_n912));
  OAI21_X1  g711(.A(G176gat), .B1(new_n909), .B2(new_n682), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1349gat));
  NOR2_X1   g713(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n907), .A2(new_n276), .A3(new_n585), .ZN(new_n916));
  OAI21_X1  g715(.A(G183gat), .B1(new_n909), .B2(new_n681), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n919));
  XOR2_X1   g718(.A(new_n918), .B(new_n919), .Z(G1350gat));
  OAI21_X1  g719(.A(G190gat), .B1(new_n909), .B2(new_n614), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT61), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT61), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n923), .B(G190gat), .C1(new_n909), .C2(new_n614), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n907), .A2(new_n277), .A3(new_n674), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT126), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n929), .A3(new_n926), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1351gat));
  NOR3_X1   g730(.A1(new_n692), .A2(new_n671), .A3(new_n432), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n895), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(G197gat), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n933), .A2(new_n934), .A3(new_n819), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n692), .A2(new_n432), .A3(new_n275), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n906), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n554), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n935), .A2(new_n939), .ZN(G1352gat));
  NOR3_X1   g739(.A1(new_n937), .A2(G204gat), .A3(new_n682), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT62), .ZN(new_n942));
  OAI21_X1  g741(.A(G204gat), .B1(new_n933), .B2(new_n682), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1353gat));
  INV_X1    g743(.A(G211gat), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n938), .A2(new_n945), .A3(new_n585), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n895), .A2(new_n585), .A3(new_n932), .ZN(new_n948));
  AND4_X1   g747(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n945), .B1(KEYINPUT127), .B2(new_n950), .ZN(new_n951));
  AOI22_X1  g750(.A1(new_n948), .A2(new_n951), .B1(new_n947), .B2(KEYINPUT63), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n946), .B1(new_n949), .B2(new_n952), .ZN(G1354gat));
  OAI21_X1  g752(.A(G218gat), .B1(new_n933), .B2(new_n614), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n614), .A2(G218gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n937), .B2(new_n955), .ZN(G1355gat));
endmodule


