

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(n722), .ZN(n737) );
  AND2_X1 U553 ( .A1(n818), .A2(n817), .ZN(n518) );
  NOR2_X1 U554 ( .A1(n662), .A2(n529), .ZN(n519) );
  XOR2_X1 U555 ( .A(KEYINPUT76), .B(n607), .Z(n520) );
  NOR2_X1 U556 ( .A1(G168), .A2(n700), .ZN(n701) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n732) );
  XNOR2_X1 U558 ( .A(n733), .B(n732), .ZN(n736) );
  NAND2_X1 U559 ( .A1(n736), .A2(n735), .ZN(n753) );
  INV_X1 U560 ( .A(KEYINPUT99), .ZN(n760) );
  XNOR2_X1 U561 ( .A(n761), .B(n760), .ZN(n777) );
  AND2_X1 U562 ( .A1(n772), .A2(n1006), .ZN(n773) );
  NOR2_X1 U563 ( .A1(G164), .A2(G1384), .ZN(n694) );
  NAND2_X1 U564 ( .A1(n774), .A2(n773), .ZN(n775) );
  INV_X1 U565 ( .A(G543), .ZN(n523) );
  NOR2_X1 U566 ( .A1(G651), .A2(G543), .ZN(n648) );
  XOR2_X1 U567 ( .A(KEYINPUT77), .B(n612), .Z(n997) );
  XNOR2_X1 U568 ( .A(n523), .B(KEYINPUT0), .ZN(n662) );
  NOR2_X1 U569 ( .A1(n556), .A2(n555), .ZN(G160) );
  INV_X1 U570 ( .A(G651), .ZN(n529) );
  NOR2_X1 U571 ( .A1(G543), .A2(n529), .ZN(n521) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n521), .Z(n661) );
  NAND2_X1 U573 ( .A1(n661), .A2(G63), .ZN(n522) );
  XOR2_X1 U574 ( .A(KEYINPUT79), .B(n522), .Z(n526) );
  NOR2_X1 U575 ( .A1(G651), .A2(n662), .ZN(n524) );
  XNOR2_X1 U576 ( .A(KEYINPUT66), .B(n524), .ZN(n656) );
  NAND2_X1 U577 ( .A1(G51), .A2(n656), .ZN(n525) );
  NAND2_X1 U578 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U579 ( .A(KEYINPUT6), .B(n527), .ZN(n535) );
  NAND2_X1 U580 ( .A1(n648), .A2(G89), .ZN(n528) );
  XNOR2_X1 U581 ( .A(n528), .B(KEYINPUT4), .ZN(n531) );
  NAND2_X1 U582 ( .A1(G76), .A2(n519), .ZN(n530) );
  NAND2_X1 U583 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U584 ( .A(KEYINPUT5), .B(n532), .Z(n533) );
  XNOR2_X1 U585 ( .A(KEYINPUT78), .B(n533), .ZN(n534) );
  NOR2_X1 U586 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U587 ( .A(n536), .B(KEYINPUT7), .Z(n537) );
  XNOR2_X1 U588 ( .A(KEYINPUT80), .B(n537), .ZN(G168) );
  INV_X1 U589 ( .A(G2104), .ZN(n538) );
  NOR2_X4 U590 ( .A1(G2105), .A2(n538), .ZN(n901) );
  NAND2_X1 U591 ( .A1(G102), .A2(n901), .ZN(n541) );
  NOR2_X1 U592 ( .A1(G2104), .A2(G2105), .ZN(n539) );
  XOR2_X2 U593 ( .A(KEYINPUT17), .B(n539), .Z(n902) );
  NAND2_X1 U594 ( .A1(G138), .A2(n902), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n548) );
  NAND2_X1 U596 ( .A1(G2105), .A2(G2104), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n542), .B(KEYINPUT69), .ZN(n907) );
  NAND2_X1 U598 ( .A1(G114), .A2(n907), .ZN(n546) );
  INV_X1 U599 ( .A(G2104), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n543), .A2(G2105), .ZN(n544) );
  XNOR2_X1 U601 ( .A(n544), .B(KEYINPUT67), .ZN(n905) );
  NAND2_X1 U602 ( .A1(G126), .A2(n905), .ZN(n545) );
  NAND2_X1 U603 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U604 ( .A1(n548), .A2(n547), .ZN(G164) );
  NAND2_X1 U605 ( .A1(G101), .A2(n901), .ZN(n549) );
  XOR2_X1 U606 ( .A(KEYINPUT23), .B(n549), .Z(n550) );
  XNOR2_X1 U607 ( .A(n550), .B(KEYINPUT68), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G113), .A2(n907), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U610 ( .A1(G137), .A2(n902), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G125), .A2(n905), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U613 ( .A(G2430), .B(G2451), .Z(n558) );
  XNOR2_X1 U614 ( .A(KEYINPUT105), .B(G2443), .ZN(n557) );
  XNOR2_X1 U615 ( .A(n558), .B(n557), .ZN(n565) );
  XOR2_X1 U616 ( .A(G2435), .B(G2446), .Z(n560) );
  XNOR2_X1 U617 ( .A(G2427), .B(G2454), .ZN(n559) );
  XNOR2_X1 U618 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U619 ( .A(n561), .B(G2438), .Z(n563) );
  XNOR2_X1 U620 ( .A(G1341), .B(G1348), .ZN(n562) );
  XNOR2_X1 U621 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U622 ( .A(n565), .B(n564), .ZN(n566) );
  AND2_X1 U623 ( .A1(n566), .A2(G14), .ZN(G401) );
  NAND2_X1 U624 ( .A1(n661), .A2(G64), .ZN(n567) );
  XOR2_X1 U625 ( .A(KEYINPUT71), .B(n567), .Z(n569) );
  NAND2_X1 U626 ( .A1(G52), .A2(n656), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U628 ( .A(KEYINPUT72), .B(n570), .ZN(n575) );
  NAND2_X1 U629 ( .A1(G77), .A2(n519), .ZN(n572) );
  NAND2_X1 U630 ( .A1(G90), .A2(n648), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U632 ( .A(KEYINPUT9), .B(n573), .Z(n574) );
  NOR2_X1 U633 ( .A1(n575), .A2(n574), .ZN(G171) );
  INV_X1 U634 ( .A(G171), .ZN(G301) );
  NAND2_X1 U635 ( .A1(G123), .A2(n905), .ZN(n576) );
  XNOR2_X1 U636 ( .A(n576), .B(KEYINPUT18), .ZN(n583) );
  NAND2_X1 U637 ( .A1(G99), .A2(n901), .ZN(n578) );
  NAND2_X1 U638 ( .A1(G135), .A2(n902), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n907), .A2(G111), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT82), .B(n579), .Z(n580) );
  NOR2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n950) );
  XNOR2_X1 U644 ( .A(G2096), .B(n950), .ZN(n584) );
  OR2_X1 U645 ( .A1(G2100), .A2(n584), .ZN(G156) );
  INV_X1 U646 ( .A(G120), .ZN(G236) );
  INV_X1 U647 ( .A(G69), .ZN(G235) );
  INV_X1 U648 ( .A(G108), .ZN(G238) );
  INV_X1 U649 ( .A(G132), .ZN(G219) );
  INV_X1 U650 ( .A(G82), .ZN(G220) );
  NAND2_X1 U651 ( .A1(G78), .A2(n519), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G91), .A2(n648), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n661), .A2(G65), .ZN(n588) );
  NAND2_X1 U655 ( .A1(G53), .A2(n656), .ZN(n587) );
  NAND2_X1 U656 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U658 ( .A(KEYINPUT74), .B(n591), .ZN(n727) );
  INV_X1 U659 ( .A(n727), .ZN(G299) );
  XOR2_X1 U660 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U661 ( .A1(G94), .A2(G452), .ZN(n592) );
  XNOR2_X1 U662 ( .A(n592), .B(KEYINPUT73), .ZN(G173) );
  NAND2_X1 U663 ( .A1(G7), .A2(G661), .ZN(n593) );
  XOR2_X1 U664 ( .A(n593), .B(KEYINPUT10), .Z(n838) );
  NAND2_X1 U665 ( .A1(n838), .A2(G567), .ZN(n594) );
  XOR2_X1 U666 ( .A(KEYINPUT11), .B(n594), .Z(G234) );
  NAND2_X1 U667 ( .A1(n648), .A2(G81), .ZN(n595) );
  XNOR2_X1 U668 ( .A(n595), .B(KEYINPUT12), .ZN(n597) );
  NAND2_X1 U669 ( .A1(G68), .A2(n519), .ZN(n596) );
  NAND2_X1 U670 ( .A1(n597), .A2(n596), .ZN(n598) );
  XOR2_X1 U671 ( .A(KEYINPUT13), .B(n598), .Z(n602) );
  NAND2_X1 U672 ( .A1(G56), .A2(n661), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n599), .B(KEYINPUT14), .ZN(n600) );
  XNOR2_X1 U674 ( .A(n600), .B(KEYINPUT75), .ZN(n601) );
  NOR2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U676 ( .A1(G43), .A2(n656), .ZN(n603) );
  NAND2_X1 U677 ( .A1(n604), .A2(n603), .ZN(n712) );
  INV_X1 U678 ( .A(n712), .ZN(n1000) );
  NAND2_X1 U679 ( .A1(n1000), .A2(G860), .ZN(G153) );
  NAND2_X1 U680 ( .A1(G868), .A2(G301), .ZN(n614) );
  NAND2_X1 U681 ( .A1(G66), .A2(n661), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G92), .A2(n648), .ZN(n606) );
  NAND2_X1 U683 ( .A1(G54), .A2(n656), .ZN(n605) );
  NAND2_X1 U684 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n519), .A2(G79), .ZN(n607) );
  NOR2_X1 U686 ( .A1(n608), .A2(n520), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U688 ( .A(n611), .B(KEYINPUT15), .ZN(n612) );
  OR2_X1 U689 ( .A1(n997), .A2(G868), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(G284) );
  NAND2_X1 U691 ( .A1(G868), .A2(G286), .ZN(n616) );
  INV_X1 U692 ( .A(G868), .ZN(n676) );
  NAND2_X1 U693 ( .A1(G299), .A2(n676), .ZN(n615) );
  NAND2_X1 U694 ( .A1(n616), .A2(n615), .ZN(G297) );
  INV_X1 U695 ( .A(G559), .ZN(n617) );
  NOR2_X1 U696 ( .A1(G860), .A2(n617), .ZN(n618) );
  XNOR2_X1 U697 ( .A(KEYINPUT81), .B(n618), .ZN(n619) );
  NAND2_X1 U698 ( .A1(n619), .A2(n997), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U700 ( .A1(G868), .A2(n712), .ZN(n623) );
  NAND2_X1 U701 ( .A1(G868), .A2(n997), .ZN(n621) );
  NOR2_X1 U702 ( .A1(G559), .A2(n621), .ZN(n622) );
  NOR2_X1 U703 ( .A1(n623), .A2(n622), .ZN(G282) );
  NAND2_X1 U704 ( .A1(G80), .A2(n519), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G93), .A2(n648), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n661), .A2(G67), .ZN(n627) );
  NAND2_X1 U708 ( .A1(G55), .A2(n656), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n628) );
  OR2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n675) );
  NAND2_X1 U711 ( .A1(G559), .A2(n997), .ZN(n630) );
  XNOR2_X1 U712 ( .A(n630), .B(KEYINPUT83), .ZN(n673) );
  XNOR2_X1 U713 ( .A(n673), .B(n1000), .ZN(n631) );
  NOR2_X1 U714 ( .A1(G860), .A2(n631), .ZN(n632) );
  XOR2_X1 U715 ( .A(n675), .B(n632), .Z(G145) );
  NAND2_X1 U716 ( .A1(G75), .A2(n519), .ZN(n634) );
  NAND2_X1 U717 ( .A1(G88), .A2(n648), .ZN(n633) );
  NAND2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G62), .A2(n661), .ZN(n635) );
  XNOR2_X1 U720 ( .A(n635), .B(KEYINPUT86), .ZN(n637) );
  NAND2_X1 U721 ( .A1(G50), .A2(n656), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U723 ( .A1(n639), .A2(n638), .ZN(G166) );
  INV_X1 U724 ( .A(G166), .ZN(G303) );
  NAND2_X1 U725 ( .A1(G73), .A2(n519), .ZN(n640) );
  XNOR2_X1 U726 ( .A(n640), .B(KEYINPUT2), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G86), .A2(n648), .ZN(n642) );
  NAND2_X1 U728 ( .A1(G48), .A2(n656), .ZN(n641) );
  NAND2_X1 U729 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U730 ( .A1(G61), .A2(n661), .ZN(n643) );
  XNOR2_X1 U731 ( .A(KEYINPUT85), .B(n643), .ZN(n644) );
  NOR2_X1 U732 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U733 ( .A1(n647), .A2(n646), .ZN(G305) );
  NAND2_X1 U734 ( .A1(G72), .A2(n519), .ZN(n650) );
  NAND2_X1 U735 ( .A1(G85), .A2(n648), .ZN(n649) );
  NAND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U737 ( .A1(G60), .A2(n661), .ZN(n651) );
  XOR2_X1 U738 ( .A(KEYINPUT70), .B(n651), .Z(n652) );
  NOR2_X1 U739 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U740 ( .A1(G47), .A2(n656), .ZN(n654) );
  NAND2_X1 U741 ( .A1(n655), .A2(n654), .ZN(G290) );
  NAND2_X1 U742 ( .A1(G651), .A2(G74), .ZN(n658) );
  NAND2_X1 U743 ( .A1(G49), .A2(n656), .ZN(n657) );
  NAND2_X1 U744 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U745 ( .A(KEYINPUT84), .B(n659), .ZN(n660) );
  NOR2_X1 U746 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U747 ( .A1(n662), .A2(G87), .ZN(n663) );
  NAND2_X1 U748 ( .A1(n664), .A2(n663), .ZN(G288) );
  XOR2_X1 U749 ( .A(G303), .B(G305), .Z(n672) );
  XOR2_X1 U750 ( .A(G290), .B(n1000), .Z(n670) );
  XOR2_X1 U751 ( .A(KEYINPUT87), .B(KEYINPUT19), .Z(n666) );
  XOR2_X1 U752 ( .A(n727), .B(KEYINPUT88), .Z(n665) );
  XNOR2_X1 U753 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U754 ( .A(n675), .B(n667), .Z(n668) );
  XNOR2_X1 U755 ( .A(n668), .B(G288), .ZN(n669) );
  XNOR2_X1 U756 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U757 ( .A(n672), .B(n671), .ZN(n868) );
  XNOR2_X1 U758 ( .A(n673), .B(n868), .ZN(n674) );
  NAND2_X1 U759 ( .A1(n674), .A2(G868), .ZN(n678) );
  NAND2_X1 U760 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U761 ( .A1(n678), .A2(n677), .ZN(G295) );
  NAND2_X1 U762 ( .A1(G2078), .A2(G2084), .ZN(n679) );
  XOR2_X1 U763 ( .A(KEYINPUT20), .B(n679), .Z(n680) );
  NAND2_X1 U764 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U765 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U766 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U767 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U768 ( .A1(G220), .A2(G219), .ZN(n683) );
  XOR2_X1 U769 ( .A(KEYINPUT22), .B(n683), .Z(n684) );
  NOR2_X1 U770 ( .A1(G218), .A2(n684), .ZN(n685) );
  XOR2_X1 U771 ( .A(KEYINPUT89), .B(n685), .Z(n686) );
  NAND2_X1 U772 ( .A1(G96), .A2(n686), .ZN(n844) );
  NAND2_X1 U773 ( .A1(n844), .A2(G2106), .ZN(n691) );
  NOR2_X1 U774 ( .A1(G235), .A2(G236), .ZN(n687) );
  XOR2_X1 U775 ( .A(KEYINPUT90), .B(n687), .Z(n688) );
  NOR2_X1 U776 ( .A1(G238), .A2(n688), .ZN(n689) );
  NAND2_X1 U777 ( .A1(G57), .A2(n689), .ZN(n843) );
  NAND2_X1 U778 ( .A1(G567), .A2(n843), .ZN(n690) );
  NAND2_X1 U779 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U780 ( .A(n692), .B(KEYINPUT91), .Z(n842) );
  NAND2_X1 U781 ( .A1(G661), .A2(G483), .ZN(n693) );
  NOR2_X1 U782 ( .A1(n842), .A2(n693), .ZN(n841) );
  NAND2_X1 U783 ( .A1(n841), .A2(G36), .ZN(G176) );
  XNOR2_X1 U784 ( .A(KEYINPUT65), .B(n694), .ZN(n787) );
  NAND2_X1 U785 ( .A1(G160), .A2(G40), .ZN(n788) );
  NOR2_X1 U786 ( .A1(n787), .A2(n788), .ZN(n695) );
  XNOR2_X2 U787 ( .A(KEYINPUT64), .B(n695), .ZN(n722) );
  NAND2_X1 U788 ( .A1(G8), .A2(n737), .ZN(n751) );
  NOR2_X1 U789 ( .A1(n751), .A2(G1966), .ZN(n698) );
  INV_X1 U790 ( .A(G8), .ZN(n696) );
  NOR2_X1 U791 ( .A1(n737), .A2(G2084), .ZN(n749) );
  OR2_X1 U792 ( .A1(n696), .A2(n749), .ZN(n697) );
  OR2_X2 U793 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U794 ( .A(KEYINPUT30), .B(n699), .ZN(n700) );
  XNOR2_X1 U795 ( .A(n701), .B(KEYINPUT97), .ZN(n706) );
  XOR2_X1 U796 ( .A(G2078), .B(KEYINPUT25), .Z(n975) );
  NAND2_X1 U797 ( .A1(n975), .A2(n722), .ZN(n703) );
  NAND2_X1 U798 ( .A1(n737), .A2(G1961), .ZN(n702) );
  NAND2_X1 U799 ( .A1(n703), .A2(n702), .ZN(n734) );
  NAND2_X1 U800 ( .A1(G301), .A2(n734), .ZN(n704) );
  XNOR2_X1 U801 ( .A(KEYINPUT98), .B(n704), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U803 ( .A(n707), .B(KEYINPUT31), .ZN(n752) );
  NAND2_X1 U804 ( .A1(n722), .A2(G1996), .ZN(n708) );
  XNOR2_X1 U805 ( .A(n708), .B(KEYINPUT26), .ZN(n710) );
  NAND2_X1 U806 ( .A1(n737), .A2(G1341), .ZN(n709) );
  NAND2_X1 U807 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U808 ( .A1(n712), .A2(n711), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n718), .A2(n997), .ZN(n717) );
  NAND2_X1 U810 ( .A1(G2067), .A2(n722), .ZN(n714) );
  NAND2_X1 U811 ( .A1(n737), .A2(G1348), .ZN(n713) );
  NAND2_X1 U812 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U813 ( .A(n715), .B(KEYINPUT96), .ZN(n716) );
  NAND2_X1 U814 ( .A1(n717), .A2(n716), .ZN(n720) );
  OR2_X1 U815 ( .A1(n997), .A2(n718), .ZN(n719) );
  NAND2_X1 U816 ( .A1(n720), .A2(n719), .ZN(n726) );
  NAND2_X1 U817 ( .A1(G2072), .A2(n722), .ZN(n721) );
  XNOR2_X1 U818 ( .A(n721), .B(KEYINPUT27), .ZN(n724) );
  XNOR2_X1 U819 ( .A(G1956), .B(KEYINPUT95), .ZN(n922) );
  NOR2_X1 U820 ( .A1(n722), .A2(n922), .ZN(n723) );
  NOR2_X1 U821 ( .A1(n724), .A2(n723), .ZN(n728) );
  NAND2_X1 U822 ( .A1(n728), .A2(n727), .ZN(n725) );
  NAND2_X1 U823 ( .A1(n726), .A2(n725), .ZN(n731) );
  NOR2_X1 U824 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U825 ( .A(n729), .B(KEYINPUT28), .Z(n730) );
  NAND2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n733) );
  OR2_X1 U827 ( .A1(G301), .A2(n734), .ZN(n735) );
  NOR2_X1 U828 ( .A1(n737), .A2(G2090), .ZN(n739) );
  INV_X1 U829 ( .A(n751), .ZN(n766) );
  NOR2_X1 U830 ( .A1(G1971), .A2(n751), .ZN(n738) );
  NOR2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U832 ( .A1(n740), .A2(G303), .ZN(n741) );
  OR2_X1 U833 ( .A1(n696), .A2(n741), .ZN(n743) );
  AND2_X1 U834 ( .A1(n753), .A2(n743), .ZN(n742) );
  NAND2_X1 U835 ( .A1(n752), .A2(n742), .ZN(n747) );
  INV_X1 U836 ( .A(n743), .ZN(n745) );
  AND2_X1 U837 ( .A1(G286), .A2(G8), .ZN(n744) );
  OR2_X1 U838 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U839 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U840 ( .A(n748), .B(KEYINPUT32), .ZN(n759) );
  NAND2_X1 U841 ( .A1(G8), .A2(n749), .ZN(n750) );
  XNOR2_X1 U842 ( .A(KEYINPUT94), .B(n750), .ZN(n757) );
  OR2_X1 U843 ( .A1(G1966), .A2(n751), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n753), .A2(n752), .ZN(n754) );
  AND2_X1 U845 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n759), .A2(n758), .ZN(n761) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n768) );
  NOR2_X1 U849 ( .A1(G1971), .A2(G303), .ZN(n762) );
  NOR2_X1 U850 ( .A1(n768), .A2(n762), .ZN(n1013) );
  XNOR2_X1 U851 ( .A(KEYINPUT100), .B(n1013), .ZN(n764) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n763) );
  AND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n777), .A2(n765), .ZN(n774) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n1012) );
  AND2_X1 U856 ( .A1(n766), .A2(n1012), .ZN(n767) );
  NOR2_X1 U857 ( .A1(KEYINPUT33), .A2(n767), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n768), .A2(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U859 ( .A1(n751), .A2(n769), .ZN(n770) );
  NOR2_X1 U860 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U861 ( .A(G1981), .B(G305), .Z(n1006) );
  XNOR2_X1 U862 ( .A(n775), .B(KEYINPUT101), .ZN(n785) );
  NOR2_X1 U863 ( .A1(G2090), .A2(G303), .ZN(n776) );
  NAND2_X1 U864 ( .A1(G8), .A2(n776), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U866 ( .A1(n779), .A2(n751), .ZN(n783) );
  NOR2_X1 U867 ( .A1(G1981), .A2(G305), .ZN(n780) );
  XOR2_X1 U868 ( .A(n780), .B(KEYINPUT24), .Z(n781) );
  OR2_X1 U869 ( .A1(n751), .A2(n781), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U871 ( .A1(n785), .A2(n784), .ZN(n786) );
  INV_X1 U872 ( .A(n786), .ZN(n819) );
  INV_X1 U873 ( .A(n787), .ZN(n789) );
  NOR2_X1 U874 ( .A1(n789), .A2(n788), .ZN(n833) );
  NAND2_X1 U875 ( .A1(G116), .A2(n907), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G128), .A2(n905), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U878 ( .A(n792), .B(KEYINPUT35), .ZN(n797) );
  NAND2_X1 U879 ( .A1(G104), .A2(n901), .ZN(n794) );
  NAND2_X1 U880 ( .A1(G140), .A2(n902), .ZN(n793) );
  NAND2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U882 ( .A(KEYINPUT34), .B(n795), .Z(n796) );
  NAND2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U884 ( .A(n798), .B(KEYINPUT36), .Z(n883) );
  XNOR2_X1 U885 ( .A(KEYINPUT37), .B(G2067), .ZN(n820) );
  NOR2_X1 U886 ( .A1(n883), .A2(n820), .ZN(n957) );
  NAND2_X1 U887 ( .A1(n833), .A2(n957), .ZN(n828) );
  NAND2_X1 U888 ( .A1(G107), .A2(n907), .ZN(n799) );
  XNOR2_X1 U889 ( .A(n799), .B(KEYINPUT92), .ZN(n802) );
  NAND2_X1 U890 ( .A1(G131), .A2(n902), .ZN(n800) );
  XOR2_X1 U891 ( .A(KEYINPUT93), .B(n800), .Z(n801) );
  NAND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n806) );
  NAND2_X1 U893 ( .A1(G95), .A2(n901), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G119), .A2(n905), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n894) );
  INV_X1 U897 ( .A(G1991), .ZN(n855) );
  NOR2_X1 U898 ( .A1(n894), .A2(n855), .ZN(n815) );
  NAND2_X1 U899 ( .A1(n901), .A2(G105), .ZN(n807) );
  XNOR2_X1 U900 ( .A(n807), .B(KEYINPUT38), .ZN(n809) );
  NAND2_X1 U901 ( .A1(G117), .A2(n907), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n813) );
  NAND2_X1 U903 ( .A1(G141), .A2(n902), .ZN(n811) );
  NAND2_X1 U904 ( .A1(G129), .A2(n905), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  OR2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n882) );
  AND2_X1 U907 ( .A1(G1996), .A2(n882), .ZN(n814) );
  NOR2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n955) );
  INV_X1 U909 ( .A(n955), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n816), .A2(n833), .ZN(n821) );
  AND2_X1 U911 ( .A1(n828), .A2(n821), .ZN(n818) );
  XNOR2_X1 U912 ( .A(G1986), .B(G290), .ZN(n999) );
  NAND2_X1 U913 ( .A1(n999), .A2(n833), .ZN(n817) );
  NAND2_X1 U914 ( .A1(n819), .A2(n518), .ZN(n836) );
  AND2_X1 U915 ( .A1(n883), .A2(n820), .ZN(n960) );
  INV_X1 U916 ( .A(n821), .ZN(n824) );
  AND2_X1 U917 ( .A1(n855), .A2(n894), .ZN(n953) );
  NOR2_X1 U918 ( .A1(G1986), .A2(G290), .ZN(n822) );
  NOR2_X1 U919 ( .A1(n953), .A2(n822), .ZN(n823) );
  NOR2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n826) );
  NOR2_X1 U921 ( .A1(n882), .A2(G1996), .ZN(n825) );
  XNOR2_X1 U922 ( .A(n825), .B(KEYINPUT102), .ZN(n963) );
  NOR2_X1 U923 ( .A1(n826), .A2(n963), .ZN(n827) );
  XNOR2_X1 U924 ( .A(n827), .B(KEYINPUT39), .ZN(n829) );
  NAND2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U926 ( .A(KEYINPUT103), .B(n830), .ZN(n831) );
  NOR2_X1 U927 ( .A1(n960), .A2(n831), .ZN(n832) );
  XOR2_X1 U928 ( .A(KEYINPUT104), .B(n832), .Z(n834) );
  NAND2_X1 U929 ( .A1(n834), .A2(n833), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U931 ( .A(n837), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n838), .ZN(G217) );
  INV_X1 U933 ( .A(n838), .ZN(G223) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U935 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U937 ( .A1(n841), .A2(n840), .ZN(G188) );
  INV_X1 U938 ( .A(n842), .ZN(G319) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  NOR2_X1 U941 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  XOR2_X1 U943 ( .A(KEYINPUT43), .B(G2678), .Z(n846) );
  XNOR2_X1 U944 ( .A(KEYINPUT107), .B(KEYINPUT106), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U946 ( .A(KEYINPUT42), .B(G2072), .Z(n848) );
  XNOR2_X1 U947 ( .A(G2067), .B(G2090), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U949 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U950 ( .A(G2096), .B(G2100), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n854) );
  XOR2_X1 U952 ( .A(G2078), .B(G2084), .Z(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(G227) );
  XOR2_X1 U954 ( .A(G1976), .B(G1971), .Z(n857) );
  XOR2_X1 U955 ( .A(G1996), .B(n855), .Z(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n867) );
  XOR2_X1 U957 ( .A(KEYINPUT110), .B(KEYINPUT108), .Z(n859) );
  XNOR2_X1 U958 ( .A(G1961), .B(G2474), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U960 ( .A(G1981), .B(G1956), .Z(n861) );
  XNOR2_X1 U961 ( .A(G1986), .B(G1966), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U963 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U964 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(G229) );
  XNOR2_X1 U967 ( .A(G286), .B(n868), .ZN(n870) );
  XOR2_X1 U968 ( .A(G301), .B(n997), .Z(n869) );
  XNOR2_X1 U969 ( .A(n870), .B(n869), .ZN(n871) );
  NOR2_X1 U970 ( .A1(G37), .A2(n871), .ZN(G397) );
  NAND2_X1 U971 ( .A1(n901), .A2(G100), .ZN(n872) );
  XNOR2_X1 U972 ( .A(KEYINPUT112), .B(n872), .ZN(n875) );
  NAND2_X1 U973 ( .A1(n907), .A2(G112), .ZN(n873) );
  XOR2_X1 U974 ( .A(KEYINPUT111), .B(n873), .Z(n874) );
  NAND2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n876), .B(KEYINPUT113), .ZN(n878) );
  NAND2_X1 U977 ( .A1(G136), .A2(n902), .ZN(n877) );
  NAND2_X1 U978 ( .A1(n878), .A2(n877), .ZN(n881) );
  NAND2_X1 U979 ( .A1(n905), .A2(G124), .ZN(n879) );
  XOR2_X1 U980 ( .A(KEYINPUT44), .B(n879), .Z(n880) );
  NOR2_X1 U981 ( .A1(n881), .A2(n880), .ZN(G162) );
  XOR2_X1 U982 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n885) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n898) );
  NAND2_X1 U985 ( .A1(G118), .A2(n907), .ZN(n887) );
  NAND2_X1 U986 ( .A1(G130), .A2(n905), .ZN(n886) );
  NAND2_X1 U987 ( .A1(n887), .A2(n886), .ZN(n893) );
  NAND2_X1 U988 ( .A1(n901), .A2(G106), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n888), .B(KEYINPUT114), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G142), .A2(n902), .ZN(n889) );
  NAND2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U992 ( .A(KEYINPUT45), .B(n891), .Z(n892) );
  NOR2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n895) );
  XOR2_X1 U994 ( .A(n895), .B(n894), .Z(n896) );
  XNOR2_X1 U995 ( .A(n896), .B(n950), .ZN(n897) );
  XOR2_X1 U996 ( .A(n898), .B(n897), .Z(n900) );
  XNOR2_X1 U997 ( .A(G164), .B(G160), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n900), .B(n899), .ZN(n914) );
  NAND2_X1 U999 ( .A1(G103), .A2(n901), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(G139), .A2(n902), .ZN(n903) );
  NAND2_X1 U1001 ( .A1(n904), .A2(n903), .ZN(n912) );
  NAND2_X1 U1002 ( .A1(n905), .A2(G127), .ZN(n906) );
  XOR2_X1 U1003 ( .A(KEYINPUT115), .B(n906), .Z(n909) );
  NAND2_X1 U1004 ( .A1(n907), .A2(G115), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1006 ( .A(KEYINPUT47), .B(n910), .Z(n911) );
  NOR2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(n945) );
  XOR2_X1 U1008 ( .A(n945), .B(G162), .Z(n913) );
  XNOR2_X1 U1009 ( .A(n914), .B(n913), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G37), .A2(n915), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(KEYINPUT116), .B(n916), .ZN(G395) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n918), .ZN(n919) );
  AND2_X1 U1015 ( .A1(G319), .A2(n919), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(G397), .A2(G395), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1020 ( .A(G20), .B(n922), .ZN(n926) );
  XNOR2_X1 U1021 ( .A(G1341), .B(G19), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(G1981), .B(G6), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n929) );
  XOR2_X1 U1025 ( .A(KEYINPUT59), .B(G1348), .Z(n927) );
  XNOR2_X1 U1026 ( .A(G4), .B(n927), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(KEYINPUT60), .B(n930), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(G1966), .B(G21), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(G1961), .B(G5), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n941) );
  XNOR2_X1 U1033 ( .A(G1971), .B(G22), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(G23), .B(G1976), .ZN(n935) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n938) );
  XOR2_X1 U1036 ( .A(G1986), .B(G24), .Z(n937) );
  NAND2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1038 ( .A(KEYINPUT58), .B(n939), .ZN(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(KEYINPUT61), .B(n942), .ZN(n943) );
  INV_X1 U1041 ( .A(G16), .ZN(n1021) );
  NAND2_X1 U1042 ( .A1(n943), .A2(n1021), .ZN(n944) );
  NAND2_X1 U1043 ( .A1(n944), .A2(G11), .ZN(n996) );
  XOR2_X1 U1044 ( .A(G2072), .B(n945), .Z(n947) );
  XOR2_X1 U1045 ( .A(G164), .B(G2078), .Z(n946) );
  NOR2_X1 U1046 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1047 ( .A(KEYINPUT118), .B(n948), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(n949), .B(KEYINPUT50), .ZN(n962) );
  XNOR2_X1 U1049 ( .A(G160), .B(G2084), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1051 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT117), .B(n958), .ZN(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n967) );
  XOR2_X1 U1057 ( .A(G2090), .B(G162), .Z(n964) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(KEYINPUT51), .B(n965), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT52), .B(n968), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n989) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n989), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n970), .A2(G29), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT120), .B(n971), .ZN(n994) );
  XOR2_X1 U1066 ( .A(G29), .B(KEYINPUT122), .Z(n992) );
  XOR2_X1 U1067 ( .A(G25), .B(G1991), .Z(n972) );
  NAND2_X1 U1068 ( .A1(n972), .A2(G28), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(G2067), .B(G26), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(G33), .B(G2072), .ZN(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(G1996), .B(G32), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(G27), .B(n975), .ZN(n976) );
  NOR2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1077 ( .A(KEYINPUT53), .B(n982), .Z(n986) );
  XNOR2_X1 U1078 ( .A(KEYINPUT54), .B(G34), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(n983), .B(KEYINPUT121), .ZN(n984) );
  XNOR2_X1 U1080 ( .A(G2084), .B(n984), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(G35), .B(G2090), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n990) );
  XOR2_X1 U1084 ( .A(n990), .B(n989), .Z(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n1026) );
  XOR2_X1 U1088 ( .A(G1348), .B(n997), .Z(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(G1341), .B(KEYINPUT125), .ZN(n1001) );
  XOR2_X1 U1091 ( .A(n1001), .B(n1000), .Z(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1009) );
  XOR2_X1 U1093 ( .A(G1966), .B(KEYINPUT123), .Z(n1004) );
  XNOR2_X1 U1094 ( .A(G168), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1096 ( .A(KEYINPUT57), .B(n1007), .Z(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1018) );
  XOR2_X1 U1098 ( .A(G299), .B(G1956), .Z(n1011) );
  NAND2_X1 U1099 ( .A1(G303), .A2(G1971), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(n1016), .B(KEYINPUT124), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(G1961), .B(G171), .Z(n1019) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(n1021), .B(KEYINPUT56), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1109 ( .A(KEYINPUT126), .B(n1024), .Z(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(n1027), .B(KEYINPUT62), .ZN(n1028) );
  XOR2_X1 U1112 ( .A(KEYINPUT127), .B(n1028), .Z(G150) );
  INV_X1 U1113 ( .A(G150), .ZN(G311) );
endmodule

