//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n524, new_n525, new_n526, new_n527,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n543, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1208,
    new_n1209, new_n1210, new_n1212, new_n1213;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT69), .Z(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(KEYINPUT70), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n455), .A2(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(new_n459), .B2(new_n460), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n465), .A2(new_n467), .A3(G137), .A4(new_n463), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n464), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n465), .A2(new_n467), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n479), .A2(new_n482), .A3(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n465), .A2(new_n467), .A3(G126), .A4(G2105), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n463), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n476), .A2(new_n494), .A3(G138), .A4(new_n463), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT6), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G651), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(G50), .A3(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n506), .A2(new_n508), .A3(new_n498), .A4(new_n500), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n510), .A2(new_n497), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n504), .A2(new_n513), .ZN(G166));
  AND2_X1   g089(.A1(new_n501), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G51), .ZN(new_n516));
  INV_X1    g091(.A(new_n512), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G89), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n516), .A2(new_n518), .A3(new_n519), .A4(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  XNOR2_X1  g098(.A(KEYINPUT72), .B(G52), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n515), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n517), .A2(G90), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n525), .B(new_n526), .C1(new_n497), .C2(new_n527), .ZN(G301));
  INV_X1    g103(.A(G301), .ZN(G171));
  NAND2_X1  g104(.A1(new_n506), .A2(new_n508), .ZN(new_n530));
  INV_X1    g105(.A(G56), .ZN(new_n531));
  INV_X1    g106(.A(G68), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n530), .A2(new_n531), .B1(new_n532), .B2(new_n505), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI221_X1 g110(.A(KEYINPUT73), .B1(new_n532), .B2(new_n505), .C1(new_n530), .C2(new_n531), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(G651), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g112(.A(KEYINPUT74), .B(G43), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n515), .A2(new_n538), .B1(G81), .B2(new_n517), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  AND3_X1   g117(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G36), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n543), .A2(new_n546), .ZN(G188));
  NAND3_X1  g122(.A1(new_n501), .A2(G53), .A3(G543), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT9), .ZN(new_n549));
  INV_X1    g124(.A(G65), .ZN(new_n550));
  INV_X1    g125(.A(G78), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n530), .A2(new_n550), .B1(new_n551), .B2(new_n505), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT76), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT76), .ZN(new_n554));
  OAI221_X1 g129(.A(new_n554), .B1(new_n551), .B2(new_n505), .C1(new_n530), .C2(new_n550), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n553), .A2(G651), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G91), .ZN(new_n557));
  OR3_X1    g132(.A1(new_n512), .A2(KEYINPUT75), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT75), .B1(new_n512), .B2(new_n557), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n549), .A2(new_n556), .A3(new_n560), .ZN(G299));
  INV_X1    g136(.A(G166), .ZN(G303));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n501), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G49), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n517), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n501), .A2(KEYINPUT77), .A3(G49), .A4(G543), .ZN(new_n569));
  NAND4_X1  g144(.A1(new_n566), .A2(new_n567), .A3(new_n568), .A4(new_n569), .ZN(G288));
  NAND4_X1  g145(.A1(new_n498), .A2(new_n500), .A3(G48), .A4(G543), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n512), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n506), .A2(new_n508), .A3(G61), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n497), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n515), .A2(G47), .B1(G85), .B2(new_n517), .ZN(new_n579));
  NAND2_X1  g154(.A1(G72), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G60), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n530), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n582), .A2(KEYINPUT78), .A3(G651), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n579), .A2(new_n585), .A3(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  INV_X1    g163(.A(G92), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n512), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n515), .A2(G54), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  INV_X1    g168(.A(G79), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n530), .A2(new_n593), .B1(new_n594), .B2(new_n505), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(KEYINPUT79), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n597));
  OAI221_X1 g172(.A(new_n597), .B1(new_n594), .B2(new_n505), .C1(new_n530), .C2(new_n593), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(G651), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n591), .A2(new_n592), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n588), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n588), .B1(new_n601), .B2(G868), .ZN(G321));
  INV_X1    g178(.A(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(G299), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(new_n604), .B2(G168), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n540), .A2(new_n604), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n600), .A2(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(new_n604), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT80), .Z(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g189(.A(new_n472), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT12), .B1(new_n480), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT12), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n476), .A2(new_n617), .A3(new_n472), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n478), .A2(G123), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n481), .A2(G135), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n463), .A2(G111), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(G2096), .Z(new_n627));
  NAND2_X1  g202(.A1(new_n621), .A2(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(KEYINPUT15), .B(G2435), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2438), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2430), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT81), .B(KEYINPUT14), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G14), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n644), .B1(new_n648), .B2(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n646), .A2(new_n647), .ZN(new_n653));
  AOI21_X1  g228(.A(KEYINPUT18), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n651), .B(new_n654), .Z(G227));
  XOR2_X1   g230(.A(G1971), .B(G1976), .Z(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  AOI22_X1  g239(.A1(new_n662), .A2(new_n663), .B1(new_n658), .B2(new_n664), .ZN(new_n665));
  OR3_X1    g240(.A1(new_n658), .A2(new_n661), .A3(new_n664), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n666), .C1(new_n663), .C2(new_n662), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  INV_X1    g245(.A(G1981), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1986), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n669), .B(new_n673), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G229));
  NAND2_X1  g250(.A1(new_n541), .A2(G16), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(G16), .B2(G19), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT87), .B(G1341), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G5), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(G171), .B2(new_n681), .ZN(new_n683));
  INV_X1    g258(.A(G1961), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n677), .A2(new_n679), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(G28), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(G28), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g266(.A1(new_n680), .A2(new_n685), .A3(new_n686), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(G162), .A2(G29), .ZN(new_n693));
  OR2_X1    g268(.A1(G29), .A2(G35), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT29), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n693), .A2(new_n697), .A3(new_n694), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G2090), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g276(.A(G29), .B1(new_n470), .B2(new_n474), .ZN(new_n702));
  INV_X1    g277(.A(G2084), .ZN(new_n703));
  OR2_X1    g278(.A1(KEYINPUT24), .A2(G34), .ZN(new_n704));
  NAND2_X1  g279(.A1(KEYINPUT24), .A2(G34), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n704), .A2(new_n690), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n702), .A2(new_n703), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n696), .A2(G2090), .A3(new_n698), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n703), .B1(new_n702), .B2(new_n706), .ZN(new_n709));
  NOR2_X1   g284(.A1(G29), .A2(G32), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n472), .A2(G105), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n476), .A2(new_n463), .ZN(new_n712));
  INV_X1    g287(.A(G141), .ZN(new_n713));
  INV_X1    g288(.A(G129), .ZN(new_n714));
  OAI221_X1 g289(.A(new_n711), .B1(new_n712), .B2(new_n713), .C1(new_n714), .C2(new_n477), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT90), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT26), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n710), .B1(new_n720), .B2(G29), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT27), .B(G1996), .Z(new_n722));
  AOI21_X1  g297(.A(new_n709), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n701), .A2(new_n707), .A3(new_n708), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(G168), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G16), .B2(G21), .ZN(new_n726));
  INV_X1    g301(.A(G1966), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g303(.A1(new_n692), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(G29), .A2(G33), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n472), .A2(G103), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT88), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT25), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NAND2_X1  g310(.A1(G115), .A2(G2104), .ZN(new_n736));
  INV_X1    g311(.A(G127), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n480), .B2(new_n737), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n738), .A2(G2105), .B1(new_n481), .B2(G139), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n734), .A2(new_n735), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n730), .B1(new_n740), .B2(new_n690), .ZN(new_n741));
  INV_X1    g316(.A(G2072), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT89), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n681), .A2(G4), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n601), .B2(new_n681), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1348), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n690), .A2(G26), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n478), .A2(G128), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n481), .A2(G140), .ZN(new_n751));
  OR2_X1    g326(.A1(G104), .A2(G2105), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n752), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n749), .B1(new_n754), .B2(new_n690), .ZN(new_n755));
  MUX2_X1   g330(.A(new_n749), .B(new_n755), .S(KEYINPUT28), .Z(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(G2067), .ZN(new_n757));
  NAND2_X1  g332(.A1(G299), .A2(G16), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n681), .A2(KEYINPUT23), .A3(G20), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT23), .ZN(new_n760));
  INV_X1    g335(.A(G20), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(G16), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n758), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G1956), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n741), .A2(new_n742), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n721), .A2(new_n722), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n756), .B2(G2067), .ZN(new_n768));
  AND4_X1   g343(.A1(new_n757), .A2(new_n765), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n726), .A2(new_n727), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT91), .Z(new_n771));
  NAND4_X1  g346(.A1(new_n729), .A2(new_n748), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT36), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT86), .ZN(new_n774));
  NOR2_X1   g349(.A1(G16), .A2(G24), .ZN(new_n775));
  INV_X1    g350(.A(G290), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(G16), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n774), .B1(new_n777), .B2(G1986), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n681), .A2(G23), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G288), .B2(G16), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT33), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n780), .A2(new_n781), .ZN(new_n784));
  OAI21_X1  g359(.A(G1976), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(new_n784), .ZN(new_n786));
  INV_X1    g361(.A(G1976), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n786), .A2(new_n787), .A3(new_n782), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n504), .A2(new_n681), .A3(new_n513), .ZN(new_n790));
  NOR2_X1   g365(.A1(G16), .A2(G22), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n792), .A2(G1971), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n681), .A2(G6), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n577), .B2(new_n681), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT32), .B(G1981), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G1971), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n790), .A2(new_n798), .A3(new_n791), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n793), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n789), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n778), .B1(new_n801), .B2(KEYINPUT34), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n777), .A2(G1986), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT34), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n789), .A2(new_n800), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n690), .A2(G25), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n807));
  INV_X1    g382(.A(G107), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G2105), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT83), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n478), .A2(G119), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n481), .A2(G131), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT84), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT84), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n811), .A2(new_n817), .A3(new_n812), .A4(new_n813), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n806), .B1(new_n820), .B2(new_n690), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT35), .B(G1991), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT85), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n821), .B(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n802), .A2(new_n803), .A3(new_n805), .A4(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n772), .B1(new_n773), .B2(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n826), .A2(new_n773), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n626), .A2(new_n690), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(G11), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n690), .A2(G27), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(G164), .B2(new_n690), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT93), .ZN(new_n835));
  INV_X1    g410(.A(G2078), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n832), .A2(new_n837), .ZN(G311));
  AND2_X1   g413(.A1(new_n826), .A2(new_n773), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n826), .A2(new_n773), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n839), .A2(new_n840), .A3(new_n772), .ZN(new_n841));
  INV_X1    g416(.A(new_n837), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n841), .A2(new_n842), .A3(new_n829), .A4(new_n831), .ZN(G150));
  NAND3_X1  g418(.A1(new_n501), .A2(G55), .A3(G543), .ZN(new_n844));
  INV_X1    g419(.A(G93), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  OAI221_X1 g421(.A(new_n844), .B1(new_n845), .B2(new_n512), .C1(new_n846), .C2(new_n497), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(G860), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT95), .B(KEYINPUT37), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n846), .A2(new_n497), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n515), .A2(G55), .B1(G93), .B2(new_n517), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n540), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n847), .A2(new_n537), .A3(new_n539), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT39), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n600), .A2(new_n608), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT94), .B(KEYINPUT38), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n856), .B(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n850), .B1(new_n860), .B2(G860), .ZN(G145));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n619), .B(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(new_n815), .B2(new_n818), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n478), .A2(G130), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n481), .A2(G142), .ZN(new_n867));
  OR2_X1    g442(.A1(G106), .A2(G2105), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(G2104), .C1(G118), .C2(new_n463), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n815), .A2(new_n818), .A3(new_n863), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n865), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n872), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n870), .B1(new_n874), .B2(new_n864), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n740), .B(KEYINPUT96), .ZN(new_n876));
  INV_X1    g451(.A(new_n715), .ZN(new_n877));
  INV_X1    g452(.A(new_n719), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n750), .A2(new_n751), .A3(new_n753), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n754), .B1(new_n715), .B2(new_n719), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n493), .A2(new_n495), .ZN(new_n882));
  INV_X1    g457(.A(new_n491), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n880), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n880), .B2(new_n881), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n876), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n740), .A2(KEYINPUT96), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n886), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n880), .A2(new_n881), .A3(new_n884), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n873), .B(new_n875), .C1(new_n887), .C2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n626), .B(G160), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G162), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT100), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n887), .A2(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n875), .A2(new_n873), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT99), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n740), .A2(KEYINPUT96), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n890), .A2(new_n889), .A3(new_n900), .A4(new_n891), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n888), .B1(new_n885), .B2(new_n886), .ZN(new_n902));
  AND4_X1   g477(.A1(KEYINPUT99), .A2(new_n898), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  OAI211_X1 g478(.A(new_n893), .B(new_n896), .C1(new_n899), .C2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n898), .A2(new_n901), .A3(new_n902), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n893), .A2(KEYINPUT98), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT98), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n897), .A2(new_n907), .A3(new_n898), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n908), .A3(new_n895), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n904), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g487(.A1(G299), .A2(KEYINPUT102), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n549), .A2(new_n914), .A3(new_n556), .A4(new_n560), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n601), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n600), .A2(G299), .A3(KEYINPUT102), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(KEYINPUT41), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n853), .B2(new_n854), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n853), .A2(new_n922), .A3(new_n854), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n611), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n925), .ZN(new_n927));
  INV_X1    g502(.A(new_n611), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n927), .A2(new_n928), .A3(new_n923), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n918), .B(new_n921), .C1(new_n926), .C2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n919), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n928), .B1(new_n927), .B2(new_n923), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n924), .A2(new_n611), .A3(new_n925), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n776), .A2(G288), .ZN(new_n938));
  INV_X1    g513(.A(G288), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(G290), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(KEYINPUT103), .A3(new_n940), .ZN(new_n944));
  XNOR2_X1  g519(.A(G166), .B(new_n577), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n945), .A2(new_n944), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n948), .A2(KEYINPUT42), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT42), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n930), .A2(KEYINPUT104), .A3(new_n934), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n937), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT104), .B1(new_n930), .B2(new_n934), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(new_n951), .A3(new_n949), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n604), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n847), .A2(G868), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(G295));
  NAND2_X1  g534(.A1(new_n953), .A2(new_n952), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n956), .B1(new_n960), .B2(new_n955), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(G868), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n963));
  INV_X1    g538(.A(new_n958), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT105), .B1(new_n957), .B2(new_n958), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(G331));
  NOR2_X1   g542(.A1(G301), .A2(KEYINPUT106), .ZN(new_n968));
  INV_X1    g543(.A(new_n854), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n847), .B1(new_n537), .B2(new_n539), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n853), .B(new_n854), .C1(KEYINPUT106), .C2(G301), .ZN(new_n972));
  AOI21_X1  g547(.A(G168), .B1(KEYINPUT106), .B2(G301), .ZN(new_n973));
  AND3_X1   g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n971), .B2(new_n972), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n931), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT107), .ZN(new_n977));
  INV_X1    g552(.A(new_n948), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n979), .B(new_n931), .C1(new_n974), .C2(new_n975), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n971), .A2(new_n972), .ZN(new_n981));
  INV_X1    g556(.A(new_n973), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n983), .A2(new_n921), .A3(new_n918), .A4(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n977), .A2(new_n978), .A3(new_n980), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n976), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n948), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n988), .A3(new_n910), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n977), .A2(new_n980), .A3(new_n985), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n948), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n993), .A2(KEYINPUT43), .A3(new_n910), .A4(new_n986), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT44), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n991), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AND4_X1   g571(.A1(KEYINPUT43), .A2(new_n986), .A3(new_n988), .A4(new_n910), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(new_n910), .A3(new_n986), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n990), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n996), .B1(new_n999), .B2(new_n995), .ZN(G397));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n879), .B(G2067), .ZN(new_n1002));
  INV_X1    g577(.A(G1996), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n720), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  OR3_X1    g580(.A1(G164), .A2(KEYINPUT108), .A3(G1384), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT108), .B1(G164), .B2(G1384), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  INV_X1    g584(.A(new_n474), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n468), .A2(new_n469), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(G2105), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1012), .A3(G40), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT109), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n1015));
  NAND3_X1  g590(.A1(G160), .A2(new_n1015), .A3(G40), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1008), .A2(KEYINPUT110), .A3(new_n1009), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1006), .A2(new_n1009), .A3(new_n1007), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1015), .B1(G160), .B2(G40), .ZN(new_n1021));
  INV_X1    g596(.A(G40), .ZN(new_n1022));
  NOR4_X1   g597(.A1(new_n470), .A2(new_n474), .A3(KEYINPUT109), .A4(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1019), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1018), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1018), .A2(KEYINPUT112), .A3(new_n1025), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1005), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1018), .A2(new_n1003), .A3(new_n1025), .ZN(new_n1031));
  INV_X1    g606(.A(new_n720), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1001), .B1(new_n1030), .B2(new_n1033), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1018), .A2(KEYINPUT112), .A3(new_n1025), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT112), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1036));
  OAI22_X1  g611(.A1(new_n1035), .A2(new_n1036), .B1(new_n1004), .B2(new_n1002), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1033), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(KEYINPUT113), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n819), .A3(new_n823), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n820), .A2(new_n824), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1034), .A2(new_n1039), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1026), .ZN(new_n1045));
  NOR2_X1   g620(.A1(G290), .A2(G1986), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(KEYINPUT111), .ZN(new_n1047));
  NAND2_X1  g622(.A1(G290), .A2(G1986), .ZN(new_n1048));
  XOR2_X1   g623(.A(new_n1047), .B(new_n1048), .Z(new_n1049));
  AOI21_X1  g624(.A(new_n1044), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1009), .B1(G164), .B2(G1384), .ZN(new_n1051));
  INV_X1    g626(.A(G1384), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n884), .A2(KEYINPUT45), .A3(new_n1052), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1051), .B(new_n1053), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT114), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1017), .A2(new_n1056), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1057));
  AOI21_X1  g632(.A(G1971), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n884), .A2(new_n1060), .A3(new_n1052), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1059), .B(new_n1061), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(G2090), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G8), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G166), .A2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT115), .B(KEYINPUT55), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1066), .B(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1064), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT118), .B1(new_n1062), .B2(G2084), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1073), .A2(new_n1074), .A3(new_n703), .A4(new_n1017), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1054), .A2(new_n727), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1077), .A2(G8), .A3(G168), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n577), .A2(new_n671), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT49), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n577), .A2(new_n671), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1081), .B1(new_n1082), .B2(KEYINPUT116), .ZN(new_n1083));
  NOR3_X1   g658(.A1(new_n573), .A2(new_n576), .A3(G1981), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1084), .A2(new_n1085), .A3(KEYINPUT49), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1080), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(G164), .A2(G1384), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1065), .B1(new_n1017), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1082), .A2(KEYINPUT116), .A3(new_n1081), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1080), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT49), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1087), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1088), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n567), .A2(new_n568), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1096), .A2(G1976), .A3(new_n566), .A4(new_n569), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(G8), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT52), .ZN(new_n1099));
  AOI21_X1  g674(.A(KEYINPUT52), .B1(G288), .B2(new_n787), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1089), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1094), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1069), .B(G8), .C1(new_n1058), .C2(new_n1063), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1071), .A2(new_n1079), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT63), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1102), .B(KEYINPUT117), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1108), .A2(KEYINPUT63), .A3(new_n1104), .A4(new_n1071), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1109), .B2(new_n1078), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1072), .A2(new_n1075), .A3(G168), .A4(new_n1076), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1065), .A2(KEYINPUT122), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT51), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1077), .A2(G8), .A3(G286), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1111), .A2(new_n1116), .A3(new_n1112), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT62), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1071), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1055), .A2(new_n836), .A3(new_n1057), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n1122));
  XNOR2_X1  g697(.A(KEYINPUT124), .B(G1961), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1121), .A2(new_n1122), .B1(new_n1062), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n1125));
  OR3_X1    g700(.A1(new_n1054), .A2(new_n1125), .A3(G2078), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1054), .B2(G2078), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(KEYINPUT53), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(G301), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1114), .A2(new_n1130), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1119), .A2(new_n1120), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1104), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1094), .A2(new_n787), .A3(new_n939), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n1082), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1108), .A2(new_n1133), .B1(new_n1089), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1110), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1137));
  XNOR2_X1  g712(.A(G301), .B(KEYINPUT54), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1013), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n836), .B1(new_n1140), .B2(KEYINPUT125), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1122), .B1(new_n1140), .B2(KEYINPUT125), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1020), .A2(new_n1053), .A3(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1124), .B(new_n1139), .C1(new_n1141), .C2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1145), .A2(new_n1138), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1120), .A2(new_n1144), .A3(new_n1146), .A4(new_n1118), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT119), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT57), .B1(G299), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1062), .A2(new_n764), .ZN(new_n1151));
  NAND3_X1  g726(.A1(G299), .A2(new_n1148), .A3(KEYINPUT57), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT56), .B(G2072), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1017), .A2(new_n1051), .A3(new_n1053), .A4(new_n1153), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .A4(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT120), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1152), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(new_n1149), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1158), .A2(new_n1159), .A3(new_n1151), .A4(new_n1154), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1150), .A2(new_n1152), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  OR2_X1    g739(.A1(new_n1095), .A2(G2067), .ZN(new_n1165));
  INV_X1    g740(.A(G1348), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1062), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n600), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1156), .B(new_n1160), .C1(new_n1164), .C2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1160), .A2(new_n1156), .A3(new_n1163), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1155), .A2(KEYINPUT61), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1170), .A2(new_n1171), .B1(new_n1163), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT121), .ZN(new_n1174));
  OR3_X1    g749(.A1(new_n1054), .A2(new_n1174), .A3(G1996), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1174), .B1(new_n1054), .B2(G1996), .ZN(new_n1176));
  XOR2_X1   g751(.A(KEYINPUT58), .B(G1341), .Z(new_n1177));
  NAND2_X1  g752(.A1(new_n1095), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(new_n541), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT59), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1179), .A2(new_n1182), .A3(new_n541), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1185));
  OR3_X1    g760(.A1(new_n1185), .A2(KEYINPUT60), .A3(new_n600), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1185), .A2(new_n601), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT60), .B1(new_n1187), .B2(new_n1168), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1173), .A2(new_n1184), .A3(new_n1186), .A4(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1147), .B1(new_n1169), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1050), .B1(new_n1137), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1034), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1192));
  OR2_X1    g767(.A1(new_n879), .A2(G2067), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1192), .A2(new_n1193), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1040), .B1(new_n1032), .B2(new_n1002), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT47), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1031), .B(KEYINPUT46), .ZN(new_n1197));
  AND3_X1   g772(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1196), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1018), .A2(new_n1025), .A3(new_n1046), .ZN(new_n1201));
  XOR2_X1   g776(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1202));
  XNOR2_X1  g777(.A(new_n1201), .B(new_n1202), .ZN(new_n1203));
  AND4_X1   g778(.A1(new_n1034), .A2(new_n1039), .A3(new_n1043), .A4(new_n1203), .ZN(new_n1204));
  NOR3_X1   g779(.A1(new_n1194), .A2(new_n1200), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1191), .A2(new_n1205), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g781(.A(G227), .ZN(new_n1208));
  NAND4_X1  g782(.A1(new_n991), .A2(new_n994), .A3(G319), .A4(new_n1208), .ZN(new_n1209));
  NAND3_X1  g783(.A1(new_n911), .A2(new_n642), .A3(new_n674), .ZN(new_n1210));
  NOR2_X1   g784(.A1(new_n1209), .A2(new_n1210), .ZN(G308));
  AND2_X1   g785(.A1(new_n991), .A2(new_n994), .ZN(new_n1212));
  AND3_X1   g786(.A1(new_n911), .A2(new_n642), .A3(new_n674), .ZN(new_n1213));
  NAND4_X1  g787(.A1(new_n1212), .A2(new_n1213), .A3(G319), .A4(new_n1208), .ZN(G225));
endmodule


