//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT14), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT14), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT87), .ZN(new_n210));
  NAND2_X1  g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n209), .A2(KEYINPUT87), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n204), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(KEYINPUT88), .B(KEYINPUT15), .Z(new_n215));
  AOI21_X1  g014(.A(new_n209), .B1(new_n202), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n211), .B(KEYINPUT89), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n216), .B(new_n217), .C1(new_n203), .C2(new_n202), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n214), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G8gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n221));
  INV_X1    g020(.A(G1gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n221), .B1(KEYINPUT91), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(KEYINPUT91), .B2(new_n222), .ZN(new_n224));
  INV_X1    g023(.A(G22gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G15gat), .ZN(new_n226));
  INV_X1    g025(.A(G15gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G22gat), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n226), .A2(new_n228), .A3(KEYINPUT90), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT90), .B1(new_n226), .B2(new_n228), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n224), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n220), .B1(new_n231), .B2(KEYINPUT92), .ZN(new_n232));
  INV_X1    g031(.A(new_n230), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n226), .A2(new_n228), .A3(KEYINPUT90), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n231), .B1(new_n235), .B2(G1gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  OAI221_X1 g036(.A(new_n231), .B1(KEYINPUT92), .B2(new_n220), .C1(new_n235), .C2(G1gat), .ZN(new_n238));
  AND3_X1   g037(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT93), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT93), .B1(new_n237), .B2(new_n238), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n219), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n219), .A2(KEYINPUT17), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT17), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n243), .B1(new_n214), .B2(new_n218), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n238), .B(new_n237), .C1(new_n242), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(G229gat), .A2(G233gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT94), .ZN(new_n248));
  INV_X1    g047(.A(new_n240), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT93), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n249), .A2(new_n250), .A3(new_n214), .A4(new_n218), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(new_n241), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n246), .B(KEYINPUT13), .Z(new_n253));
  AOI22_X1  g052(.A1(new_n248), .A2(KEYINPUT18), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(G197gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT11), .B(G169gat), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n256), .B(new_n257), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT12), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n247), .A2(KEYINPUT94), .A3(new_n260), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n254), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n259), .B1(new_n254), .B2(new_n261), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G227gat), .A2(G233gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n265), .B(KEYINPUT64), .Z(new_n266));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n267));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT24), .ZN(new_n270));
  NOR2_X1   g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  AOI22_X1  g070(.A1(new_n269), .A2(new_n270), .B1(new_n271), .B2(KEYINPUT23), .ZN(new_n272));
  INV_X1    g071(.A(G183gat), .ZN(new_n273));
  INV_X1    g072(.A(G190gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(KEYINPUT24), .A3(new_n268), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n271), .B2(KEYINPUT23), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n267), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n271), .A2(KEYINPUT23), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n281), .A2(new_n267), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n278), .B(KEYINPUT65), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n280), .B1(new_n277), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT27), .B(G183gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n274), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n269), .B1(new_n287), .B2(KEYINPUT28), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT26), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n289), .A2(KEYINPUT26), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n290), .B1(new_n291), .B2(new_n271), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n289), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n278), .A3(new_n293), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n273), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT27), .B1(new_n273), .B2(KEYINPUT66), .ZN(new_n296));
  NOR2_X1   g095(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n288), .B(new_n294), .C1(new_n295), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n285), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT69), .ZN(new_n301));
  XNOR2_X1  g100(.A(G127gat), .B(G134gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G134gat), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT68), .B1(new_n305), .B2(G127gat), .ZN(new_n306));
  INV_X1    g105(.A(G120gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(G113gat), .ZN(new_n308));
  INV_X1    g107(.A(G113gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G120gat), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI22_X1  g110(.A1(new_n304), .A2(new_n306), .B1(KEYINPUT1), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n311), .A2(KEYINPUT1), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n302), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n285), .A2(new_n316), .A3(new_n299), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n315), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n300), .A2(KEYINPUT69), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n266), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT71), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n266), .A3(new_n320), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT32), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT33), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G71gat), .B(G99gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT70), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(new_n227), .ZN(new_n329));
  INV_X1    g128(.A(G43gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n324), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n331), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n323), .B(KEYINPUT32), .C1(new_n325), .C2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT34), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n321), .B2(KEYINPUT71), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n332), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n332), .B2(new_n334), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n322), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n339), .ZN(new_n341));
  INV_X1    g140(.A(new_n322), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n342), .A3(new_n337), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT36), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n340), .A2(new_n343), .A3(KEYINPUT36), .ZN(new_n347));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT22), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT72), .B(G218gat), .ZN(new_n353));
  INV_X1    g152(.A(G211gat), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G197gat), .B(G204gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G211gat), .B(G218gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n300), .A2(new_n364), .B1(G226gat), .B2(G233gat), .ZN(new_n365));
  INV_X1    g164(.A(G226gat), .ZN(new_n366));
  INV_X1    g165(.A(G233gat), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n366), .B(new_n367), .C1(new_n285), .C2(new_n299), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n363), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n365), .A2(new_n368), .A3(new_n363), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n351), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OR3_X1    g171(.A1(new_n365), .A2(new_n368), .A3(new_n363), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(new_n369), .A3(new_n350), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(KEYINPUT30), .A3(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n373), .A2(new_n369), .A3(new_n376), .A4(new_n350), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(G225gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n315), .B(KEYINPUT74), .ZN(new_n383));
  AND2_X1   g182(.A1(G155gat), .A2(G162gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(G155gat), .A2(G162gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XOR2_X1   g185(.A(G141gat), .B(G148gat), .Z(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n387), .B2(KEYINPUT73), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT2), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n389), .B2(new_n384), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  OAI221_X1 g190(.A(new_n387), .B1(new_n389), .B2(new_n384), .C1(new_n386), .C2(KEYINPUT73), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n382), .B1(new_n383), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n315), .A2(KEYINPUT74), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT74), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n312), .B2(new_n314), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n382), .B(new_n393), .C1(new_n395), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n391), .A2(new_n392), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n319), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n381), .B1(new_n394), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT78), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(KEYINPUT78), .B(new_n381), .C1(new_n394), .C2(new_n401), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n391), .A2(KEYINPUT3), .A3(new_n392), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n407), .B(new_n408), .C1(new_n395), .C2(new_n397), .ZN(new_n409));
  XOR2_X1   g208(.A(KEYINPUT75), .B(KEYINPUT4), .Z(new_n410));
  NAND2_X1  g209(.A1(new_n400), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n319), .A2(KEYINPUT4), .A3(new_n399), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n409), .A2(new_n411), .A3(new_n380), .A4(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT76), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT5), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n413), .B2(new_n414), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n404), .A2(new_n405), .A3(new_n415), .A4(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n393), .B2(new_n315), .ZN(new_n420));
  INV_X1    g219(.A(new_n410), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n319), .A2(new_n399), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n423), .A2(new_n416), .A3(new_n380), .A4(new_n409), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G1gat), .B(G29gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT0), .ZN(new_n427));
  XNOR2_X1  g226(.A(G57gat), .B(G85gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n418), .A2(new_n429), .A3(new_n424), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI211_X1 g233(.A(new_n432), .B(new_n429), .C1(new_n418), .C2(new_n424), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n379), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT29), .B1(new_n360), .B2(new_n361), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n439), .A2(KEYINPUT3), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT29), .B1(new_n399), .B2(new_n406), .ZN(new_n441));
  OAI22_X1  g240(.A1(new_n440), .A2(new_n399), .B1(new_n362), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(G228gat), .A2(G233gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n363), .B1(new_n441), .B2(KEYINPUT81), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT82), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(KEYINPUT81), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n448), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT82), .B1(new_n450), .B2(new_n445), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n362), .A2(new_n364), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n406), .B1(new_n439), .B2(KEYINPUT80), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n393), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(G228gat), .A3(G233gat), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n444), .B1(new_n452), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n438), .B1(new_n459), .B2(G22gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(G78gat), .B(G106gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n461), .B(KEYINPUT79), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT31), .ZN(new_n463));
  INV_X1    g262(.A(G50gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n458), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n451), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n469), .A2(new_n225), .A3(new_n444), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n225), .B1(new_n469), .B2(new_n444), .ZN(new_n471));
  OAI22_X1  g270(.A1(new_n460), .A2(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n471), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n469), .A2(new_n225), .A3(new_n444), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n438), .A4(new_n465), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n346), .B(new_n347), .C1(new_n437), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT84), .ZN(new_n478));
  INV_X1    g277(.A(new_n347), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT36), .B1(new_n340), .B2(new_n343), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n433), .A2(new_n432), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n429), .B1(new_n418), .B2(new_n424), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n378), .B1(new_n484), .B2(new_n435), .ZN(new_n485));
  INV_X1    g284(.A(new_n476), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n481), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT37), .B1(new_n370), .B2(new_n371), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT37), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n373), .A2(new_n369), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n351), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT38), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n374), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n493), .A2(KEYINPUT38), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n434), .A3(new_n436), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n380), .B1(new_n423), .B2(new_n409), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT39), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n430), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n409), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n420), .A2(new_n422), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n381), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n393), .B1(new_n395), .B2(new_n397), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT77), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n506), .A2(new_n380), .A3(new_n400), .A4(new_n398), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT39), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n501), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT40), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n501), .A2(new_n508), .A3(KEYINPUT40), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n511), .A2(new_n377), .A3(new_n375), .A4(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT85), .B1(new_n513), .B2(new_n483), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n501), .A2(new_n508), .A3(KEYINPUT40), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT40), .B1(new_n501), .B2(new_n508), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT85), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n431), .A2(new_n379), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n498), .A2(new_n520), .A3(new_n476), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n478), .A2(new_n489), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT86), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n476), .A2(new_n344), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT35), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n476), .A2(new_n344), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n525), .B(new_n526), .C1(new_n527), .C2(new_n485), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n475), .A2(new_n472), .B1(new_n340), .B2(new_n343), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n529), .B(new_n437), .C1(new_n524), .C2(KEYINPUT35), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n264), .B1(new_n523), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n434), .A2(new_n436), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G71gat), .A2(G78gat), .ZN(new_n536));
  INV_X1    g335(.A(G71gat), .ZN(new_n537));
  INV_X1    g336(.A(G78gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT9), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n536), .B(new_n539), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G57gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(G64gat), .ZN(new_n544));
  INV_X1    g343(.A(G64gat), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(G57gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n539), .A2(new_n536), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n536), .A2(new_n541), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n542), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT95), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n542), .A2(KEYINPUT95), .A3(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT21), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G127gat), .B(G155gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT20), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G183gat), .B(G211gat), .Z(new_n564));
  NOR2_X1   g363(.A1(new_n559), .A2(new_n561), .ZN(new_n565));
  OR3_X1    g364(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n249), .B(new_n250), .C1(new_n556), .C2(new_n555), .ZN(new_n569));
  XNOR2_X1  g368(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n571), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(KEYINPUT98), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n578));
  AND2_X1   g377(.A1(G99gat), .A2(G106gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G92gat), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n583), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n584));
  NAND2_X1  g383(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(G92gat), .ZN(new_n586));
  NOR2_X1   g385(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n576), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(KEYINPUT97), .A2(G99gat), .A3(G106gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(KEYINPUT8), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n582), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n581), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n595), .A2(new_n592), .A3(new_n588), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n594), .A2(KEYINPUT99), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n593), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(KEYINPUT100), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n599), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT100), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n600), .B(new_n603), .C1(new_n242), .C2(new_n244), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n597), .A2(KEYINPUT100), .A3(new_n599), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT100), .B1(new_n597), .B2(new_n599), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n219), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n604), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G190gat), .B(G218gat), .Z(new_n610));
  AND2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n609), .A2(new_n610), .ZN(new_n612));
  XNOR2_X1  g411(.A(G134gat), .B(G162gat), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  OR3_X1    g415(.A1(new_n611), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n616), .B1(new_n611), .B2(new_n612), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n574), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G230gat), .A2(G233gat), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT7), .ZN(new_n623));
  INV_X1    g422(.A(G85gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(G92gat), .A3(new_n585), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT8), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(new_n576), .B2(new_n589), .ZN(new_n628));
  AOI22_X1  g427(.A1(new_n626), .A2(new_n584), .B1(new_n628), .B2(new_n591), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n542), .B(new_n550), .C1(new_n629), .C2(new_n595), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n582), .A2(new_n593), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT101), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n551), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n633), .A2(new_n594), .A3(new_n634), .A4(new_n596), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT10), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n555), .A2(new_n599), .A3(new_n597), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n553), .A2(KEYINPUT10), .A3(new_n554), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n640), .B1(new_n603), .B2(new_n600), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n622), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n622), .B1(new_n636), .B2(new_n638), .ZN(new_n644));
  XOR2_X1   g443(.A(G120gat), .B(G148gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT102), .ZN(new_n646));
  XNOR2_X1  g445(.A(G176gat), .B(G204gat), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n646), .B(new_n647), .Z(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n622), .B(KEYINPUT103), .Z(new_n653));
  INV_X1    g452(.A(new_n640), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(new_n605), .B2(new_n606), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n653), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n649), .B1(new_n657), .B2(new_n644), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n621), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n533), .A2(new_n535), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(G1gat), .ZN(G1324gat));
  INV_X1    g463(.A(new_n533), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(new_n378), .A3(new_n661), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT16), .B(G8gat), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(new_n220), .B2(new_n666), .ZN(new_n669));
  MUX2_X1   g468(.A(new_n668), .B(new_n669), .S(KEYINPUT42), .Z(G1325gat));
  NAND4_X1  g469(.A1(new_n533), .A2(new_n227), .A3(new_n344), .A4(new_n662), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n665), .A2(new_n481), .A3(new_n661), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n672), .B2(new_n227), .ZN(G1326gat));
  NOR2_X1   g472(.A1(new_n665), .A2(new_n661), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n674), .A2(new_n486), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT104), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n677), .A3(new_n486), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n679), .B(new_n681), .ZN(G1327gat));
  INV_X1    g481(.A(new_n574), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n683), .A2(new_n619), .A3(new_n659), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n533), .A2(new_n684), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n685), .A2(G29gat), .A3(new_n534), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT45), .Z(new_n687));
  NAND2_X1  g486(.A1(new_n523), .A2(new_n532), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n619), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n528), .B(new_n530), .C1(new_n477), .C2(new_n521), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n620), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n689), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n574), .B(KEYINPUT105), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n696), .A2(new_n264), .A3(new_n659), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(G29gat), .B1(new_n698), .B2(new_n534), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n687), .A2(new_n699), .ZN(G1328gat));
  NOR3_X1   g499(.A1(new_n685), .A2(G36gat), .A3(new_n378), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT46), .ZN(new_n702));
  OAI21_X1  g501(.A(G36gat), .B1(new_n698), .B2(new_n378), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(G1329gat));
  OAI21_X1  g503(.A(G43gat), .B1(new_n698), .B2(new_n481), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n533), .A2(new_n330), .A3(new_n344), .A4(new_n684), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1330gat));
  INV_X1    g511(.A(KEYINPUT48), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n691), .A2(new_n694), .A3(new_n486), .A4(new_n697), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G50gat), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n715), .B2(KEYINPUT107), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n685), .A2(G50gat), .A3(new_n476), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n717), .B1(G50gat), .B2(new_n714), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n716), .B(new_n718), .ZN(G1331gat));
  INV_X1    g518(.A(new_n264), .ZN(new_n720));
  NOR4_X1   g519(.A1(new_n574), .A2(new_n720), .A3(new_n620), .A4(new_n660), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n692), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n692), .A2(KEYINPUT108), .A3(new_n721), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n534), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(new_n543), .ZN(G1332gat));
  XNOR2_X1  g527(.A(KEYINPUT109), .B(KEYINPUT110), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n726), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n378), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n733), .A2(new_n734), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n730), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n737), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n739), .A2(new_n729), .A3(new_n735), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(G1333gat));
  NAND2_X1  g540(.A1(new_n346), .A2(new_n347), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n731), .A2(G71gat), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n744));
  INV_X1    g543(.A(new_n344), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n726), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n537), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n726), .A2(new_n744), .A3(new_n745), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n743), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT50), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n751), .B(new_n743), .C1(new_n747), .C2(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1334gat));
  NOR2_X1   g552(.A1(new_n726), .A2(new_n476), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(new_n538), .ZN(G1335gat));
  NOR3_X1   g554(.A1(new_n683), .A2(new_n720), .A3(new_n660), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n691), .A2(new_n694), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758), .B2(new_n534), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n683), .A2(new_n720), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n692), .A2(new_n620), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n692), .A2(KEYINPUT51), .A3(new_n620), .A4(new_n760), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n535), .A2(new_n624), .A3(new_n659), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n759), .B1(new_n766), .B2(new_n767), .ZN(G1336gat));
  NAND2_X1  g567(.A1(new_n757), .A2(new_n379), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n660), .A2(G92gat), .A3(new_n378), .ZN(new_n770));
  AOI22_X1  g569(.A1(new_n769), .A2(G92gat), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1337gat));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n481), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT112), .B(G99gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n344), .A2(new_n659), .A3(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT113), .ZN(new_n777));
  OAI22_X1  g576(.A1(new_n774), .A2(new_n775), .B1(new_n766), .B2(new_n777), .ZN(G1338gat));
  NAND4_X1  g577(.A1(new_n691), .A2(new_n694), .A3(new_n486), .A4(new_n756), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(G106gat), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n476), .A2(G106gat), .A3(new_n660), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT53), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(KEYINPUT114), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n765), .A2(new_n787), .A3(new_n781), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n779), .B2(G106gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n785), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n787), .B1(new_n765), .B2(new_n781), .ZN(new_n793));
  INV_X1    g592(.A(new_n781), .ZN(new_n794));
  AOI211_X1 g593(.A(KEYINPUT114), .B(new_n794), .C1(new_n763), .C2(new_n764), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n791), .B(new_n785), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n784), .B1(new_n792), .B2(new_n797), .ZN(G1339gat));
  NAND2_X1  g597(.A1(new_n535), .A2(new_n378), .ZN(new_n799));
  INV_X1    g598(.A(new_n696), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT54), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n648), .B1(new_n657), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n655), .A2(new_n656), .A3(new_n653), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n642), .A2(KEYINPUT54), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n655), .A2(new_n656), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n801), .B1(new_n808), .B2(new_n622), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(KEYINPUT117), .A3(new_n804), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n803), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT118), .B1(new_n811), .B2(KEYINPUT55), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n651), .B1(new_n811), .B2(KEYINPUT55), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n809), .A2(KEYINPUT117), .A3(new_n804), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT117), .B1(new_n809), .B2(new_n804), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n802), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n812), .A2(new_n813), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n812), .A2(new_n813), .A3(new_n819), .A4(KEYINPUT119), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n720), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n254), .A2(new_n259), .A3(new_n261), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n252), .A2(new_n253), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n246), .B1(new_n241), .B2(new_n245), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n258), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n659), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n620), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n620), .A2(new_n825), .A3(new_n828), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n822), .A2(new_n831), .A3(new_n823), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n800), .B1(new_n830), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n661), .A2(new_n720), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  AOI211_X1 g635(.A(new_n486), .B(new_n799), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n344), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(new_n309), .A3(new_n264), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n534), .B1(new_n834), .B2(new_n836), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n529), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n378), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n720), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n839), .B1(new_n843), .B2(new_n309), .ZN(G1340gat));
  AOI21_X1  g643(.A(G120gat), .B1(new_n842), .B2(new_n659), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n745), .A2(new_n307), .A3(new_n660), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n837), .B2(new_n846), .ZN(G1341gat));
  INV_X1    g646(.A(G127gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n842), .A2(new_n848), .A3(new_n683), .ZN(new_n849));
  OAI21_X1  g648(.A(G127gat), .B1(new_n838), .B2(new_n800), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1342gat));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n620), .A2(new_n378), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(G134gat), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n841), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT120), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n855), .A2(KEYINPUT120), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n852), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(G134gat), .B1(new_n838), .B2(new_n619), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n855), .A2(KEYINPUT120), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(KEYINPUT56), .A3(new_n856), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(G1343gat));
  NAND2_X1  g662(.A1(new_n829), .A2(KEYINPUT121), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n825), .A2(new_n659), .A3(new_n865), .A4(new_n828), .ZN(new_n866));
  XOR2_X1   g665(.A(KEYINPUT122), .B(KEYINPUT55), .Z(new_n867));
  OAI22_X1  g666(.A1(new_n262), .A2(new_n263), .B1(new_n811), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n652), .B1(new_n816), .B2(new_n818), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n864), .B(new_n866), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n619), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n832), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(KEYINPUT123), .A3(new_n574), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n836), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT123), .B1(new_n872), .B2(new_n574), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n486), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT57), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n476), .B1(new_n834), .B2(new_n836), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n799), .A2(new_n742), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n877), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G141gat), .B1(new_n882), .B2(new_n264), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n742), .A2(new_n476), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n840), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n379), .ZN(new_n886));
  INV_X1    g685(.A(G141gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n720), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n890), .B1(new_n888), .B2(KEYINPUT124), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n883), .B(new_n888), .C1(KEYINPUT124), .C2(new_n890), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(G1344gat));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n880), .A3(new_n659), .A4(new_n881), .ZN(new_n895));
  INV_X1    g694(.A(G148gat), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(KEYINPUT59), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n831), .A2(new_n819), .A3(new_n813), .A4(new_n812), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n683), .B1(new_n871), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n879), .B(new_n486), .C1(new_n899), .C2(new_n835), .ZN(new_n900));
  NOR3_X1   g699(.A1(new_n799), .A2(new_n742), .A3(new_n660), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n900), .B(new_n901), .C1(new_n878), .C2(new_n879), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G148gat), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n895), .A2(new_n897), .B1(new_n903), .B2(KEYINPUT59), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n896), .A3(new_n659), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT125), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n895), .A2(new_n897), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT59), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n902), .B2(G148gat), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n908), .B(new_n905), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n907), .A2(new_n912), .ZN(G1345gat));
  OAI21_X1  g712(.A(G155gat), .B1(new_n882), .B2(new_n800), .ZN(new_n914));
  INV_X1    g713(.A(G155gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n886), .A2(new_n915), .A3(new_n683), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1346gat));
  OAI21_X1  g716(.A(G162gat), .B1(new_n882), .B2(new_n619), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n853), .A2(G162gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n885), .B2(new_n919), .ZN(G1347gat));
  AOI21_X1  g719(.A(new_n486), .B1(new_n834), .B2(new_n836), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n534), .A2(new_n379), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n745), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(G169gat), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n924), .A2(new_n925), .A3(new_n264), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n535), .B1(new_n834), .B2(new_n836), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(new_n379), .A3(new_n529), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n720), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n926), .B1(new_n925), .B2(new_n929), .ZN(G1348gat));
  INV_X1    g729(.A(G176gat), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n924), .A2(new_n931), .A3(new_n660), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n659), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n931), .B2(new_n933), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n286), .A3(new_n683), .ZN(new_n935));
  OAI21_X1  g734(.A(G183gat), .B1(new_n924), .B2(new_n800), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g737(.A1(new_n921), .A2(new_n620), .A3(new_n923), .ZN(new_n939));
  AND2_X1   g738(.A1(new_n939), .A2(G190gat), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n940), .A2(KEYINPUT126), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(KEYINPUT126), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(KEYINPUT61), .A3(new_n942), .ZN(new_n943));
  OR3_X1    g742(.A1(new_n940), .A2(KEYINPUT126), .A3(KEYINPUT61), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n928), .A2(new_n274), .A3(new_n620), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(G1351gat));
  NOR3_X1   g745(.A1(new_n742), .A2(new_n378), .A3(new_n476), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n927), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  XNOR2_X1  g748(.A(KEYINPUT127), .B(G197gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n949), .A2(new_n720), .A3(new_n950), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n878), .A2(new_n879), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n742), .A2(new_n922), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n900), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(new_n264), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n951), .B1(new_n955), .B2(new_n950), .ZN(G1352gat));
  OR3_X1    g755(.A1(new_n948), .A2(G204gat), .A3(new_n660), .ZN(new_n957));
  OR2_X1    g756(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n958));
  OAI21_X1  g757(.A(G204gat), .B1(new_n954), .B2(new_n660), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(G1353gat));
  NAND3_X1  g760(.A1(new_n949), .A2(new_n354), .A3(new_n683), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n952), .A2(new_n683), .A3(new_n900), .A4(new_n953), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n963), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G1354gat));
  OR2_X1    g766(.A1(new_n619), .A2(new_n353), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n948), .A2(new_n619), .ZN(new_n969));
  OAI22_X1  g768(.A1(new_n954), .A2(new_n968), .B1(G218gat), .B2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(G1355gat));
endmodule


