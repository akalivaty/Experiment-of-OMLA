//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT0), .A3(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G125), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G128), .Z(new_n200));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(G143), .B2(new_n187), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n191), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G125), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n195), .A2(new_n201), .A3(G128), .ZN(new_n205));
  AND3_X1   g019(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n199), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G953), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G224), .ZN(new_n209));
  XOR2_X1   g023(.A(new_n209), .B(KEYINPUT92), .Z(new_n210));
  XNOR2_X1  g024(.A(new_n207), .B(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT70), .ZN(new_n212));
  NAND2_X1  g026(.A1(KEYINPUT2), .A2(G113), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n215));
  INV_X1    g029(.A(G113), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT67), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT67), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(KEYINPUT2), .B2(G113), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n214), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(KEYINPUT69), .A2(G116), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT69), .A2(G116), .ZN(new_n222));
  INV_X1    g036(.A(G119), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G116), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(G119), .ZN(new_n226));
  OAI22_X1  g040(.A1(new_n220), .A2(KEYINPUT68), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n228));
  AOI211_X1 g042(.A(new_n228), .B(new_n214), .C1(new_n217), .C2(new_n219), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n212), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n224), .A2(new_n226), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n220), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n218), .A2(KEYINPUT2), .A3(G113), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT67), .B1(new_n215), .B2(new_n216), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n213), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n228), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n220), .A2(KEYINPUT68), .ZN(new_n237));
  INV_X1    g051(.A(new_n222), .ZN(new_n238));
  NAND2_X1  g052(.A1(KEYINPUT69), .A2(G116), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(G119), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n226), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n236), .A2(KEYINPUT70), .A3(new_n237), .A4(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n230), .A2(new_n232), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G104), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT3), .B1(new_n245), .B2(G107), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g061(.A(G107), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(G104), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(G107), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n246), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n246), .A2(new_n249), .A3(KEYINPUT80), .A4(new_n250), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n253), .A2(new_n254), .A3(G101), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(KEYINPUT82), .ZN(new_n257));
  INV_X1    g071(.A(G101), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n251), .B2(new_n252), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT82), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n259), .A2(new_n260), .A3(new_n254), .A4(new_n255), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n253), .A2(G101), .A3(new_n255), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n246), .A2(new_n249), .A3(new_n258), .A4(new_n250), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n264), .A2(KEYINPUT4), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT81), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AND3_X1   g080(.A1(new_n263), .A2(KEYINPUT81), .A3(new_n265), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n244), .B(new_n262), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT83), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n248), .A3(G104), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT83), .B1(new_n245), .B2(G107), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n248), .A2(G104), .ZN(new_n272));
  OAI211_X1 g086(.A(G101), .B(new_n270), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(new_n264), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT86), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n240), .A2(KEYINPUT5), .A3(new_n241), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n216), .B1(new_n226), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n264), .A3(KEYINPUT86), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n276), .A2(new_n280), .A3(new_n232), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT90), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n277), .A2(new_n279), .B1(new_n231), .B2(new_n220), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT90), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n276), .A4(new_n281), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n268), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT91), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT91), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n268), .A2(new_n291), .A3(new_n287), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G122), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n289), .A2(new_n290), .A3(new_n292), .A4(new_n294), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n268), .A2(new_n291), .A3(new_n287), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n291), .B1(new_n268), .B2(new_n287), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n296), .A2(new_n297), .A3(new_n293), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n268), .A2(new_n287), .A3(new_n293), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT6), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n211), .B(new_n295), .C1(new_n298), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n209), .A2(KEYINPUT7), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n302), .B1(new_n199), .B2(new_n206), .ZN(new_n303));
  INV_X1    g117(.A(new_n302), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n203), .A2(new_n205), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n198), .B(new_n304), .C1(G125), .C2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(new_n293), .B(KEYINPUT8), .Z(new_n308));
  NAND2_X1  g122(.A1(new_n280), .A2(new_n232), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n274), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n308), .B1(new_n310), .B2(new_n282), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n299), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT93), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT93), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n317), .A3(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G210), .B1(G237), .B2(G902), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n301), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n320), .B1(new_n301), .B2(new_n319), .ZN(new_n322));
  OR3_X1    g136(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT94), .ZN(new_n323));
  OAI21_X1  g137(.A(G214), .B1(G237), .B2(G902), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(KEYINPUT94), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n238), .A2(G122), .A3(new_n239), .ZN(new_n327));
  OR2_X1    g141(.A1(new_n225), .A2(G122), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n248), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n200), .A2(G143), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n189), .A2(G128), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT64), .B(G134), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n331), .B2(new_n332), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT14), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(G107), .B1(new_n327), .B2(new_n336), .ZN(new_n338));
  OAI221_X1 g152(.A(new_n330), .B1(new_n334), .B2(new_n335), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n334), .ZN(new_n340));
  INV_X1    g154(.A(new_n331), .ZN(new_n341));
  XOR2_X1   g155(.A(new_n332), .B(KEYINPUT13), .Z(new_n342));
  OAI21_X1  g156(.A(G134), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n330), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n329), .A2(new_n248), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n340), .B(new_n343), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT9), .B(G234), .ZN(new_n347));
  INV_X1    g161(.A(G217), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n347), .A2(new_n348), .A3(G953), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n339), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT99), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n339), .A2(new_n346), .ZN(new_n353));
  INV_X1    g167(.A(new_n349), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n339), .A2(KEYINPUT99), .A3(new_n346), .A4(new_n349), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n352), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n314), .ZN(new_n358));
  INV_X1    g172(.A(G478), .ZN(new_n359));
  OR2_X1    g173(.A1(new_n359), .A2(KEYINPUT15), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n358), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n208), .A3(G214), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT95), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(new_n189), .ZN(new_n366));
  NOR2_X1   g180(.A1(G237), .A2(G953), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n367), .B(G214), .C1(KEYINPUT95), .C2(G143), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  AND2_X1   g183(.A1(KEYINPUT18), .A2(G131), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(KEYINPUT96), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n370), .ZN(new_n373));
  XNOR2_X1  g187(.A(G125), .B(G140), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n374), .A2(new_n187), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n374), .A2(new_n187), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n372), .B(new_n373), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G113), .B(G122), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(new_n245), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n374), .A2(KEYINPUT16), .ZN(new_n380));
  OR3_X1    g194(.A1(new_n204), .A2(KEYINPUT16), .A3(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n187), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(G146), .A3(new_n381), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n369), .A2(KEYINPUT17), .A3(G131), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n369), .B(G131), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n385), .B(new_n386), .C1(KEYINPUT17), .C2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n377), .A2(new_n379), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n379), .B1(new_n377), .B2(new_n388), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n314), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G475), .ZN(new_n393));
  NAND2_X1  g207(.A1(G234), .A2(G237), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(G952), .A3(new_n208), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(G902), .A3(G953), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT21), .B(G898), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT97), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n374), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(KEYINPUT19), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n387), .B(new_n384), .C1(G146), .C2(new_n404), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n377), .A2(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n389), .B1(new_n406), .B2(new_n379), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT20), .ZN(new_n408));
  NOR2_X1   g222(.A1(G475), .A2(G902), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(KEYINPUT98), .Z(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n408), .B1(new_n407), .B2(new_n410), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n393), .B(new_n401), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(KEYINPUT100), .B1(new_n362), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n413), .ZN(new_n416));
  AOI22_X1  g230(.A1(new_n416), .A2(new_n411), .B1(G475), .B2(new_n392), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT100), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n417), .A2(new_n361), .A3(new_n418), .A4(new_n401), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n326), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT71), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT11), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n333), .B2(G137), .ZN(new_n425));
  INV_X1    g239(.A(G137), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n426), .A2(G134), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n427), .B1(new_n333), .B2(G137), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n425), .B1(new_n428), .B2(new_n424), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G131), .ZN(new_n430));
  INV_X1    g244(.A(G131), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n431), .B(new_n425), .C1(new_n428), .C2(new_n424), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n197), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n333), .A2(G137), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n426), .A2(G134), .ZN(new_n435));
  OAI21_X1  g249(.A(G131), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n305), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n433), .A2(new_n244), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n423), .B1(new_n439), .B2(KEYINPUT28), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT28), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n430), .A2(new_n432), .ZN(new_n442));
  INV_X1    g256(.A(new_n197), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n437), .ZN(new_n445));
  OAI211_X1 g259(.A(KEYINPUT71), .B(new_n441), .C1(new_n445), .C2(new_n244), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n439), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n445), .A2(new_n244), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n447), .B1(KEYINPUT28), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n367), .A2(G210), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n452), .B(KEYINPUT27), .Z(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT26), .B(G101), .ZN(new_n454));
  XOR2_X1   g268(.A(new_n453), .B(new_n454), .Z(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT29), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(G902), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n444), .A2(KEYINPUT30), .A3(new_n437), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT65), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n433), .A2(new_n462), .ZN(new_n463));
  AOI211_X1 g277(.A(KEYINPUT65), .B(new_n197), .C1(new_n430), .C2(new_n432), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n437), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT30), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n439), .B1(new_n467), .B2(new_n244), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n457), .B1(new_n468), .B2(new_n455), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n244), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n441), .B1(new_n470), .B2(new_n448), .ZN(new_n471));
  NOR3_X1   g285(.A1(new_n471), .A2(new_n447), .A3(new_n456), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n459), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G472), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n444), .A2(KEYINPUT65), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n433), .A2(new_n462), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n438), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n244), .B(new_n460), .C1(new_n477), .C2(KEYINPUT30), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n448), .A3(new_n455), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT31), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n456), .B1(new_n471), .B2(new_n447), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT31), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n478), .A2(new_n482), .A3(new_n448), .A4(new_n455), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT32), .ZN(new_n485));
  NOR2_X1   g299(.A1(G472), .A2(G902), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n485), .B1(new_n484), .B2(new_n486), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n474), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G221), .B1(new_n347), .B2(G902), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(KEYINPUT79), .ZN(new_n491));
  INV_X1    g305(.A(G469), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n305), .B1(new_n276), .B2(new_n281), .ZN(new_n493));
  INV_X1    g307(.A(G128), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT84), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n494), .B1(new_n202), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT84), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n191), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n274), .B1(new_n500), .B2(new_n205), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n442), .B1(new_n493), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT12), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT88), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT88), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n502), .A2(new_n506), .A3(new_n503), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n442), .B(KEYINPUT12), .C1(new_n493), .C2(new_n501), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(KEYINPUT87), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n510), .A3(KEYINPUT89), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT89), .B1(new_n508), .B2(new_n510), .ZN(new_n513));
  AND4_X1   g327(.A1(KEYINPUT10), .A2(new_n276), .A3(new_n305), .A4(new_n281), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT85), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n515), .B1(new_n501), .B2(KEYINPUT10), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT10), .ZN(new_n517));
  INV_X1    g331(.A(new_n205), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n499), .B2(new_n191), .ZN(new_n519));
  OAI211_X1 g333(.A(KEYINPUT85), .B(new_n517), .C1(new_n519), .C2(new_n274), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n514), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n262), .B(new_n443), .C1(new_n266), .C2(new_n267), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n521), .A2(new_n432), .A3(new_n430), .A4(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(G110), .B(G140), .ZN(new_n524));
  INV_X1    g338(.A(G227), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(G953), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n524), .B(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n512), .A2(new_n513), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n521), .A2(new_n522), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n442), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n523), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n527), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n492), .B(new_n314), .C1(new_n530), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n508), .A2(new_n510), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n528), .B1(new_n537), .B2(new_n523), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n533), .A2(new_n527), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(G469), .B1(new_n540), .B2(G902), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n491), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n348), .B1(G234), .B2(new_n314), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT76), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n545));
  AOI21_X1  g359(.A(G902), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G110), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT23), .B1(new_n494), .B2(G119), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n494), .A2(G119), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n200), .A2(G119), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT23), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n548), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT72), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT66), .B(G128), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(new_n223), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT23), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT72), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n558), .A2(new_n559), .A3(new_n548), .A4(new_n551), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT73), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n557), .A2(new_n550), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT24), .B(G110), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n561), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(KEYINPUT73), .B(new_n563), .C1(new_n557), .C2(new_n550), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n555), .A2(new_n560), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n384), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(new_n375), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n383), .A2(new_n384), .B1(new_n562), .B2(new_n564), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n558), .A2(new_n551), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G110), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT22), .B(G137), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n208), .A2(G221), .A3(G234), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n570), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT75), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n567), .A2(new_n569), .B1(new_n571), .B2(new_n573), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n577), .B(KEYINPUT74), .Z(new_n581));
  OAI211_X1 g395(.A(new_n578), .B(new_n579), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(KEYINPUT75), .A3(new_n577), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n547), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n544), .A2(new_n545), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n543), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  AOI211_X1 g401(.A(new_n585), .B(new_n547), .C1(new_n582), .C2(new_n583), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n582), .A2(new_n583), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n543), .A2(G902), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT77), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT77), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n594), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT78), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n589), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n582), .A2(new_n583), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n585), .B1(new_n599), .B2(new_n547), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n584), .A2(new_n586), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n601), .A3(new_n543), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n590), .A2(new_n594), .A3(new_n591), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n594), .B1(new_n590), .B2(new_n591), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT78), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n598), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n422), .A2(new_n489), .A3(new_n542), .A4(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(G101), .ZN(G3));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n610));
  INV_X1    g424(.A(G472), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n484), .B2(new_n314), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n484), .A2(new_n486), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n610), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n612), .A2(KEYINPUT101), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(new_n542), .A3(new_n607), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n324), .B1(new_n321), .B2(new_n322), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT102), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n621), .B(new_n324), .C1(new_n321), .C2(new_n322), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n393), .B1(new_n412), .B2(new_n413), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n358), .A2(new_n359), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n357), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n355), .A2(KEYINPUT33), .A3(new_n350), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n359), .A2(G902), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n624), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n400), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n620), .A2(new_n622), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT103), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n620), .A2(KEYINPUT103), .A3(new_n622), .A4(new_n633), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n618), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  XOR2_X1   g454(.A(new_n400), .B(KEYINPUT104), .Z(new_n641));
  NOR2_X1   g455(.A1(new_n623), .A2(new_n361), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n620), .A2(new_n622), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n618), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT35), .B(G107), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  INV_X1    g460(.A(KEYINPUT36), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n581), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n580), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n591), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n602), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n422), .A2(new_n617), .A3(new_n542), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n398), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n395), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n623), .A2(new_n361), .A3(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n489), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n620), .A2(new_n622), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n542), .A2(new_n651), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XNOR2_X1  g478(.A(new_n657), .B(KEYINPUT39), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n542), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(KEYINPUT40), .ZN(new_n668));
  INV_X1    g482(.A(new_n651), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n417), .A2(new_n361), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n324), .A3(new_n670), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n667), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n323), .A2(new_n325), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT38), .Z(new_n674));
  NOR2_X1   g488(.A1(new_n468), .A2(new_n456), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n314), .B1(new_n450), .B2(new_n455), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n487), .B2(new_n488), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT105), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n614), .A2(KEYINPUT32), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n683), .A3(new_n677), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n672), .A2(new_n674), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G143), .ZN(G45));
  NOR2_X1   g501(.A1(new_n632), .A2(new_n658), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n682), .B2(new_n474), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n661), .A3(new_n662), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n636), .A2(new_n637), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT89), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n529), .B1(new_n537), .B2(new_n695), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n696), .A2(new_n511), .B1(new_n533), .B2(new_n527), .ZN(new_n697));
  OAI21_X1  g511(.A(G469), .B1(new_n697), .B2(G902), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n698), .A2(new_n490), .A3(new_n536), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n489), .A2(new_n607), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n693), .B1(new_n694), .B2(new_n701), .ZN(new_n702));
  AOI211_X1 g516(.A(KEYINPUT106), .B(new_n700), .C1(new_n636), .C2(new_n637), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT41), .B(G113), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  OR2_X1    g520(.A1(new_n700), .A2(new_n643), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  NAND3_X1  g522(.A1(new_n489), .A2(new_n420), .A3(new_n651), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n699), .A2(new_n620), .A3(new_n622), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G119), .ZN(G21));
  NAND3_X1  g526(.A1(new_n620), .A2(new_n622), .A3(new_n670), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n699), .A2(new_n641), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n589), .A2(new_n596), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n480), .B(new_n483), .C1(new_n455), .C2(new_n451), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n486), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n613), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n713), .A2(new_n714), .A3(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n719), .B(G122), .Z(G24));
  AND4_X1   g534(.A1(new_n613), .A2(new_n688), .A3(new_n651), .A4(new_n717), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n661), .A2(new_n721), .A3(new_n699), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  INV_X1    g537(.A(new_n324), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n323), .B2(new_n325), .ZN(new_n725));
  INV_X1    g539(.A(new_n490), .ZN(new_n726));
  NAND2_X1  g540(.A1(G469), .A2(G902), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT107), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n696), .A2(new_n511), .ZN(new_n730));
  AOI21_X1  g544(.A(G902), .B1(new_n730), .B2(new_n534), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n729), .B1(new_n731), .B2(new_n492), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n538), .A2(KEYINPUT108), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT108), .B1(new_n538), .B2(new_n539), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(G469), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n726), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n725), .A2(new_n688), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n489), .A2(new_n715), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT42), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n489), .A2(new_n607), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n689), .A2(KEYINPUT42), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n725), .A3(new_n736), .A4(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n739), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n431), .ZN(G33));
  NAND4_X1  g559(.A1(new_n741), .A2(new_n659), .A3(new_n725), .A4(new_n736), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G134), .ZN(G36));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(new_n623), .B2(KEYINPUT109), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n417), .A2(new_n631), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n617), .A2(new_n669), .A3(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(KEYINPUT44), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n540), .A2(KEYINPUT45), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n492), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n733), .A2(new_n734), .A3(KEYINPUT45), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n729), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n757), .A2(KEYINPUT46), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n536), .B1(new_n757), .B2(KEYINPUT46), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n490), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n665), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n753), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n752), .A2(KEYINPUT44), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n763), .A2(KEYINPUT110), .A3(new_n725), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT110), .B1(new_n763), .B2(new_n725), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n762), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  OR3_X1    g581(.A1(new_n489), .A2(new_n607), .A3(new_n689), .ZN(new_n768));
  INV_X1    g582(.A(new_n725), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n760), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n771), .A2(KEYINPUT47), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(KEYINPUT47), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(G140), .Z(G42));
  NAND2_X1  g589(.A1(new_n698), .A2(new_n536), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT111), .ZN(new_n777));
  XOR2_X1   g591(.A(new_n777), .B(KEYINPUT49), .Z(new_n778));
  INV_X1    g592(.A(new_n674), .ZN(new_n779));
  INV_X1    g593(.A(new_n685), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n750), .A2(new_n724), .A3(new_n491), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(new_n715), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n778), .A2(new_n779), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  OAI22_X1  g597(.A1(new_n643), .A2(new_n700), .B1(new_n709), .B2(new_n710), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(new_n719), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(new_n702), .B2(new_n703), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(KEYINPUT112), .ZN(new_n787));
  INV_X1    g601(.A(new_n632), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n641), .B1(new_n788), .B2(new_n642), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n326), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n617), .A3(new_n542), .A4(new_n607), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n652), .A2(new_n791), .A3(new_n608), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n613), .A2(new_n651), .A3(new_n717), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n725), .A2(new_n793), .A3(new_n688), .A4(new_n736), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n669), .A2(new_n362), .A3(new_n623), .A4(new_n658), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n725), .A2(new_n795), .A3(new_n489), .A4(new_n542), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n746), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n792), .A2(new_n744), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n799), .B(new_n785), .C1(new_n702), .C2(new_n703), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n663), .A2(new_n691), .A3(new_n722), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n657), .B(KEYINPUT113), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n650), .B(new_n803), .C1(new_n587), .C2(new_n588), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT114), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n736), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n713), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n685), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n801), .B1(new_n802), .B2(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n661), .B(new_n662), .C1(new_n660), .C2(new_n690), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n685), .A2(new_n806), .A3(new_n807), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT52), .A4(new_n722), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n787), .A2(new_n798), .A3(new_n800), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n792), .A2(new_n744), .A3(new_n797), .A4(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n786), .B1(new_n809), .B2(new_n812), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n814), .A2(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n816), .A2(new_n787), .A3(new_n800), .A4(new_n813), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(KEYINPUT115), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n814), .A2(new_n815), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n822), .B1(new_n825), .B2(new_n821), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n820), .B1(new_n826), .B2(new_n819), .ZN(new_n827));
  INV_X1    g641(.A(new_n699), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n769), .A2(new_n395), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n607), .A3(new_n780), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT117), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n829), .A2(new_n832), .A3(new_n607), .A4(new_n780), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n623), .A2(new_n631), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT118), .Z(new_n836));
  NOR3_X1   g650(.A1(new_n751), .A2(new_n395), .A3(new_n718), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n724), .A3(new_n699), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n839), .A2(new_n779), .A3(new_n840), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n769), .A2(new_n828), .A3(new_n751), .A4(new_n395), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n793), .ZN(new_n843));
  OAI22_X1  g657(.A1(new_n838), .A2(new_n674), .B1(KEYINPUT116), .B2(KEYINPUT50), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n491), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n772), .B(new_n773), .C1(new_n846), .C2(new_n777), .ZN(new_n847));
  INV_X1    g661(.A(new_n837), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n769), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n845), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n836), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n738), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n842), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n856), .A2(KEYINPUT48), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n208), .A2(G952), .ZN(new_n860));
  INV_X1    g674(.A(new_n710), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n860), .B1(new_n837), .B2(new_n861), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n859), .B(new_n862), .C1(new_n855), .C2(new_n857), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n831), .A2(new_n833), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n863), .B1(new_n788), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n853), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n851), .A2(new_n852), .ZN(new_n867));
  NOR3_X1   g681(.A1(new_n827), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(G952), .A2(G953), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n783), .B1(new_n868), .B2(new_n869), .ZN(G75));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n817), .A2(new_n816), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n823), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(G902), .ZN(new_n874));
  INV_X1    g688(.A(G210), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n871), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n298), .A2(new_n300), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n290), .B2(new_n298), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n211), .ZN(new_n879));
  XNOR2_X1  g693(.A(KEYINPUT120), .B(KEYINPUT55), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n879), .B(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n876), .A2(new_n881), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n208), .A2(G952), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G51));
  AND4_X1   g699(.A1(G902), .A2(new_n873), .A3(new_n756), .A4(new_n755), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n873), .A2(KEYINPUT54), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n820), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n728), .B(KEYINPUT57), .Z(new_n889));
  AOI21_X1  g703(.A(new_n697), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n889), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n887), .B2(new_n820), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT121), .B1(new_n894), .B2(new_n697), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n884), .B1(new_n892), .B2(new_n895), .ZN(G54));
  NAND4_X1  g710(.A1(new_n873), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n897));
  INV_X1    g711(.A(new_n407), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n884), .ZN(G60));
  INV_X1    g715(.A(new_n884), .ZN(new_n902));
  INV_X1    g716(.A(new_n888), .ZN(new_n903));
  XNOR2_X1  g717(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n359), .A2(new_n314), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n626), .A2(new_n627), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n902), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n827), .A2(new_n906), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n628), .B2(new_n909), .ZN(G63));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n911));
  NAND2_X1  g725(.A1(G217), .A2(G902), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT60), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n818), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n590), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n911), .B1(new_n915), .B2(KEYINPUT124), .ZN(new_n916));
  INV_X1    g730(.A(new_n913), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n873), .A2(new_n649), .A3(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n914), .B2(new_n590), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n916), .A2(new_n902), .A3(new_n918), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n918), .A2(new_n902), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n911), .B1(new_n922), .B2(new_n915), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT123), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT123), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n925), .B(new_n911), .C1(new_n922), .C2(new_n915), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n921), .A2(new_n924), .A3(new_n926), .ZN(G66));
  INV_X1    g741(.A(new_n399), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n208), .B1(new_n928), .B2(G224), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n787), .A2(new_n800), .ZN(new_n930));
  INV_X1    g744(.A(new_n792), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n929), .B1(new_n932), .B2(new_n208), .ZN(new_n933));
  INV_X1    g747(.A(G898), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n878), .B1(new_n934), .B2(G953), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G69));
  INV_X1    g750(.A(new_n774), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n766), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n771), .A2(new_n665), .A3(new_n807), .A4(new_n854), .ZN(new_n939));
  INV_X1    g753(.A(new_n802), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n746), .A3(new_n940), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n938), .A2(new_n744), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n208), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n467), .B(new_n404), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(G900), .B2(G953), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n788), .A2(new_n642), .ZN(new_n946));
  NOR4_X1   g760(.A1(new_n769), .A2(new_n740), .A3(new_n666), .A4(new_n946), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n947), .B(KEYINPUT125), .Z(new_n948));
  NAND2_X1  g762(.A1(new_n686), .A2(new_n940), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n949), .B2(KEYINPUT62), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n949), .A2(KEYINPUT62), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n950), .A2(new_n766), .A3(new_n937), .A4(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n208), .ZN(new_n953));
  AOI22_X1  g767(.A1(new_n943), .A2(new_n945), .B1(new_n953), .B2(new_n944), .ZN(new_n954));
  OAI21_X1  g768(.A(G953), .B1(new_n525), .B2(new_n655), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G72));
  NAND2_X1  g770(.A1(G472), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n952), .B2(new_n932), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT126), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(new_n675), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n960), .B1(new_n959), .B2(new_n675), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n675), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n468), .A2(new_n456), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n964), .A2(new_n965), .A3(new_n958), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n826), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n942), .A2(new_n931), .A3(new_n930), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n965), .B1(new_n968), .B2(new_n958), .ZN(new_n969));
  NOR4_X1   g783(.A1(new_n963), .A2(new_n884), .A3(new_n967), .A4(new_n969), .ZN(G57));
endmodule


