

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U549 ( .A1(n535), .A2(n533), .ZN(n532) );
  OR2_X2 U550 ( .A1(n641), .A2(n640), .ZN(n518) );
  AND2_X2 U551 ( .A1(n639), .A2(G114), .ZN(n640) );
  AND2_X1 U552 ( .A1(n1011), .A2(n521), .ZN(n728) );
  NAND2_X1 U553 ( .A1(n633), .A2(n632), .ZN(n999) );
  AND2_X2 U554 ( .A1(n581), .A2(G2104), .ZN(n911) );
  NOR2_X2 U555 ( .A1(G651), .A2(G543), .ZN(n820) );
  XNOR2_X2 U556 ( .A(n710), .B(KEYINPUT32), .ZN(n719) );
  AND2_X1 U557 ( .A1(n712), .A2(n706), .ZN(n705) );
  INV_X1 U558 ( .A(KEYINPUT65), .ZN(n652) );
  NOR2_X1 U559 ( .A1(n999), .A2(n651), .ZN(n653) );
  NAND2_X1 U560 ( .A1(n672), .A2(n554), .ZN(n678) );
  XNOR2_X1 U561 ( .A(n556), .B(n555), .ZN(n554) );
  INV_X1 U562 ( .A(KEYINPUT27), .ZN(n555) );
  OR2_X1 U563 ( .A1(n707), .A2(G286), .ZN(n708) );
  NAND2_X1 U564 ( .A1(n1006), .A2(n545), .ZN(n544) );
  XOR2_X1 U565 ( .A(KEYINPUT98), .B(n686), .Z(n687) );
  NOR2_X1 U566 ( .A1(n726), .A2(n720), .ZN(n1007) );
  NAND2_X1 U567 ( .A1(G1976), .A2(G288), .ZN(n1006) );
  NAND2_X1 U568 ( .A1(n532), .A2(n530), .ZN(n710) );
  NAND2_X1 U569 ( .A1(n531), .A2(KEYINPUT102), .ZN(n530) );
  NAND2_X1 U570 ( .A1(G160), .A2(G40), .ZN(n741) );
  NAND2_X1 U571 ( .A1(n629), .A2(n548), .ZN(n547) );
  XNOR2_X1 U572 ( .A(n628), .B(n549), .ZN(n548) );
  XNOR2_X1 U573 ( .A(KEYINPUT12), .B(KEYINPUT70), .ZN(n549) );
  INV_X1 U574 ( .A(KEYINPUT13), .ZN(n546) );
  NAND2_X1 U575 ( .A1(n528), .A2(n525), .ZN(n634) );
  AND2_X1 U576 ( .A1(n527), .A2(n526), .ZN(n525) );
  NAND2_X1 U577 ( .A1(G2105), .A2(KEYINPUT17), .ZN(n526) );
  AND2_X1 U578 ( .A1(G2105), .A2(G126), .ZN(n557) );
  INV_X1 U579 ( .A(G2104), .ZN(n588) );
  INV_X1 U580 ( .A(KEYINPUT0), .ZN(n560) );
  XNOR2_X1 U581 ( .A(KEYINPUT68), .B(G543), .ZN(n561) );
  AND2_X1 U582 ( .A1(n588), .A2(G2105), .ZN(n916) );
  XNOR2_X1 U583 ( .A(n582), .B(KEYINPUT23), .ZN(n583) );
  INV_X1 U584 ( .A(KEYINPUT66), .ZN(n582) );
  NAND2_X1 U585 ( .A1(n671), .A2(G2072), .ZN(n556) );
  NAND2_X1 U586 ( .A1(n657), .A2(n656), .ZN(n670) );
  INV_X1 U587 ( .A(n711), .ZN(n691) );
  XOR2_X1 U588 ( .A(KEYINPUT28), .B(n679), .Z(n680) );
  XNOR2_X1 U589 ( .A(n699), .B(n698), .ZN(n712) );
  NOR2_X1 U590 ( .A1(n697), .A2(n696), .ZN(n699) );
  AND2_X1 U591 ( .A1(n708), .A2(n709), .ZN(n536) );
  AND2_X1 U592 ( .A1(n534), .A2(G8), .ZN(n533) );
  OR2_X1 U593 ( .A1(n708), .A2(n709), .ZN(n534) );
  AND2_X1 U594 ( .A1(n538), .A2(n519), .ZN(n542) );
  AND2_X1 U595 ( .A1(n1007), .A2(KEYINPUT103), .ZN(n541) );
  INV_X1 U596 ( .A(KEYINPUT33), .ZN(n724) );
  NOR2_X1 U597 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n529) );
  NAND2_X1 U598 ( .A1(G2104), .A2(KEYINPUT17), .ZN(n527) );
  INV_X1 U599 ( .A(KEYINPUT105), .ZN(n551) );
  NOR2_X1 U600 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U601 ( .A1(n631), .A2(n630), .ZN(n633) );
  XNOR2_X1 U602 ( .A(n547), .B(n546), .ZN(n630) );
  NAND2_X1 U603 ( .A1(G102), .A2(n911), .ZN(n635) );
  XNOR2_X1 U604 ( .A(n638), .B(KEYINPUT85), .ZN(n641) );
  NAND2_X1 U605 ( .A1(n588), .A2(n557), .ZN(n638) );
  NOR2_X2 U606 ( .A1(n593), .A2(n592), .ZN(G160) );
  OR2_X1 U607 ( .A1(n1006), .A2(n545), .ZN(n517) );
  AND2_X1 U608 ( .A1(n543), .A2(n517), .ZN(n519) );
  AND2_X1 U609 ( .A1(n718), .A2(n539), .ZN(n520) );
  XNOR2_X1 U610 ( .A(n667), .B(KEYINPUT15), .ZN(n795) );
  OR2_X1 U611 ( .A1(n727), .A2(n740), .ZN(n521) );
  XOR2_X1 U612 ( .A(n775), .B(KEYINPUT96), .Z(n522) );
  NOR2_X1 U613 ( .A1(n740), .A2(n739), .ZN(n523) );
  AND2_X1 U614 ( .A1(n552), .A2(n790), .ZN(n524) );
  INV_X1 U615 ( .A(KEYINPUT102), .ZN(n709) );
  NAND2_X1 U616 ( .A1(n529), .A2(n581), .ZN(n528) );
  INV_X1 U617 ( .A(n537), .ZN(n531) );
  NAND2_X1 U618 ( .A1(n537), .A2(n536), .ZN(n535) );
  NAND2_X1 U619 ( .A1(n713), .A2(n705), .ZN(n537) );
  NAND2_X1 U620 ( .A1(n719), .A2(n718), .ZN(n731) );
  NAND2_X1 U621 ( .A1(n719), .A2(n520), .ZN(n538) );
  INV_X1 U622 ( .A(n544), .ZN(n539) );
  NAND2_X1 U623 ( .A1(n542), .A2(n540), .ZN(n722) );
  NAND2_X1 U624 ( .A1(n731), .A2(n541), .ZN(n540) );
  OR2_X1 U625 ( .A1(n1007), .A2(n544), .ZN(n543) );
  INV_X1 U626 ( .A(KEYINPUT103), .ZN(n545) );
  NAND2_X1 U627 ( .A1(n550), .A2(n558), .ZN(n553) );
  XNOR2_X1 U628 ( .A(n737), .B(n551), .ZN(n550) );
  NAND2_X1 U629 ( .A1(n553), .A2(n524), .ZN(n791) );
  NAND2_X1 U630 ( .A1(n558), .A2(n523), .ZN(n552) );
  BUF_X1 U631 ( .A(n655), .Z(n742) );
  AND2_X1 U632 ( .A1(n655), .A2(n646), .ZN(n648) );
  AND2_X1 U633 ( .A1(n655), .A2(n654), .ZN(n671) );
  AND2_X1 U634 ( .A1(n522), .A2(n776), .ZN(n558) );
  INV_X1 U635 ( .A(KEYINPUT26), .ZN(n647) );
  BUF_X1 U636 ( .A(n690), .Z(n700) );
  INV_X1 U637 ( .A(KEYINPUT31), .ZN(n698) );
  INV_X1 U638 ( .A(G2105), .ZN(n581) );
  XNOR2_X1 U639 ( .A(n584), .B(n583), .ZN(n587) );
  INV_X1 U640 ( .A(G651), .ZN(n567) );
  NOR2_X1 U641 ( .A1(G543), .A2(n567), .ZN(n559) );
  XOR2_X2 U642 ( .A(KEYINPUT1), .B(n559), .Z(n819) );
  NAND2_X1 U643 ( .A1(G63), .A2(n819), .ZN(n563) );
  XNOR2_X2 U644 ( .A(n561), .B(n560), .ZN(n578) );
  NOR2_X2 U645 ( .A1(G651), .A2(n578), .ZN(n827) );
  NAND2_X1 U646 ( .A1(G51), .A2(n827), .ZN(n562) );
  NAND2_X1 U647 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U648 ( .A(KEYINPUT6), .B(n564), .ZN(n572) );
  NAND2_X1 U649 ( .A1(G89), .A2(n820), .ZN(n565) );
  XNOR2_X1 U650 ( .A(n565), .B(KEYINPUT4), .ZN(n566) );
  XNOR2_X1 U651 ( .A(n566), .B(KEYINPUT74), .ZN(n569) );
  NOR2_X4 U652 ( .A1(n578), .A2(n567), .ZN(n823) );
  NAND2_X1 U653 ( .A1(G76), .A2(n823), .ZN(n568) );
  NAND2_X1 U654 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U655 ( .A(n570), .B(KEYINPUT5), .Z(n571) );
  NOR2_X1 U656 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U657 ( .A(KEYINPUT75), .B(n573), .Z(n574) );
  XOR2_X1 U658 ( .A(KEYINPUT7), .B(n574), .Z(G168) );
  XOR2_X1 U659 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U660 ( .A1(G49), .A2(n827), .ZN(n576) );
  NAND2_X1 U661 ( .A1(G74), .A2(G651), .ZN(n575) );
  NAND2_X1 U662 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U663 ( .A1(n819), .A2(n577), .ZN(n580) );
  NAND2_X1 U664 ( .A1(G87), .A2(n578), .ZN(n579) );
  NAND2_X1 U665 ( .A1(n580), .A2(n579), .ZN(G288) );
  NAND2_X1 U666 ( .A1(G101), .A2(n911), .ZN(n584) );
  INV_X1 U667 ( .A(n634), .ZN(n585) );
  INV_X1 U668 ( .A(n585), .ZN(n743) );
  NAND2_X1 U669 ( .A1(G137), .A2(n743), .ZN(n586) );
  NAND2_X1 U670 ( .A1(n587), .A2(n586), .ZN(n593) );
  NAND2_X1 U671 ( .A1(G125), .A2(n916), .ZN(n591) );
  NAND2_X1 U672 ( .A1(G2104), .A2(G2105), .ZN(n589) );
  XNOR2_X2 U673 ( .A(n589), .B(KEYINPUT67), .ZN(n639) );
  NAND2_X1 U674 ( .A1(G113), .A2(n639), .ZN(n590) );
  NAND2_X1 U675 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U676 ( .A1(G65), .A2(n819), .ZN(n595) );
  NAND2_X1 U677 ( .A1(G91), .A2(n820), .ZN(n594) );
  NAND2_X1 U678 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U679 ( .A1(G78), .A2(n823), .ZN(n597) );
  NAND2_X1 U680 ( .A1(G53), .A2(n827), .ZN(n596) );
  NAND2_X1 U681 ( .A1(n597), .A2(n596), .ZN(n598) );
  OR2_X1 U682 ( .A1(n599), .A2(n598), .ZN(G299) );
  NAND2_X1 U683 ( .A1(G90), .A2(n820), .ZN(n601) );
  NAND2_X1 U684 ( .A1(G77), .A2(n823), .ZN(n600) );
  NAND2_X1 U685 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U686 ( .A(KEYINPUT9), .B(n602), .ZN(n606) );
  NAND2_X1 U687 ( .A1(G64), .A2(n819), .ZN(n604) );
  NAND2_X1 U688 ( .A1(G52), .A2(n827), .ZN(n603) );
  AND2_X1 U689 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U690 ( .A1(n606), .A2(n605), .ZN(G301) );
  INV_X1 U691 ( .A(G301), .ZN(G171) );
  NAND2_X1 U692 ( .A1(G88), .A2(n820), .ZN(n608) );
  NAND2_X1 U693 ( .A1(G75), .A2(n823), .ZN(n607) );
  NAND2_X1 U694 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U695 ( .A1(G62), .A2(n819), .ZN(n610) );
  NAND2_X1 U696 ( .A1(G50), .A2(n827), .ZN(n609) );
  NAND2_X1 U697 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U698 ( .A1(n612), .A2(n611), .ZN(G166) );
  XOR2_X1 U699 ( .A(KEYINPUT88), .B(G166), .Z(G303) );
  NAND2_X1 U700 ( .A1(n827), .A2(G48), .ZN(n619) );
  NAND2_X1 U701 ( .A1(G61), .A2(n819), .ZN(n614) );
  NAND2_X1 U702 ( .A1(G86), .A2(n820), .ZN(n613) );
  NAND2_X1 U703 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U704 ( .A1(n823), .A2(G73), .ZN(n615) );
  XOR2_X1 U705 ( .A(KEYINPUT2), .B(n615), .Z(n616) );
  NOR2_X1 U706 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U707 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U708 ( .A(KEYINPUT81), .B(n620), .Z(G305) );
  AND2_X1 U709 ( .A1(n819), .A2(G60), .ZN(n624) );
  NAND2_X1 U710 ( .A1(G85), .A2(n820), .ZN(n622) );
  NAND2_X1 U711 ( .A1(G72), .A2(n823), .ZN(n621) );
  NAND2_X1 U712 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U713 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U714 ( .A1(n827), .A2(G47), .ZN(n625) );
  NAND2_X1 U715 ( .A1(n626), .A2(n625), .ZN(G290) );
  NAND2_X1 U716 ( .A1(G56), .A2(n819), .ZN(n627) );
  XOR2_X1 U717 ( .A(KEYINPUT14), .B(n627), .Z(n631) );
  NAND2_X1 U718 ( .A1(G81), .A2(n820), .ZN(n628) );
  NAND2_X1 U719 ( .A1(G68), .A2(n823), .ZN(n629) );
  NAND2_X1 U720 ( .A1(n827), .A2(G43), .ZN(n632) );
  NAND2_X1 U721 ( .A1(n634), .A2(G138), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U723 ( .A(n637), .B(KEYINPUT86), .ZN(n642) );
  NOR2_X1 U724 ( .A1(n642), .A2(n518), .ZN(n644) );
  INV_X1 U725 ( .A(KEYINPUT87), .ZN(n643) );
  XNOR2_X1 U726 ( .A(n644), .B(n643), .ZN(G164) );
  NOR2_X2 U727 ( .A1(G164), .A2(G1384), .ZN(n655) );
  INV_X1 U728 ( .A(G1996), .ZN(n645) );
  NOR2_X1 U729 ( .A1(n741), .A2(n645), .ZN(n646) );
  XNOR2_X1 U730 ( .A(n648), .B(n647), .ZN(n650) );
  INV_X1 U731 ( .A(n741), .ZN(n654) );
  NAND2_X2 U732 ( .A1(n742), .A2(n654), .ZN(n690) );
  NAND2_X1 U733 ( .A1(n690), .A2(G1341), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U735 ( .A(n653), .B(n652), .ZN(n669) );
  NAND2_X1 U736 ( .A1(G1348), .A2(n690), .ZN(n657) );
  NAND2_X1 U737 ( .A1(G2067), .A2(n671), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n823), .A2(G79), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n658), .B(KEYINPUT72), .ZN(n660) );
  NAND2_X1 U740 ( .A1(G54), .A2(n827), .ZN(n659) );
  NAND2_X1 U741 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U742 ( .A(n661), .B(KEYINPUT73), .ZN(n663) );
  NAND2_X1 U743 ( .A1(G92), .A2(n820), .ZN(n662) );
  NAND2_X1 U744 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U745 ( .A1(G66), .A2(n819), .ZN(n664) );
  XNOR2_X1 U746 ( .A(KEYINPUT71), .B(n664), .ZN(n665) );
  NAND2_X1 U747 ( .A1(n670), .A2(n795), .ZN(n668) );
  NAND2_X1 U748 ( .A1(n669), .A2(n668), .ZN(n676) );
  NOR2_X1 U749 ( .A1(n795), .A2(n670), .ZN(n674) );
  NAND2_X1 U750 ( .A1(G1956), .A2(n690), .ZN(n672) );
  NOR2_X1 U751 ( .A1(G299), .A2(n678), .ZN(n673) );
  NOR2_X1 U752 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U754 ( .A(n677), .B(KEYINPUT99), .ZN(n681) );
  NAND2_X1 U755 ( .A1(G299), .A2(n678), .ZN(n679) );
  NOR2_X2 U756 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U757 ( .A(n682), .B(KEYINPUT29), .ZN(n688) );
  XOR2_X1 U758 ( .A(G2078), .B(KEYINPUT25), .Z(n982) );
  NOR2_X1 U759 ( .A1(n982), .A2(n690), .ZN(n683) );
  XNOR2_X1 U760 ( .A(n683), .B(KEYINPUT97), .ZN(n685) );
  INV_X1 U761 ( .A(G1961), .ZN(n1023) );
  NAND2_X1 U762 ( .A1(n1023), .A2(n700), .ZN(n684) );
  NAND2_X1 U763 ( .A1(n685), .A2(n684), .ZN(n695) );
  AND2_X1 U764 ( .A1(n695), .A2(G171), .ZN(n686) );
  NAND2_X1 U765 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U766 ( .A(n689), .B(KEYINPUT100), .ZN(n713) );
  NAND2_X1 U767 ( .A1(G8), .A2(n690), .ZN(n740) );
  NOR2_X1 U768 ( .A1(G1966), .A2(n740), .ZN(n715) );
  NOR2_X1 U769 ( .A1(G2084), .A2(n690), .ZN(n711) );
  NAND2_X1 U770 ( .A1(n691), .A2(G8), .ZN(n692) );
  OR2_X1 U771 ( .A1(n715), .A2(n692), .ZN(n693) );
  XNOR2_X1 U772 ( .A(KEYINPUT30), .B(n693), .ZN(n694) );
  NOR2_X1 U773 ( .A1(G168), .A2(n694), .ZN(n697) );
  NOR2_X1 U774 ( .A1(G171), .A2(n695), .ZN(n696) );
  NOR2_X1 U775 ( .A1(G1971), .A2(n740), .ZN(n702) );
  NOR2_X1 U776 ( .A1(G2090), .A2(n700), .ZN(n701) );
  NOR2_X1 U777 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U778 ( .A1(G303), .A2(n703), .ZN(n704) );
  XOR2_X1 U779 ( .A(KEYINPUT101), .B(n704), .Z(n706) );
  INV_X1 U780 ( .A(n706), .ZN(n707) );
  NAND2_X1 U781 ( .A1(G8), .A2(n711), .ZN(n717) );
  AND2_X1 U782 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U783 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U784 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U785 ( .A1(G1976), .A2(G288), .ZN(n726) );
  NOR2_X1 U786 ( .A1(G303), .A2(G1971), .ZN(n720) );
  INV_X1 U787 ( .A(n740), .ZN(n721) );
  NAND2_X1 U788 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U789 ( .A(n723), .B(KEYINPUT64), .ZN(n725) );
  NAND2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n729) );
  XOR2_X1 U791 ( .A(G1981), .B(G305), .Z(n1011) );
  NAND2_X1 U792 ( .A1(n726), .A2(KEYINPUT33), .ZN(n727) );
  NAND2_X1 U793 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U794 ( .A(n730), .B(KEYINPUT104), .ZN(n736) );
  NOR2_X1 U795 ( .A1(G2090), .A2(G303), .ZN(n732) );
  NAND2_X1 U796 ( .A1(G8), .A2(n732), .ZN(n733) );
  NAND2_X1 U797 ( .A1(n731), .A2(n733), .ZN(n734) );
  NAND2_X1 U798 ( .A1(n734), .A2(n740), .ZN(n735) );
  NAND2_X1 U799 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U800 ( .A1(G1981), .A2(G305), .ZN(n738) );
  XOR2_X1 U801 ( .A(n738), .B(KEYINPUT24), .Z(n739) );
  NOR2_X1 U802 ( .A1(n742), .A2(n741), .ZN(n788) );
  NAND2_X1 U803 ( .A1(G104), .A2(n911), .ZN(n746) );
  NAND2_X1 U804 ( .A1(n743), .A2(G140), .ZN(n744) );
  XOR2_X1 U805 ( .A(KEYINPUT89), .B(n744), .Z(n745) );
  NAND2_X1 U806 ( .A1(n746), .A2(n745), .ZN(n749) );
  XOR2_X1 U807 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n747) );
  XNOR2_X1 U808 ( .A(KEYINPUT34), .B(n747), .ZN(n748) );
  XNOR2_X1 U809 ( .A(n749), .B(n748), .ZN(n754) );
  NAND2_X1 U810 ( .A1(G128), .A2(n916), .ZN(n751) );
  NAND2_X1 U811 ( .A1(G116), .A2(n639), .ZN(n750) );
  NAND2_X1 U812 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U813 ( .A(KEYINPUT35), .B(n752), .Z(n753) );
  NOR2_X1 U814 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U815 ( .A(KEYINPUT36), .B(n755), .ZN(n926) );
  XNOR2_X1 U816 ( .A(G2067), .B(KEYINPUT37), .ZN(n777) );
  NOR2_X1 U817 ( .A1(n926), .A2(n777), .ZN(n967) );
  NAND2_X1 U818 ( .A1(n788), .A2(n967), .ZN(n785) );
  XOR2_X1 U819 ( .A(KEYINPUT95), .B(KEYINPUT38), .Z(n757) );
  NAND2_X1 U820 ( .A1(G105), .A2(n911), .ZN(n756) );
  XNOR2_X1 U821 ( .A(n757), .B(n756), .ZN(n764) );
  NAND2_X1 U822 ( .A1(G141), .A2(n743), .ZN(n759) );
  NAND2_X1 U823 ( .A1(G117), .A2(n639), .ZN(n758) );
  NAND2_X1 U824 ( .A1(n759), .A2(n758), .ZN(n762) );
  NAND2_X1 U825 ( .A1(n916), .A2(G129), .ZN(n760) );
  XOR2_X1 U826 ( .A(KEYINPUT94), .B(n760), .Z(n761) );
  NOR2_X1 U827 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U828 ( .A1(n764), .A2(n763), .ZN(n893) );
  NAND2_X1 U829 ( .A1(G1996), .A2(n893), .ZN(n774) );
  NAND2_X1 U830 ( .A1(G107), .A2(n639), .ZN(n765) );
  XNOR2_X1 U831 ( .A(n765), .B(KEYINPUT92), .ZN(n772) );
  NAND2_X1 U832 ( .A1(G95), .A2(n911), .ZN(n767) );
  NAND2_X1 U833 ( .A1(G119), .A2(n916), .ZN(n766) );
  NAND2_X1 U834 ( .A1(n767), .A2(n766), .ZN(n770) );
  NAND2_X1 U835 ( .A1(G131), .A2(n743), .ZN(n768) );
  XNOR2_X1 U836 ( .A(KEYINPUT93), .B(n768), .ZN(n769) );
  NOR2_X1 U837 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U838 ( .A1(n772), .A2(n771), .ZN(n923) );
  NAND2_X1 U839 ( .A1(G1991), .A2(n923), .ZN(n773) );
  NAND2_X1 U840 ( .A1(n774), .A2(n773), .ZN(n959) );
  NAND2_X1 U841 ( .A1(n788), .A2(n959), .ZN(n781) );
  NAND2_X1 U842 ( .A1(n785), .A2(n781), .ZN(n775) );
  XNOR2_X1 U843 ( .A(G1986), .B(G290), .ZN(n1005) );
  NAND2_X1 U844 ( .A1(n1005), .A2(n788), .ZN(n776) );
  NAND2_X1 U845 ( .A1(n926), .A2(n777), .ZN(n970) );
  NOR2_X1 U846 ( .A1(n923), .A2(G1991), .ZN(n778) );
  XNOR2_X1 U847 ( .A(n778), .B(KEYINPUT107), .ZN(n964) );
  NOR2_X1 U848 ( .A1(G1986), .A2(G290), .ZN(n779) );
  XOR2_X1 U849 ( .A(n779), .B(KEYINPUT106), .Z(n780) );
  NAND2_X1 U850 ( .A1(n964), .A2(n780), .ZN(n782) );
  NAND2_X1 U851 ( .A1(n782), .A2(n781), .ZN(n783) );
  OR2_X1 U852 ( .A1(n893), .A2(G1996), .ZN(n955) );
  NAND2_X1 U853 ( .A1(n783), .A2(n955), .ZN(n784) );
  XOR2_X1 U854 ( .A(KEYINPUT39), .B(n784), .Z(n786) );
  NAND2_X1 U855 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U856 ( .A1(n970), .A2(n787), .ZN(n789) );
  NAND2_X1 U857 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U858 ( .A(n791), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U859 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U860 ( .A(G57), .ZN(G237) );
  INV_X1 U861 ( .A(G132), .ZN(G219) );
  INV_X1 U862 ( .A(G82), .ZN(G220) );
  NAND2_X1 U863 ( .A1(G7), .A2(G661), .ZN(n793) );
  XNOR2_X1 U864 ( .A(n793), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U865 ( .A(G223), .B(KEYINPUT69), .ZN(n859) );
  NAND2_X1 U866 ( .A1(n859), .A2(G567), .ZN(n794) );
  XOR2_X1 U867 ( .A(KEYINPUT11), .B(n794), .Z(G234) );
  INV_X1 U868 ( .A(G860), .ZN(n801) );
  OR2_X1 U869 ( .A1(n999), .A2(n801), .ZN(G153) );
  NAND2_X1 U870 ( .A1(G868), .A2(G301), .ZN(n797) );
  INV_X1 U871 ( .A(G868), .ZN(n840) );
  NAND2_X1 U872 ( .A1(n795), .A2(n840), .ZN(n796) );
  NAND2_X1 U873 ( .A1(n797), .A2(n796), .ZN(G284) );
  XNOR2_X1 U874 ( .A(KEYINPUT76), .B(n840), .ZN(n798) );
  NOR2_X1 U875 ( .A1(G286), .A2(n798), .ZN(n800) );
  NOR2_X1 U876 ( .A1(G868), .A2(G299), .ZN(n799) );
  NOR2_X1 U877 ( .A1(n800), .A2(n799), .ZN(G297) );
  NAND2_X1 U878 ( .A1(n801), .A2(G559), .ZN(n802) );
  INV_X1 U879 ( .A(n795), .ZN(n929) );
  NAND2_X1 U880 ( .A1(n802), .A2(n929), .ZN(n803) );
  XNOR2_X1 U881 ( .A(n803), .B(KEYINPUT77), .ZN(n804) );
  XOR2_X1 U882 ( .A(KEYINPUT16), .B(n804), .Z(G148) );
  NOR2_X1 U883 ( .A1(G868), .A2(n999), .ZN(n807) );
  NAND2_X1 U884 ( .A1(G868), .A2(n929), .ZN(n805) );
  NOR2_X1 U885 ( .A1(G559), .A2(n805), .ZN(n806) );
  NOR2_X1 U886 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U887 ( .A(KEYINPUT78), .B(n808), .ZN(G282) );
  NAND2_X1 U888 ( .A1(G123), .A2(n916), .ZN(n809) );
  XNOR2_X1 U889 ( .A(n809), .B(KEYINPUT18), .ZN(n811) );
  NAND2_X1 U890 ( .A1(n911), .A2(G99), .ZN(n810) );
  NAND2_X1 U891 ( .A1(n811), .A2(n810), .ZN(n815) );
  NAND2_X1 U892 ( .A1(G135), .A2(n743), .ZN(n813) );
  NAND2_X1 U893 ( .A1(G111), .A2(n639), .ZN(n812) );
  NAND2_X1 U894 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U895 ( .A1(n815), .A2(n814), .ZN(n963) );
  XNOR2_X1 U896 ( .A(G2096), .B(n963), .ZN(n817) );
  INV_X1 U897 ( .A(G2100), .ZN(n816) );
  NAND2_X1 U898 ( .A1(n817), .A2(n816), .ZN(G156) );
  NAND2_X1 U899 ( .A1(G559), .A2(n929), .ZN(n818) );
  XNOR2_X1 U900 ( .A(n999), .B(n818), .ZN(n837) );
  NOR2_X1 U901 ( .A1(n837), .A2(G860), .ZN(n831) );
  NAND2_X1 U902 ( .A1(G67), .A2(n819), .ZN(n822) );
  NAND2_X1 U903 ( .A1(G93), .A2(n820), .ZN(n821) );
  NAND2_X1 U904 ( .A1(n822), .A2(n821), .ZN(n826) );
  NAND2_X1 U905 ( .A1(G80), .A2(n823), .ZN(n824) );
  XNOR2_X1 U906 ( .A(KEYINPUT79), .B(n824), .ZN(n825) );
  NOR2_X1 U907 ( .A1(n826), .A2(n825), .ZN(n829) );
  NAND2_X1 U908 ( .A1(n827), .A2(G55), .ZN(n828) );
  NAND2_X1 U909 ( .A1(n829), .A2(n828), .ZN(n839) );
  XOR2_X1 U910 ( .A(n839), .B(KEYINPUT80), .Z(n830) );
  XNOR2_X1 U911 ( .A(n831), .B(n830), .ZN(G145) );
  XNOR2_X1 U912 ( .A(KEYINPUT19), .B(G288), .ZN(n836) );
  XNOR2_X1 U913 ( .A(G290), .B(G299), .ZN(n834) );
  XOR2_X1 U914 ( .A(G166), .B(G305), .Z(n832) );
  XNOR2_X1 U915 ( .A(n839), .B(n832), .ZN(n833) );
  XNOR2_X1 U916 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U917 ( .A(n836), .B(n835), .ZN(n932) );
  XOR2_X1 U918 ( .A(n837), .B(n932), .Z(n838) );
  NAND2_X1 U919 ( .A1(n838), .A2(G868), .ZN(n842) );
  NAND2_X1 U920 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U921 ( .A1(n842), .A2(n841), .ZN(G295) );
  NAND2_X1 U922 ( .A1(G2084), .A2(G2078), .ZN(n843) );
  XOR2_X1 U923 ( .A(KEYINPUT20), .B(n843), .Z(n844) );
  NAND2_X1 U924 ( .A1(G2090), .A2(n844), .ZN(n845) );
  XNOR2_X1 U925 ( .A(KEYINPUT21), .B(n845), .ZN(n846) );
  NAND2_X1 U926 ( .A1(n846), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U927 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U928 ( .A1(G220), .A2(G219), .ZN(n847) );
  XNOR2_X1 U929 ( .A(KEYINPUT22), .B(n847), .ZN(n848) );
  NAND2_X1 U930 ( .A1(n848), .A2(G96), .ZN(n849) );
  NOR2_X1 U931 ( .A1(G218), .A2(n849), .ZN(n850) );
  XOR2_X1 U932 ( .A(KEYINPUT82), .B(n850), .Z(n865) );
  NAND2_X1 U933 ( .A1(n865), .A2(G2106), .ZN(n854) );
  NAND2_X1 U934 ( .A1(G69), .A2(G120), .ZN(n851) );
  NOR2_X1 U935 ( .A1(G237), .A2(n851), .ZN(n852) );
  NAND2_X1 U936 ( .A1(G108), .A2(n852), .ZN(n864) );
  NAND2_X1 U937 ( .A1(G567), .A2(n864), .ZN(n853) );
  NAND2_X1 U938 ( .A1(n854), .A2(n853), .ZN(n855) );
  XNOR2_X1 U939 ( .A(KEYINPUT83), .B(n855), .ZN(G319) );
  NAND2_X1 U940 ( .A1(G661), .A2(G483), .ZN(n857) );
  INV_X1 U941 ( .A(G319), .ZN(n856) );
  NOR2_X1 U942 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U943 ( .A(n858), .B(KEYINPUT84), .ZN(n863) );
  NAND2_X1 U944 ( .A1(G36), .A2(n863), .ZN(G176) );
  NAND2_X1 U945 ( .A1(n859), .A2(G2106), .ZN(n860) );
  XNOR2_X1 U946 ( .A(n860), .B(KEYINPUT108), .ZN(G217) );
  AND2_X1 U947 ( .A1(G15), .A2(G2), .ZN(n861) );
  NAND2_X1 U948 ( .A1(G661), .A2(n861), .ZN(G259) );
  NAND2_X1 U949 ( .A1(G3), .A2(G1), .ZN(n862) );
  NAND2_X1 U950 ( .A1(n863), .A2(n862), .ZN(G188) );
  XNOR2_X1 U951 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  INV_X1 U953 ( .A(G120), .ZN(G236) );
  INV_X1 U954 ( .A(G69), .ZN(G235) );
  NOR2_X1 U955 ( .A1(n865), .A2(n864), .ZN(G325) );
  INV_X1 U956 ( .A(G325), .ZN(G261) );
  XOR2_X1 U957 ( .A(G2096), .B(KEYINPUT43), .Z(n867) );
  XNOR2_X1 U958 ( .A(G2072), .B(G2678), .ZN(n866) );
  XNOR2_X1 U959 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U960 ( .A(n868), .B(KEYINPUT110), .Z(n870) );
  XNOR2_X1 U961 ( .A(G2067), .B(G2090), .ZN(n869) );
  XNOR2_X1 U962 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U963 ( .A(KEYINPUT42), .B(G2100), .Z(n872) );
  XNOR2_X1 U964 ( .A(G2084), .B(G2078), .ZN(n871) );
  XNOR2_X1 U965 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U966 ( .A(n874), .B(n873), .ZN(G227) );
  XOR2_X1 U967 ( .A(G1971), .B(G1956), .Z(n876) );
  XNOR2_X1 U968 ( .A(G1986), .B(G1961), .ZN(n875) );
  XNOR2_X1 U969 ( .A(n876), .B(n875), .ZN(n880) );
  XOR2_X1 U970 ( .A(G1966), .B(G1981), .Z(n878) );
  XNOR2_X1 U971 ( .A(G1996), .B(G1991), .ZN(n877) );
  XNOR2_X1 U972 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U973 ( .A(n880), .B(n879), .Z(n882) );
  XNOR2_X1 U974 ( .A(KEYINPUT111), .B(G2474), .ZN(n881) );
  XNOR2_X1 U975 ( .A(n882), .B(n881), .ZN(n884) );
  XOR2_X1 U976 ( .A(G1976), .B(KEYINPUT41), .Z(n883) );
  XNOR2_X1 U977 ( .A(n884), .B(n883), .ZN(G229) );
  NAND2_X1 U978 ( .A1(G124), .A2(n916), .ZN(n885) );
  XNOR2_X1 U979 ( .A(n885), .B(KEYINPUT44), .ZN(n888) );
  NAND2_X1 U980 ( .A1(G136), .A2(n743), .ZN(n886) );
  XNOR2_X1 U981 ( .A(n886), .B(KEYINPUT112), .ZN(n887) );
  NAND2_X1 U982 ( .A1(n888), .A2(n887), .ZN(n892) );
  NAND2_X1 U983 ( .A1(G100), .A2(n911), .ZN(n890) );
  NAND2_X1 U984 ( .A1(G112), .A2(n639), .ZN(n889) );
  NAND2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n891) );
  NOR2_X1 U986 ( .A1(n892), .A2(n891), .ZN(G162) );
  XOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n895) );
  XOR2_X1 U988 ( .A(n893), .B(n963), .Z(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n907) );
  NAND2_X1 U990 ( .A1(n639), .A2(G118), .ZN(n896) );
  XOR2_X1 U991 ( .A(KEYINPUT113), .B(n896), .Z(n898) );
  NAND2_X1 U992 ( .A1(n916), .A2(G130), .ZN(n897) );
  NAND2_X1 U993 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U994 ( .A(KEYINPUT114), .B(n899), .ZN(n905) );
  NAND2_X1 U995 ( .A1(G142), .A2(n743), .ZN(n901) );
  NAND2_X1 U996 ( .A1(G106), .A2(n911), .ZN(n900) );
  NAND2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U998 ( .A(KEYINPUT115), .B(n902), .ZN(n903) );
  XNOR2_X1 U999 ( .A(KEYINPUT45), .B(n903), .ZN(n904) );
  NOR2_X1 U1000 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1001 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1002 ( .A(G164), .B(G160), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1004 ( .A(G162), .B(n910), .ZN(n925) );
  NAND2_X1 U1005 ( .A1(G103), .A2(n911), .ZN(n912) );
  XNOR2_X1 U1006 ( .A(n912), .B(KEYINPUT116), .ZN(n915) );
  NAND2_X1 U1007 ( .A1(G139), .A2(n743), .ZN(n913) );
  XOR2_X1 U1008 ( .A(KEYINPUT117), .B(n913), .Z(n914) );
  NAND2_X1 U1009 ( .A1(n915), .A2(n914), .ZN(n922) );
  NAND2_X1 U1010 ( .A1(n916), .A2(G127), .ZN(n917) );
  XNOR2_X1 U1011 ( .A(n917), .B(KEYINPUT118), .ZN(n919) );
  NAND2_X1 U1012 ( .A1(G115), .A2(n639), .ZN(n918) );
  NAND2_X1 U1013 ( .A1(n919), .A2(n918), .ZN(n920) );
  XOR2_X1 U1014 ( .A(KEYINPUT47), .B(n920), .Z(n921) );
  NOR2_X1 U1015 ( .A1(n922), .A2(n921), .ZN(n951) );
  XNOR2_X1 U1016 ( .A(n923), .B(n951), .ZN(n924) );
  XNOR2_X1 U1017 ( .A(n925), .B(n924), .ZN(n927) );
  XOR2_X1 U1018 ( .A(n927), .B(n926), .Z(n928) );
  NOR2_X1 U1019 ( .A1(G37), .A2(n928), .ZN(G395) );
  XNOR2_X1 U1020 ( .A(n999), .B(KEYINPUT119), .ZN(n931) );
  XNOR2_X1 U1021 ( .A(G171), .B(n929), .ZN(n930) );
  XNOR2_X1 U1022 ( .A(n931), .B(n930), .ZN(n934) );
  XOR2_X1 U1023 ( .A(n932), .B(G286), .Z(n933) );
  XNOR2_X1 U1024 ( .A(n934), .B(n933), .ZN(n935) );
  NOR2_X1 U1025 ( .A1(G37), .A2(n935), .ZN(G397) );
  XOR2_X1 U1026 ( .A(G2451), .B(G2430), .Z(n937) );
  XNOR2_X1 U1027 ( .A(G2438), .B(G2443), .ZN(n936) );
  XNOR2_X1 U1028 ( .A(n937), .B(n936), .ZN(n943) );
  XOR2_X1 U1029 ( .A(G2435), .B(G2454), .Z(n939) );
  XNOR2_X1 U1030 ( .A(G1348), .B(G1341), .ZN(n938) );
  XNOR2_X1 U1031 ( .A(n939), .B(n938), .ZN(n941) );
  XOR2_X1 U1032 ( .A(G2446), .B(G2427), .Z(n940) );
  XNOR2_X1 U1033 ( .A(n941), .B(n940), .ZN(n942) );
  XOR2_X1 U1034 ( .A(n943), .B(n942), .Z(n944) );
  NAND2_X1 U1035 ( .A1(G14), .A2(n944), .ZN(n950) );
  NAND2_X1 U1036 ( .A1(G319), .A2(n950), .ZN(n947) );
  NOR2_X1 U1037 ( .A1(G227), .A2(G229), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(KEYINPUT49), .B(n945), .ZN(n946) );
  NOR2_X1 U1039 ( .A1(n947), .A2(n946), .ZN(n949) );
  NOR2_X1 U1040 ( .A1(G395), .A2(G397), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n949), .A2(n948), .ZN(G225) );
  INV_X1 U1042 ( .A(G225), .ZN(G308) );
  INV_X1 U1043 ( .A(G108), .ZN(G238) );
  INV_X1 U1044 ( .A(n950), .ZN(G401) );
  XOR2_X1 U1045 ( .A(G2072), .B(n951), .Z(n953) );
  XOR2_X1 U1046 ( .A(G164), .B(G2078), .Z(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(KEYINPUT50), .B(n954), .ZN(n961) );
  XNOR2_X1 U1049 ( .A(G162), .B(G2090), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1051 ( .A(KEYINPUT51), .B(n957), .Z(n958) );
  NOR2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n972) );
  XOR2_X1 U1054 ( .A(G2084), .B(G160), .Z(n962) );
  NOR2_X1 U1055 ( .A1(n963), .A2(n962), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1057 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(n968), .B(KEYINPUT120), .ZN(n969) );
  NAND2_X1 U1059 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1060 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1061 ( .A(KEYINPUT52), .B(n973), .ZN(n974) );
  INV_X1 U1062 ( .A(KEYINPUT55), .ZN(n995) );
  NAND2_X1 U1063 ( .A1(n974), .A2(n995), .ZN(n975) );
  NAND2_X1 U1064 ( .A1(n975), .A2(G29), .ZN(n1054) );
  XNOR2_X1 U1065 ( .A(G2090), .B(G35), .ZN(n990) );
  XOR2_X1 U1066 ( .A(G1991), .B(G25), .Z(n976) );
  NAND2_X1 U1067 ( .A1(G28), .A2(n976), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(n977), .B(KEYINPUT121), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(G1996), .B(G32), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(G2072), .B(G33), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n987) );
  XOR2_X1 U1073 ( .A(n982), .B(G27), .Z(n985) );
  XOR2_X1 U1074 ( .A(G26), .B(KEYINPUT122), .Z(n983) );
  XNOR2_X1 U1075 ( .A(G2067), .B(n983), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(KEYINPUT53), .B(n988), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1080 ( .A(G2084), .B(G34), .Z(n991) );
  XNOR2_X1 U1081 ( .A(KEYINPUT54), .B(n991), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(n995), .B(n994), .ZN(n997) );
  INV_X1 U1084 ( .A(G29), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1086 ( .A1(G11), .A2(n998), .ZN(n1052) );
  XNOR2_X1 U1087 ( .A(G16), .B(KEYINPUT56), .ZN(n1022) );
  XNOR2_X1 U1088 ( .A(G171), .B(G1961), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(n999), .B(G1341), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(G299), .B(G1956), .ZN(n1000) );
  NOR2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1020) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  AND2_X1 U1095 ( .A1(G303), .A2(G1971), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(KEYINPUT124), .B(n1010), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G168), .ZN(n1012) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(n1013), .B(KEYINPUT57), .ZN(n1014) );
  NAND2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(n795), .B(G1348), .Z(n1016) );
  XNOR2_X1 U1103 ( .A(KEYINPUT123), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1050) );
  INV_X1 U1107 ( .A(G16), .ZN(n1048) );
  XNOR2_X1 U1108 ( .A(n1023), .B(G5), .ZN(n1044) );
  XOR2_X1 U1109 ( .A(G1966), .B(G21), .Z(n1034) );
  XNOR2_X1 U1110 ( .A(G1348), .B(KEYINPUT59), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(n1024), .B(G4), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(G1981), .B(G6), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(G1341), .B(G19), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(KEYINPUT125), .B(G1956), .Z(n1029) );
  XNOR2_X1 U1117 ( .A(G20), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1119 ( .A(KEYINPUT60), .B(n1032), .ZN(n1033) );
  NAND2_X1 U1120 ( .A1(n1034), .A2(n1033), .ZN(n1042) );
  XNOR2_X1 U1121 ( .A(G1986), .B(G24), .ZN(n1036) );
  XNOR2_X1 U1122 ( .A(G23), .B(G1976), .ZN(n1035) );
  NOR2_X1 U1123 ( .A1(n1036), .A2(n1035), .ZN(n1039) );
  XOR2_X1 U1124 ( .A(G1971), .B(KEYINPUT126), .Z(n1037) );
  XNOR2_X1 U1125 ( .A(G22), .B(n1037), .ZN(n1038) );
  NAND2_X1 U1126 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1127 ( .A(KEYINPUT58), .B(n1040), .ZN(n1041) );
  NOR2_X1 U1128 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NAND2_X1 U1129 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XNOR2_X1 U1130 ( .A(n1045), .B(KEYINPUT127), .ZN(n1046) );
  XNOR2_X1 U1131 ( .A(KEYINPUT61), .B(n1046), .ZN(n1047) );
  NAND2_X1 U1132 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  NAND2_X1 U1133 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  NOR2_X1 U1134 ( .A1(n1052), .A2(n1051), .ZN(n1053) );
  NAND2_X1 U1135 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
  XOR2_X1 U1136 ( .A(KEYINPUT62), .B(n1055), .Z(G311) );
  INV_X1 U1137 ( .A(G311), .ZN(G150) );
endmodule

