//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1039, new_n1040, new_n1041, new_n1042, new_n1044,
    new_n1045;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204));
  AND2_X1   g003(.A1(G113gat), .A2(G120gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(G113gat), .A2(G120gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G134gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G127gat), .ZN(new_n209));
  INV_X1    g008(.A(G127gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G134gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT69), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n204), .B(new_n207), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G113gat), .ZN(new_n215));
  INV_X1    g014(.A(G120gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G113gat), .A2(G120gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n217), .A2(new_n204), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n213), .A3(new_n218), .ZN(new_n220));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n214), .A2(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G141gat), .B(G148gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g027(.A(G155gat), .B(G162gat), .ZN(new_n229));
  OR2_X1    g028(.A1(G141gat), .A2(G148gat), .ZN(new_n230));
  INV_X1    g029(.A(G155gat), .ZN(new_n231));
  INV_X1    g030(.A(G162gat), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT2), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G141gat), .A2(G148gat), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n229), .A2(new_n230), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n228), .B2(new_n235), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT74), .ZN(new_n239));
  OAI211_X1 g038(.A(new_n223), .B(new_n237), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  AOI211_X1 g039(.A(KEYINPUT74), .B(new_n236), .C1(new_n228), .C2(new_n235), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n203), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n237), .A2(new_n214), .A3(new_n222), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n228), .A2(new_n235), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT74), .B1(new_n245), .B2(new_n236), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(new_n239), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n244), .A2(new_n246), .A3(KEYINPUT75), .A4(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n214), .A2(new_n222), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT4), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n245), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n228), .A2(new_n235), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n223), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n254), .B1(new_n214), .B2(new_n222), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n253), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n252), .B1(new_n258), .B2(new_n251), .ZN(new_n259));
  NAND2_X1  g058(.A1(G225gat), .A2(G233gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n249), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT5), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n223), .A2(new_n253), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n245), .A2(new_n250), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n260), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n262), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n250), .A2(KEYINPUT70), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n251), .B(new_n245), .C1(new_n269), .C2(new_n256), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n264), .A2(KEYINPUT4), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n266), .A2(KEYINPUT5), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n249), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT76), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n242), .A2(new_n248), .B1(new_n271), .B2(new_n270), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT76), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n273), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n268), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G1gat), .B(G29gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT0), .ZN(new_n281));
  XNOR2_X1  g080(.A(G57gat), .B(G85gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n279), .A2(KEYINPUT6), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n279), .A2(new_n283), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n286));
  INV_X1    g085(.A(new_n283), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n268), .A2(new_n275), .A3(new_n287), .A4(new_n278), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G197gat), .B(G204gat), .ZN(new_n290));
  INV_X1    g089(.A(G211gat), .ZN(new_n291));
  INV_X1    g090(.A(G218gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n290), .B1(KEYINPUT22), .B2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G211gat), .B(G218gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n294), .B(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G226gat), .ZN(new_n298));
  INV_X1    g097(.A(G233gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G183gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT65), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT65), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G183gat), .ZN(new_n305));
  INV_X1    g104(.A(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT66), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(G190gat), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n303), .A2(new_n305), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(KEYINPUT24), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT24), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n313), .A2(G183gat), .A3(G190gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n317), .A2(G169gat), .A3(G176gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT23), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n318), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n316), .A2(KEYINPUT67), .A3(KEYINPUT25), .A4(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT25), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n322), .ZN(new_n326));
  INV_X1    g125(.A(new_n318), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n312), .A2(new_n314), .B1(new_n302), .B2(new_n306), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n325), .B1(new_n310), .B2(new_n315), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT67), .B1(new_n332), .B2(new_n323), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT66), .B(G190gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT27), .B(G183gat), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n334), .A2(new_n335), .A3(KEYINPUT28), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT27), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(new_n303), .B2(new_n305), .ZN(new_n338));
  NOR2_X1   g137(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n334), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT28), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n336), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR3_X1   g141(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT26), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n321), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n343), .B1(new_n320), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n311), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT68), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT68), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n319), .B1(new_n344), .B2(new_n321), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n349), .B(new_n311), .C1(new_n350), .C2(new_n343), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  OAI22_X1  g151(.A1(new_n331), .A2(new_n333), .B1(new_n342), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n316), .A2(KEYINPUT25), .A3(new_n323), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT67), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(new_n324), .A3(new_n330), .ZN(new_n359));
  INV_X1    g158(.A(new_n339), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT65), .B(G183gat), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n360), .B1(new_n361), .B2(new_n337), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT28), .B1(new_n362), .B2(new_n334), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n348), .B(new_n351), .C1(new_n363), .C2(new_n336), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n359), .A2(KEYINPUT72), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n301), .B1(new_n355), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n300), .A2(KEYINPUT29), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT73), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n359), .A2(KEYINPUT73), .A3(new_n364), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n297), .B1(new_n366), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n367), .A3(new_n365), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n370), .A2(new_n300), .A3(new_n371), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n375), .A3(new_n296), .ZN(new_n376));
  XNOR2_X1  g175(.A(G8gat), .B(G36gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n373), .A2(new_n376), .A3(new_n380), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n381), .A2(KEYINPUT30), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n353), .A2(new_n354), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT72), .B1(new_n359), .B2(new_n364), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n300), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n353), .A2(new_n369), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT73), .B1(new_n359), .B2(new_n364), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n367), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n296), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n374), .A2(new_n375), .A3(new_n296), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n379), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(KEYINPUT30), .A3(new_n381), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n284), .A2(new_n289), .B1(new_n382), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n255), .A2(new_n257), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n353), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n359), .A2(new_n257), .A3(new_n255), .A4(new_n364), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT34), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n398), .B(KEYINPUT64), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(KEYINPUT34), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n400), .A2(KEYINPUT71), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT71), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n399), .A2(new_n404), .A3(KEYINPUT34), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n395), .A2(new_n396), .A3(new_n401), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT33), .ZN(new_n407));
  XOR2_X1   g206(.A(G15gat), .B(G43gat), .Z(new_n408));
  XNOR2_X1  g207(.A(G71gat), .B(G99gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n406), .B(KEYINPUT32), .C1(new_n407), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n406), .A2(new_n407), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n406), .A2(KEYINPUT32), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n414), .A3(new_n410), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n403), .A2(new_n405), .A3(new_n412), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n412), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n395), .A2(new_n396), .B1(G227gat), .B2(G233gat), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT34), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT71), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n397), .A2(new_n402), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n237), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n296), .B1(new_n424), .B2(KEYINPUT29), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT3), .B1(new_n297), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n425), .B1(new_n427), .B2(new_n245), .ZN(new_n428));
  XOR2_X1   g227(.A(G78gat), .B(G106gat), .Z(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT31), .B(G50gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n429), .B(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n428), .B(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G228gat), .A2(G233gat), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n433), .B(G22gat), .Z(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n432), .B(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n416), .A2(new_n423), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n202), .B1(new_n393), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n382), .A2(new_n392), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XOR2_X1   g239(.A(new_n283), .B(KEYINPUT77), .Z(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n279), .A2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n443), .A2(new_n286), .A3(new_n288), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n284), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n202), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT82), .B1(new_n440), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n381), .A2(KEYINPUT30), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n381), .A2(KEYINPUT30), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n448), .B1(new_n449), .B2(new_n391), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n416), .A2(new_n436), .A3(new_n423), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT82), .ZN(new_n453));
  AOI21_X1  g252(.A(KEYINPUT35), .B1(new_n444), .B2(new_n284), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n438), .B1(new_n447), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n416), .A2(KEYINPUT36), .A3(new_n423), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT36), .B1(new_n416), .B2(new_n423), .ZN(new_n459));
  OAI22_X1  g258(.A1(new_n393), .A2(new_n436), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT78), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n461), .A2(KEYINPUT40), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n276), .A2(new_n260), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT39), .B1(new_n265), .B2(new_n266), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n441), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n249), .A2(new_n272), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(new_n266), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n467), .A2(KEYINPUT39), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n462), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n464), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n442), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT39), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n463), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n462), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n471), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n469), .A2(new_n475), .A3(new_n443), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n436), .B1(new_n439), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT37), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n373), .A2(new_n478), .A3(new_n376), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(new_n379), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n478), .B1(new_n373), .B2(new_n376), .ZN(new_n481));
  OAI211_X1 g280(.A(KEYINPUT80), .B(KEYINPUT38), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT37), .B1(new_n389), .B2(new_n390), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(new_n379), .A3(new_n479), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT80), .B1(new_n485), .B2(KEYINPUT38), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n444), .A2(new_n284), .A3(new_n381), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT38), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n479), .A2(new_n489), .A3(new_n379), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n385), .A2(new_n388), .A3(new_n296), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT79), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n385), .A2(new_n388), .A3(KEYINPUT79), .A4(new_n296), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n374), .A2(new_n375), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n297), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n490), .B1(KEYINPUT37), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n488), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n477), .B1(new_n487), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT81), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n460), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n488), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n497), .A2(KEYINPUT37), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n479), .A2(new_n489), .A3(new_n379), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(KEYINPUT38), .B1(new_n480), .B2(new_n481), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT80), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n503), .A2(new_n506), .A3(new_n509), .A4(new_n482), .ZN(new_n510));
  INV_X1    g309(.A(new_n436), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n469), .A2(new_n443), .A3(new_n475), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n450), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT81), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n456), .B1(new_n502), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(G8gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n518), .A2(G1gat), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n517), .B1(new_n519), .B2(KEYINPUT84), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n518), .B1(new_n521), .B2(G1gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n520), .B(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G29gat), .A2(G36gat), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR3_X1   g326(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n530));
  INV_X1    g329(.A(G43gat), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT83), .B1(new_n531), .B2(G50gat), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n529), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n529), .A2(new_n530), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n524), .A2(new_n535), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT85), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT17), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n520), .B(new_n523), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n539), .A2(new_n544), .A3(KEYINPUT18), .A4(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT11), .ZN(new_n548));
  INV_X1    g347(.A(G169gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(G197gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT12), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n543), .A2(new_n540), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT86), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n556), .A2(new_n539), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n545), .B(KEYINPUT13), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n546), .B(new_n554), .C1(new_n557), .C2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n539), .A2(new_n544), .A3(new_n545), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT87), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n561), .A2(KEYINPUT87), .A3(new_n562), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n561), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n556), .A2(new_n539), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n568), .A2(KEYINPUT18), .B1(new_n569), .B2(new_n558), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n554), .B1(new_n570), .B2(new_n563), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n516), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G71gat), .B(G78gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT88), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT9), .ZN(new_n576));
  INV_X1    g375(.A(G71gat), .ZN(new_n577));
  INV_X1    g376(.A(G78gat), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(G57gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n580), .A2(G64gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n580), .A2(G64gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n575), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n581), .B1(new_n583), .B2(KEYINPUT89), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n586), .B1(KEYINPUT89), .B2(new_n581), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(new_n579), .A3(new_n574), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT90), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n585), .A2(KEYINPUT90), .A3(new_n588), .ZN(new_n592));
  AND2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n524), .B1(new_n594), .B2(KEYINPUT21), .ZN(new_n595));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT91), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT91), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n593), .A2(new_n601), .A3(new_n598), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n603), .A2(new_n604), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n597), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n603), .A2(new_n604), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n609), .A2(new_n605), .A3(new_n596), .ZN(new_n610));
  XOR2_X1   g409(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n608), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n608), .B2(new_n610), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n595), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n608), .A2(new_n610), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(new_n611), .ZN(new_n618));
  INV_X1    g417(.A(new_n595), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(new_n619), .A3(new_n613), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G183gat), .B(G211gat), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n616), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G134gat), .B(G162gat), .Z(new_n626));
  NAND2_X1  g425(.A1(G85gat), .A2(G92gat), .ZN(new_n627));
  NAND2_X1  g426(.A1(KEYINPUT92), .A2(KEYINPUT7), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n627), .B(new_n628), .Z(new_n629));
  INV_X1    g428(.A(KEYINPUT8), .ZN(new_n630));
  AND2_X1   g429(.A1(G99gat), .A2(G106gat), .ZN(new_n631));
  OAI221_X1 g430(.A(new_n629), .B1(new_n630), .B2(new_n631), .C1(G85gat), .C2(G92gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G99gat), .B(G106gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT93), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n632), .B(new_n634), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n542), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT41), .ZN(new_n637));
  NAND2_X1  g436(.A1(G232gat), .A2(G233gat), .ZN(new_n638));
  OAI22_X1  g437(.A1(new_n635), .A2(new_n540), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G190gat), .B(G218gat), .ZN(new_n640));
  OR3_X1    g439(.A1(new_n636), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n637), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n640), .B1(new_n636), .B2(new_n639), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n642), .B1(new_n641), .B2(new_n643), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n626), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n646), .ZN(new_n648));
  INV_X1    g447(.A(new_n626), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n644), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT94), .B1(new_n635), .B2(new_n589), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n635), .A2(new_n592), .A3(new_n591), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT10), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n593), .A2(KEYINPUT94), .A3(new_n635), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n593), .A2(new_n658), .A3(new_n635), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n654), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT96), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n657), .A2(new_n659), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n654), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(KEYINPUT95), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT95), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n668), .A2(new_n671), .A3(new_n654), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n667), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n668), .B2(new_n654), .ZN(new_n674));
  AOI211_X1 g473(.A(KEYINPUT95), .B(new_n653), .C1(new_n657), .C2(new_n659), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n674), .A2(new_n675), .A3(KEYINPUT96), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n666), .B1(new_n673), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(KEYINPUT97), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n670), .A2(new_n667), .A3(new_n672), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT96), .B1(new_n674), .B2(new_n675), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT97), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n666), .ZN(new_n683));
  INV_X1    g482(.A(new_n662), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n672), .A3(new_n670), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n678), .A2(new_n683), .B1(new_n665), .B2(new_n685), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n623), .A2(new_n625), .A3(new_n652), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT98), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n616), .A2(new_n620), .A3(new_n624), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n624), .B1(new_n616), .B2(new_n620), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT98), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n691), .A2(new_n692), .A3(new_n652), .A4(new_n686), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n573), .A2(new_n688), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n289), .A2(new_n284), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT100), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT99), .B(G1gat), .Z(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1324gat));
  NOR2_X1   g498(.A1(new_n694), .A2(new_n439), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT16), .B(G8gat), .Z(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(KEYINPUT42), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n704), .B1(new_n703), .B2(new_n705), .ZN(new_n708));
  OAI221_X1 g507(.A(new_n702), .B1(new_n517), .B2(new_n700), .C1(new_n707), .C2(new_n708), .ZN(G1325gat));
  NOR2_X1   g508(.A1(new_n458), .A2(new_n459), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G15gat), .B1(new_n694), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n423), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n417), .A2(new_n422), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n716), .A2(G15gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n712), .B1(new_n694), .B2(new_n717), .ZN(G1326gat));
  NOR2_X1   g517(.A1(new_n694), .A2(new_n436), .ZN(new_n719));
  XOR2_X1   g518(.A(KEYINPUT43), .B(G22gat), .Z(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1327gat));
  NAND2_X1  g520(.A1(new_n685), .A2(new_n665), .ZN(new_n722));
  INV_X1    g521(.A(new_n683), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n682), .B1(new_n681), .B2(new_n666), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n691), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n572), .ZN(new_n727));
  INV_X1    g526(.A(new_n438), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n453), .B1(new_n452), .B2(new_n454), .ZN(new_n729));
  AND4_X1   g528(.A1(new_n453), .A2(new_n454), .A3(new_n437), .A4(new_n439), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n509), .A2(new_n482), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n506), .A2(new_n284), .A3(new_n444), .A4(new_n381), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n501), .B(new_n513), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n393), .ZN(new_n735));
  INV_X1    g534(.A(new_n459), .ZN(new_n736));
  AOI22_X1  g535(.A1(new_n735), .A2(new_n511), .B1(new_n736), .B2(new_n457), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n501), .B1(new_n510), .B2(new_n513), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n731), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n726), .A2(new_n727), .A3(new_n740), .A4(new_n651), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(G29gat), .A3(new_n695), .ZN(new_n742));
  XNOR2_X1  g541(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n740), .A2(KEYINPUT44), .A3(new_n651), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT44), .B1(new_n740), .B2(new_n651), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT103), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n567), .B2(new_n571), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n565), .A2(new_n566), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(new_n570), .A3(new_n554), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n546), .B1(new_n557), .B2(new_n559), .ZN(new_n752));
  INV_X1    g551(.A(new_n563), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n553), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(KEYINPUT103), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n749), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n691), .A2(new_n725), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n747), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G29gat), .B1(new_n758), .B2(new_n695), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n759), .ZN(G1328gat));
  NOR3_X1   g559(.A1(new_n741), .A2(G36gat), .A3(new_n439), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT46), .ZN(new_n762));
  OAI21_X1  g561(.A(G36gat), .B1(new_n758), .B2(new_n439), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(G1329gat));
  OAI21_X1  g563(.A(G43gat), .B1(new_n758), .B2(new_n711), .ZN(new_n765));
  OR3_X1    g564(.A1(new_n741), .A2(G43gat), .A3(new_n716), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT104), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n758), .B2(new_n711), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n747), .A2(KEYINPUT104), .A3(new_n710), .A4(new_n757), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n531), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n766), .A2(KEYINPUT47), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n767), .A2(KEYINPUT47), .B1(new_n771), .B2(new_n772), .ZN(G1330gat));
  INV_X1    g572(.A(G50gat), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT107), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n747), .A2(new_n775), .A3(new_n511), .A4(new_n757), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n777), .B1(new_n516), .B2(new_n652), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n740), .A2(KEYINPUT44), .A3(new_n651), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n778), .A2(new_n511), .A3(new_n779), .A4(new_n757), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT107), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n774), .B1(new_n776), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n741), .A2(KEYINPUT106), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT106), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n573), .A2(new_n784), .A3(new_n651), .A4(new_n726), .ZN(new_n785));
  AOI211_X1 g584(.A(G50gat), .B(new_n436), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT48), .B1(new_n782), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n783), .A2(new_n785), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n436), .A2(G50gat), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT48), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n780), .A2(G50gat), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT105), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT105), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n780), .A2(new_n794), .A3(G50gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n791), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n787), .A2(new_n788), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n788), .B1(new_n787), .B2(new_n796), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(G1331gat));
  NAND2_X1  g598(.A1(new_n623), .A2(new_n625), .ZN(new_n800));
  INV_X1    g599(.A(new_n756), .ZN(new_n801));
  NOR4_X1   g600(.A1(new_n800), .A2(new_n651), .A3(new_n686), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(new_n740), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n695), .B(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(new_n580), .ZN(G1332gat));
  INV_X1    g607(.A(new_n803), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n450), .ZN(new_n810));
  NOR2_X1   g609(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n811));
  AND2_X1   g610(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n811), .B2(new_n810), .ZN(G1333gat));
  XNOR2_X1  g613(.A(new_n715), .B(KEYINPUT110), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n803), .A2(G71gat), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n809), .A2(new_n710), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(G71gat), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g618(.A1(new_n809), .A2(new_n511), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT112), .ZN(new_n821));
  XNOR2_X1  g620(.A(KEYINPUT111), .B(G78gat), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n821), .B(new_n822), .ZN(G1335gat));
  OAI211_X1 g622(.A(new_n725), .B(new_n756), .C1(new_n689), .C2(new_n690), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n747), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G85gat), .B1(new_n826), .B2(new_n695), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n740), .A2(new_n651), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n800), .A2(new_n756), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n691), .A2(new_n801), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n832), .A2(KEYINPUT51), .A3(new_n740), .A4(new_n651), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(KEYINPUT113), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(KEYINPUT113), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n725), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n695), .A2(G85gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n827), .B1(new_n837), .B2(new_n838), .ZN(G1336gat));
  NAND3_X1  g638(.A1(new_n747), .A2(new_n450), .A3(new_n825), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G92gat), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n686), .A2(G92gat), .A3(new_n439), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT52), .B1(new_n834), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n842), .B(KEYINPUT114), .Z(new_n845));
  AOI22_X1  g644(.A1(new_n840), .A2(G92gat), .B1(new_n834), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT52), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(G1337gat));
  OAI21_X1  g647(.A(G99gat), .B1(new_n826), .B2(new_n711), .ZN(new_n849));
  OR2_X1    g648(.A1(new_n716), .A2(G99gat), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n849), .B1(new_n837), .B2(new_n850), .ZN(G1338gat));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n778), .A2(new_n511), .A3(new_n779), .A4(new_n825), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(G106gat), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n686), .A2(G106gat), .A3(new_n436), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n834), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n855), .B1(new_n834), .B2(new_n856), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n852), .B(new_n854), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n853), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n861), .A2(new_n862), .B1(new_n834), .B2(new_n856), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n859), .B1(new_n863), .B2(new_n852), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n859), .B(KEYINPUT117), .C1(new_n863), .C2(new_n852), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1339gat));
  NAND2_X1  g667(.A1(new_n557), .A2(new_n559), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n539), .A2(new_n544), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(G229gat), .A3(G233gat), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n552), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n567), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n725), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n678), .A2(new_n683), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n660), .A2(new_n654), .A3(new_n661), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n684), .A2(KEYINPUT54), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n665), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n662), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n877), .A2(KEYINPUT55), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT55), .B1(new_n877), .B2(new_n880), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n875), .A2(new_n749), .A3(new_n883), .A4(new_n755), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n651), .B1(new_n874), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n886));
  INV_X1    g685(.A(new_n872), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n751), .B2(new_n887), .ZN(new_n888));
  NOR3_X1   g687(.A1(new_n567), .A2(KEYINPUT118), .A3(new_n872), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n883), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n890), .A2(new_n891), .A3(new_n652), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n800), .B1(new_n885), .B2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n691), .A2(new_n652), .A3(new_n686), .A4(new_n756), .ZN(new_n894));
  AOI211_X1 g693(.A(new_n716), .B(new_n511), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n695), .A2(new_n450), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(new_n215), .A3(new_n572), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n895), .A2(new_n805), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n899), .A2(new_n450), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n801), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n898), .B1(new_n901), .B2(new_n215), .ZN(G1340gat));
  OAI21_X1  g701(.A(G120gat), .B1(new_n897), .B2(new_n686), .ZN(new_n903));
  INV_X1    g702(.A(new_n900), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n686), .A2(G120gat), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT119), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(G1341gat));
  NAND3_X1  g706(.A1(new_n900), .A2(new_n210), .A3(new_n691), .ZN(new_n908));
  OAI21_X1  g707(.A(G127gat), .B1(new_n897), .B2(new_n800), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n908), .A2(KEYINPUT120), .A3(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1342gat));
  NOR4_X1   g713(.A1(new_n899), .A2(G134gat), .A3(new_n450), .A4(new_n652), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT56), .ZN(new_n916));
  OAI21_X1  g715(.A(G134gat), .B1(new_n897), .B2(new_n652), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1343gat));
  AOI21_X1  g717(.A(new_n436), .B1(new_n893), .B2(new_n894), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n806), .A2(new_n710), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n572), .A2(G141gat), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n919), .A2(KEYINPUT122), .A3(new_n920), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n923), .A2(new_n439), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT58), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n711), .A2(new_n896), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n893), .A2(new_n894), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT57), .B1(new_n931), .B2(new_n511), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n436), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n727), .A2(new_n875), .A3(new_n883), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n651), .B1(new_n874), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n800), .B1(new_n937), .B2(new_n892), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n935), .B1(new_n938), .B2(new_n894), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n727), .B(new_n930), .C1(new_n932), .C2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT123), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n938), .A2(new_n894), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(new_n934), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n944), .B1(KEYINPUT57), .B2(new_n919), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n945), .A2(KEYINPUT123), .A3(new_n727), .A4(new_n930), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n946), .A3(G141gat), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n928), .A2(new_n947), .ZN(new_n948));
  NOR4_X1   g747(.A1(new_n921), .A2(G141gat), .A3(new_n572), .A4(new_n450), .ZN(new_n949));
  INV_X1    g748(.A(new_n873), .ZN(new_n950));
  OAI22_X1  g749(.A1(new_n891), .A2(new_n756), .B1(new_n686), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n652), .ZN(new_n952));
  INV_X1    g751(.A(new_n890), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n953), .A2(new_n651), .A3(new_n875), .A4(new_n883), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n691), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n687), .A2(new_n801), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n511), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n939), .B1(new_n957), .B2(new_n933), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT121), .B1(new_n958), .B2(new_n929), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT121), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n960), .A3(new_n930), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n801), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n949), .B1(new_n962), .B2(G141gat), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n948), .B1(new_n963), .B2(new_n927), .ZN(G1344gat));
  NAND3_X1  g763(.A1(new_n959), .A2(new_n725), .A3(new_n961), .ZN(new_n965));
  INV_X1    g764(.A(G148gat), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n966), .A2(KEYINPUT59), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n693), .A2(new_n688), .A3(new_n572), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(new_n938), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n970), .A2(new_n933), .A3(new_n511), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n957), .A2(KEYINPUT57), .ZN(new_n972));
  NAND4_X1  g771(.A1(new_n971), .A2(new_n972), .A3(new_n725), .A4(new_n930), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(G148gat), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(KEYINPUT59), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n968), .A2(new_n975), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n923), .A2(new_n439), .A3(new_n925), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n977), .A2(new_n966), .A3(new_n725), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1345gat));
  NAND2_X1  g778(.A1(new_n959), .A2(new_n961), .ZN(new_n980));
  OAI21_X1  g779(.A(G155gat), .B1(new_n980), .B2(new_n800), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n977), .A2(new_n231), .A3(new_n691), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1346gat));
  OAI21_X1  g782(.A(G162gat), .B1(new_n980), .B2(new_n652), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n652), .A2(G162gat), .A3(new_n450), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n923), .A2(new_n925), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT124), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n986), .A2(KEYINPUT124), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(G1347gat));
  AND2_X1   g788(.A1(new_n931), .A2(new_n695), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n990), .A2(new_n450), .A3(new_n437), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n756), .A2(G169gat), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(KEYINPUT125), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n806), .A2(new_n450), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n995), .A2(new_n815), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n931), .A2(new_n436), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n997), .A2(KEYINPUT126), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT126), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n931), .A2(new_n999), .A3(new_n436), .A4(new_n996), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n998), .A2(new_n727), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1001), .A2(G169gat), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n994), .A2(new_n1002), .ZN(G1348gat));
  INV_X1    g802(.A(G176gat), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n991), .A2(new_n1004), .A3(new_n725), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n998), .A2(new_n725), .A3(new_n1000), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1005), .B1(new_n1004), .B2(new_n1006), .ZN(G1349gat));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n335), .A3(new_n691), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n998), .A2(new_n691), .A3(new_n1000), .ZN(new_n1009));
  INV_X1    g808(.A(new_n361), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(KEYINPUT60), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT60), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1008), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1013), .A2(new_n1015), .ZN(G1350gat));
  NAND3_X1  g815(.A1(new_n991), .A2(new_n334), .A3(new_n651), .ZN(new_n1017));
  NAND3_X1  g816(.A1(new_n998), .A2(new_n651), .A3(new_n1000), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT61), .ZN(new_n1019));
  AND3_X1   g818(.A1(new_n1018), .A2(new_n1019), .A3(G190gat), .ZN(new_n1020));
  AOI21_X1  g819(.A(new_n1019), .B1(new_n1018), .B2(G190gat), .ZN(new_n1021));
  OAI21_X1  g820(.A(new_n1017), .B1(new_n1020), .B2(new_n1021), .ZN(G1351gat));
  AND2_X1   g821(.A1(new_n971), .A2(new_n972), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n995), .A2(new_n710), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NOR3_X1   g824(.A1(new_n1025), .A2(new_n551), .A3(new_n572), .ZN(new_n1026));
  NOR3_X1   g825(.A1(new_n710), .A2(new_n439), .A3(new_n436), .ZN(new_n1027));
  AND2_X1   g826(.A1(new_n990), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g827(.A(G197gat), .B1(new_n1028), .B2(new_n801), .ZN(new_n1029));
  NOR2_X1   g828(.A1(new_n1026), .A2(new_n1029), .ZN(G1352gat));
  NOR2_X1   g829(.A1(new_n686), .A2(G204gat), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n990), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1032), .A2(KEYINPUT62), .ZN(new_n1033));
  XOR2_X1   g832(.A(new_n1033), .B(KEYINPUT127), .Z(new_n1034));
  NOR2_X1   g833(.A1(new_n1032), .A2(KEYINPUT62), .ZN(new_n1035));
  NAND3_X1  g834(.A1(new_n1023), .A2(new_n725), .A3(new_n1024), .ZN(new_n1036));
  AOI21_X1  g835(.A(new_n1035), .B1(new_n1036), .B2(G204gat), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1034), .A2(new_n1037), .ZN(G1353gat));
  NAND3_X1  g837(.A1(new_n1028), .A2(new_n291), .A3(new_n691), .ZN(new_n1039));
  NAND4_X1  g838(.A1(new_n971), .A2(new_n972), .A3(new_n691), .A4(new_n1024), .ZN(new_n1040));
  AND3_X1   g839(.A1(new_n1040), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1041));
  AOI21_X1  g840(.A(KEYINPUT63), .B1(new_n1040), .B2(G211gat), .ZN(new_n1042));
  OAI21_X1  g841(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(G1354gat));
  OAI21_X1  g842(.A(G218gat), .B1(new_n1025), .B2(new_n652), .ZN(new_n1044));
  NAND3_X1  g843(.A1(new_n1028), .A2(new_n292), .A3(new_n651), .ZN(new_n1045));
  NAND2_X1  g844(.A1(new_n1044), .A2(new_n1045), .ZN(G1355gat));
endmodule


