//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n593, new_n594, new_n596,
    new_n597, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n630,
    new_n631, new_n632, new_n633, new_n636, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND3_X1  g035(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT66), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G137), .A3(new_n460), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n468), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n460), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR3_X1   g048(.A1(new_n463), .A2(new_n466), .A3(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n468), .A2(new_n470), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT67), .ZN(new_n476));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n464), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n476), .A2(new_n478), .A3(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n476), .A2(new_n478), .A3(new_n460), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n481), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  AND2_X1   g063(.A1(new_n464), .A2(G126), .ZN(new_n489));
  AND2_X1   g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  OAI21_X1  g065(.A(G2105), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n467), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G102), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(KEYINPUT68), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n495), .A2(new_n468), .A3(new_n470), .A4(new_n460), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n464), .A2(KEYINPUT4), .A3(new_n460), .A4(new_n495), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n491), .A2(new_n493), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT69), .A3(KEYINPUT5), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n504), .A2(new_n506), .B1(new_n503), .B2(G543), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(G88), .A3(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n512), .A2(new_n505), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT70), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT70), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n509), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n504), .A2(new_n506), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n503), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(KEYINPUT71), .A3(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n516), .A2(new_n518), .B1(new_n522), .B2(new_n529), .ZN(G166));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT73), .B(G51), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT72), .B1(new_n512), .B2(new_n505), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n534), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n532), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n531), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n534), .B1(new_n508), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(new_n535), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g117(.A(KEYINPUT74), .B(new_n539), .C1(new_n542), .C2(new_n532), .ZN(new_n543));
  NAND4_X1  g118(.A1(new_n524), .A2(G89), .A3(new_n525), .A4(new_n508), .ZN(new_n544));
  NAND3_X1  g119(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT75), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT75), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n547), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(KEYINPUT7), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n548), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT7), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n544), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT76), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n555));
  NAND4_X1  g130(.A1(new_n544), .A2(new_n552), .A3(new_n555), .A4(new_n549), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n538), .A2(new_n543), .B1(new_n554), .B2(new_n556), .ZN(G168));
  AOI22_X1  g132(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n558));
  OR2_X1    g133(.A1(new_n558), .A2(new_n521), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n507), .A2(new_n508), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(KEYINPUT78), .B(G90), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n533), .A2(new_n535), .ZN(new_n564));
  XOR2_X1   g139(.A(KEYINPUT77), .B(G52), .Z(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n559), .A2(new_n563), .A3(new_n566), .ZN(G301));
  INV_X1    g142(.A(G301), .ZN(G171));
  INV_X1    g143(.A(G43), .ZN(new_n569));
  INV_X1    g144(.A(G81), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n542), .A2(new_n569), .B1(new_n570), .B2(new_n560), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n521), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G860), .ZN(G153));
  AND3_X1   g150(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G36), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(G188));
  NAND3_X1  g155(.A1(new_n507), .A2(G91), .A3(new_n508), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n507), .A2(KEYINPUT79), .A3(G91), .A4(new_n508), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G78), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G65), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n526), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n508), .A2(G53), .A3(G543), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT9), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n585), .A2(new_n589), .A3(new_n591), .ZN(G299));
  NAND2_X1  g167(.A1(new_n538), .A2(new_n543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n554), .A2(new_n556), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G286));
  NAND2_X1  g170(.A1(new_n516), .A2(new_n518), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n522), .A2(new_n529), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G303));
  OAI21_X1  g173(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n513), .A2(G49), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n507), .A2(G87), .A3(new_n508), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G288));
  NAND2_X1  g178(.A1(new_n507), .A2(G86), .ZN(new_n604));
  NAND2_X1  g179(.A1(G48), .A2(G543), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(new_n508), .ZN(new_n607));
  NAND2_X1  g182(.A1(G73), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G61), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n526), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G651), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n607), .A2(new_n611), .ZN(G305));
  AOI22_X1  g187(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(new_n521), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n564), .A2(G47), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n561), .A2(G85), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(G290));
  NAND2_X1  g192(.A1(G301), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G92), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n560), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT10), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n564), .A2(G54), .ZN(new_n622));
  NAND2_X1  g197(.A1(G79), .A2(G543), .ZN(new_n623));
  INV_X1    g198(.A(G66), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n526), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G651), .ZN(new_n626));
  AND3_X1   g201(.A1(new_n621), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n618), .B1(new_n627), .B2(G868), .ZN(G284));
  OAI21_X1  g203(.A(new_n618), .B1(new_n627), .B2(G868), .ZN(G321));
  INV_X1    g204(.A(G868), .ZN(new_n630));
  NOR2_X1   g205(.A1(G168), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT80), .ZN(new_n632));
  INV_X1    g207(.A(G299), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(G868), .B2(new_n633), .ZN(G297));
  OAI21_X1  g209(.A(new_n632), .B1(G868), .B2(new_n633), .ZN(G280));
  XNOR2_X1  g210(.A(KEYINPUT81), .B(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n627), .B1(G860), .B2(new_n636), .ZN(G148));
  NAND2_X1  g212(.A1(new_n627), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n574), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n464), .A2(new_n492), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(KEYINPUT12), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2100), .Z(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT82), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  OAI211_X1 g224(.A(new_n648), .B(new_n649), .C1(G111), .C2(new_n460), .ZN(new_n650));
  INV_X1    g225(.A(G123), .ZN(new_n651));
  INV_X1    g226(.A(G135), .ZN(new_n652));
  OAI221_X1 g227(.A(new_n650), .B1(new_n479), .B2(new_n651), .C1(new_n652), .C2(new_n482), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(G2096), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n645), .A2(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT83), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT16), .ZN(new_n658));
  XOR2_X1   g233(.A(G2443), .B(G2446), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1341), .B(G1348), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2427), .B(G2438), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2430), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT15), .B(G2435), .Z(new_n665));
  XOR2_X1   g240(.A(new_n664), .B(new_n665), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT14), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n662), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G14), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G401));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2067), .B(G2678), .Z(new_n673));
  OR2_X1    g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(new_n675), .A3(KEYINPUT17), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT18), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n674), .A2(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2072), .B(G2078), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(new_n680), .B2(new_n678), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2096), .B(G2100), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n686), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  AOI22_X1  g267(.A1(new_n690), .A2(KEYINPUT20), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n694), .A2(new_n686), .A3(new_n689), .ZN(new_n695));
  OAI211_X1 g270(.A(new_n693), .B(new_n695), .C1(KEYINPUT20), .C2(new_n690), .ZN(new_n696));
  XOR2_X1   g271(.A(G1991), .B(G1996), .Z(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n696), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT84), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1981), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  OR2_X1    g279(.A1(G95), .A2(G2105), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n705), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n706));
  INV_X1    g281(.A(G119), .ZN(new_n707));
  INV_X1    g282(.A(G131), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n706), .B1(new_n479), .B2(new_n707), .C1(new_n708), .C2(new_n482), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n480), .A2(G119), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n483), .A2(G131), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n712), .A2(new_n713), .A3(KEYINPUT85), .A4(new_n706), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G29), .ZN(new_n716));
  OR2_X1    g291(.A1(G25), .A2(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(KEYINPUT86), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT86), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n716), .A2(new_n720), .A3(new_n717), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT35), .B(G1991), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n719), .A2(new_n723), .A3(new_n721), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  MUX2_X1   g302(.A(G6), .B(G305), .S(G16), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT89), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT32), .B(G1981), .Z(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT89), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n728), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n730), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G16), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G23), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n602), .B2(new_n737), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT90), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT33), .B(G1976), .Z(new_n741));
  AND2_X1   g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n737), .A2(G22), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G166), .B2(new_n737), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n745), .A2(G1971), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n742), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT34), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n745), .A2(G1971), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n736), .A2(new_n747), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G16), .A2(G24), .ZN(new_n751));
  XOR2_X1   g326(.A(G290), .B(KEYINPUT87), .Z(new_n752));
  AOI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT88), .B(G1986), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n727), .A2(new_n750), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(KEYINPUT91), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n736), .A2(new_n747), .A3(new_n749), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(KEYINPUT34), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n727), .A2(new_n750), .A3(new_n760), .A4(new_n755), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n757), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n763));
  OR2_X1    g338(.A1(KEYINPUT92), .A2(KEYINPUT36), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n763), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n757), .A2(new_n759), .A3(new_n761), .A4(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(KEYINPUT99), .B1(G5), .B2(G16), .ZN(new_n768));
  OR3_X1    g343(.A1(KEYINPUT99), .A2(G5), .A3(G16), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n768), .B(new_n769), .C1(G301), .C2(new_n737), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1961), .ZN(new_n771));
  AND2_X1   g346(.A1(KEYINPUT24), .A2(G34), .ZN(new_n772));
  NOR2_X1   g347(.A1(KEYINPUT24), .A2(G34), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n772), .A2(new_n773), .A3(G29), .ZN(new_n774));
  INV_X1    g349(.A(new_n473), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n775), .A2(new_n462), .A3(new_n465), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n774), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2084), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G29), .ZN(new_n780));
  AND2_X1   g355(.A1(KEYINPUT30), .A2(G28), .ZN(new_n781));
  NOR2_X1   g356(.A1(KEYINPUT30), .A2(G28), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n653), .B2(new_n780), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(G29), .A2(G32), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n483), .A2(G141), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n480), .A2(G129), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT26), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n492), .A2(G105), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n787), .A2(new_n788), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n786), .B1(new_n792), .B2(new_n780), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT27), .B(G1996), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n771), .B(new_n785), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n780), .A2(G35), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G162), .B2(new_n780), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT29), .B(G2090), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n780), .A2(G33), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n492), .A2(G103), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT25), .Z(new_n802));
  AOI22_X1  g377(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n803));
  AOI21_X1  g378(.A(KEYINPUT94), .B1(new_n483), .B2(G139), .ZN(new_n804));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n805));
  INV_X1    g380(.A(G139), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n482), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n802), .B1(new_n460), .B2(new_n803), .C1(new_n804), .C2(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n800), .B1(new_n808), .B2(G29), .ZN(new_n809));
  INV_X1    g384(.A(G2072), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n799), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n780), .A2(G27), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G164), .B2(new_n780), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(G2078), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n737), .A2(G19), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n574), .B2(new_n737), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(G1341), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(G1341), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n815), .A2(G2078), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n795), .A2(new_n813), .A3(new_n816), .A4(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G1966), .ZN(new_n824));
  NAND2_X1  g399(.A1(G168), .A2(G16), .ZN(new_n825));
  OR2_X1    g400(.A1(new_n825), .A2(KEYINPUT96), .ZN(new_n826));
  OAI211_X1 g401(.A(new_n825), .B(KEYINPUT96), .C1(G16), .C2(G21), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT97), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n828), .B1(new_n826), .B2(new_n827), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n824), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n780), .A2(G26), .ZN(new_n832));
  OR2_X1    g407(.A1(G104), .A2(G2105), .ZN(new_n833));
  OAI211_X1 g408(.A(new_n833), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT93), .ZN(new_n835));
  INV_X1    g410(.A(G128), .ZN(new_n836));
  INV_X1    g411(.A(G140), .ZN(new_n837));
  OAI221_X1 g412(.A(new_n835), .B1(new_n479), .B2(new_n836), .C1(new_n837), .C2(new_n482), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n832), .B1(new_n838), .B2(G29), .ZN(new_n839));
  MUX2_X1   g414(.A(new_n832), .B(new_n839), .S(KEYINPUT28), .Z(new_n840));
  INV_X1    g415(.A(G2067), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n737), .A2(G4), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n627), .B2(new_n737), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G1348), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n793), .A2(new_n794), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT95), .Z(new_n847));
  NOR3_X1   g422(.A1(new_n842), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT100), .B(KEYINPUT23), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n737), .A2(G20), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n633), .B2(new_n737), .ZN(new_n852));
  INV_X1    g427(.A(G1956), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n823), .A2(new_n831), .A3(new_n848), .A4(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT31), .B(G11), .Z(new_n856));
  NOR3_X1   g431(.A1(new_n829), .A2(new_n830), .A3(new_n824), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT98), .ZN(new_n858));
  NOR3_X1   g433(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n765), .A2(new_n767), .A3(new_n859), .ZN(G311));
  NAND3_X1  g435(.A1(new_n765), .A2(new_n859), .A3(new_n767), .ZN(G150));
  AOI22_X1  g436(.A1(new_n561), .A2(G93), .B1(new_n564), .B2(G55), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(new_n521), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n865), .A2(G860), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT37), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n627), .A2(G559), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT38), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n574), .A2(new_n865), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n574), .A2(new_n865), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT39), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n869), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n867), .B1(new_n875), .B2(G860), .ZN(G145));
  XNOR2_X1  g451(.A(new_n838), .B(G164), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n792), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n808), .B(KEYINPUT101), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n808), .A2(KEYINPUT101), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n880), .B1(new_n882), .B2(new_n878), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n480), .A2(G130), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n483), .A2(G142), .ZN(new_n886));
  OR2_X1    g461(.A1(G106), .A2(G2105), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n887), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n711), .A2(new_n714), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n711), .B2(new_n714), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT102), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n892), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n895), .A3(new_n890), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n893), .A2(new_n896), .A3(new_n643), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n643), .B1(new_n893), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g473(.A(G160), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n893), .A2(new_n896), .ZN(new_n900));
  INV_X1    g475(.A(new_n643), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n893), .A2(new_n896), .A3(new_n643), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(new_n776), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n487), .B(new_n653), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n899), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(new_n899), .B2(new_n904), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n884), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n905), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n897), .A2(new_n898), .A3(G160), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n776), .B1(new_n902), .B2(new_n903), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n899), .A2(new_n904), .A3(new_n905), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n912), .A2(new_n883), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G37), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n908), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g492(.A1(new_n865), .A2(new_n630), .ZN(new_n918));
  AND2_X1   g493(.A1(G290), .A2(new_n602), .ZN(new_n919));
  NOR2_X1   g494(.A1(G290), .A2(new_n602), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n921));
  OR3_X1    g496(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n919), .B2(new_n920), .ZN(new_n923));
  XNOR2_X1  g498(.A(G166), .B(G305), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n924), .A2(new_n923), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT42), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n873), .B(new_n638), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n621), .A2(new_n622), .A3(new_n626), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n930), .A2(G299), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n620), .A2(KEYINPUT10), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n620), .A2(KEYINPUT10), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n932), .A2(new_n933), .B1(G651), .B2(new_n625), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n633), .B1(new_n934), .B2(new_n622), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n929), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n627), .A2(new_n633), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n930), .A2(G299), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(KEYINPUT41), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT41), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n942), .B1(new_n931), .B2(new_n935), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n938), .B1(new_n929), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n928), .B(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n918), .B1(new_n946), .B2(new_n630), .ZN(G295));
  OAI21_X1  g522(.A(new_n918), .B1(new_n946), .B2(new_n630), .ZN(G331));
  NOR3_X1   g523(.A1(new_n871), .A2(new_n872), .A3(G171), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n574), .A2(new_n865), .ZN(new_n950));
  AOI21_X1  g525(.A(G301), .B1(new_n950), .B2(new_n870), .ZN(new_n951));
  OAI21_X1  g526(.A(G286), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(G171), .B1(new_n871), .B2(new_n872), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(G301), .A3(new_n870), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n954), .A3(G168), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n944), .ZN(new_n957));
  INV_X1    g532(.A(new_n927), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n957), .B(new_n958), .C1(new_n937), .C2(new_n956), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n941), .A2(new_n943), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n952), .B2(new_n955), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n952), .A2(new_n955), .A3(new_n936), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n927), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n959), .A2(new_n963), .A3(new_n915), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n959), .A2(new_n963), .A3(new_n966), .A4(new_n915), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n968), .B(new_n969), .ZN(G397));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n490), .B1(new_n464), .B2(G126), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n493), .B1(new_n972), .B2(new_n460), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n498), .A2(new_n499), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT50), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n775), .A2(G40), .A3(new_n462), .A4(new_n465), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n979), .B(new_n971), .C1(new_n973), .C2(new_n974), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n976), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G1348), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n500), .A2(G160), .A3(G40), .A4(new_n971), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT118), .B1(new_n984), .B2(G2067), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n975), .A2(new_n977), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n841), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n983), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n930), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n983), .A2(new_n627), .A3(new_n985), .A4(new_n988), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(KEYINPUT60), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n981), .A2(new_n853), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n975), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g570(.A(KEYINPUT45), .B(new_n971), .C1(new_n973), .C2(new_n974), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT56), .B(G2072), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n995), .A2(new_n978), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n993), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n585), .A2(KEYINPUT116), .A3(new_n589), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT57), .ZN(new_n1001));
  NAND3_X1  g576(.A1(G299), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n583), .A2(new_n584), .B1(new_n588), .B2(G651), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1003), .B(new_n591), .C1(KEYINPUT116), .C2(KEYINPUT57), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n999), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1007), .A2(new_n993), .A3(new_n998), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(KEYINPUT61), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n992), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT117), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1007), .A2(new_n993), .A3(KEYINPUT117), .A4(new_n998), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT61), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1010), .A2(new_n1014), .ZN(new_n1015));
  OR2_X1    g590(.A1(new_n991), .A2(KEYINPUT60), .ZN(new_n1016));
  AND2_X1   g591(.A1(new_n995), .A2(new_n996), .ZN(new_n1017));
  INV_X1    g592(.A(G1996), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(KEYINPUT119), .A3(new_n1018), .A4(new_n978), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT58), .B(G1341), .Z(new_n1020));
  NAND2_X1  g595(.A1(new_n984), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n995), .A2(new_n978), .A3(new_n996), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(G1996), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(new_n1021), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT59), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n574), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n1025), .B2(new_n574), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT120), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1025), .A2(new_n574), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(KEYINPUT59), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1025), .A2(new_n1026), .A3(new_n574), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1015), .A2(new_n1016), .A3(new_n1029), .A4(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n989), .A2(new_n627), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1006), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1012), .B(new_n1013), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT125), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n602), .B2(G1976), .ZN(new_n1042));
  INV_X1    g617(.A(G1976), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G288), .A2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(G8), .B1(new_n975), .B2(new_n977), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(KEYINPUT110), .B(G8), .C1(new_n975), .C2(new_n977), .ZN(new_n1048));
  AOI211_X1 g623(.A(new_n1042), .B(new_n1044), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1044), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT52), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1049), .B1(new_n1053), .B2(KEYINPUT111), .ZN(new_n1054));
  INV_X1    g629(.A(G1981), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n607), .A2(new_n611), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n507), .A2(G61), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n521), .B1(new_n1057), .B2(new_n608), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n512), .B1(new_n604), .B2(new_n605), .ZN(new_n1059));
  OAI21_X1  g634(.A(G1981), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1056), .A2(new_n1060), .A3(KEYINPUT49), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT49), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT112), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI211_X1 g639(.A(KEYINPUT112), .B(KEYINPUT49), .C1(new_n1056), .C2(new_n1060), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1050), .B(new_n1061), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1042), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(KEYINPUT111), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1054), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G8), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT55), .B1(G166), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n1074));
  NAND3_X1  g649(.A1(G303), .A2(new_n1074), .A3(G8), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n981), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT108), .B(G2090), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1971), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1023), .A2(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1076), .B1(new_n1082), .B2(new_n1072), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1023), .A2(G2078), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(KEYINPUT123), .B2(KEYINPUT53), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1077), .A2(G1961), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1023), .B2(G2078), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(KEYINPUT124), .A2(KEYINPUT54), .ZN(new_n1090));
  MUX2_X1   g665(.A(new_n1090), .B(KEYINPUT54), .S(G301), .Z(new_n1091));
  OR2_X1    g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1081), .A2(KEYINPUT107), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT107), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1023), .A2(new_n1094), .A3(new_n1080), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n1079), .A3(new_n1095), .ZN(new_n1096));
  NOR3_X1   g671(.A1(G166), .A2(KEYINPUT55), .A3(new_n1072), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1074), .B1(G303), .B2(G8), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT109), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT109), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1073), .A2(new_n1075), .A3(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1096), .A2(G8), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1071), .A2(new_n1083), .A3(new_n1092), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1023), .A2(new_n824), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n976), .A2(new_n778), .A3(new_n978), .A4(new_n980), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(G8), .ZN(new_n1107));
  NAND3_X1  g682(.A1(G286), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1109), .B1(G168), .B2(new_n1072), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1107), .A2(new_n1111), .A3(KEYINPUT51), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1072), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1115), .A2(new_n1106), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n1115), .B2(new_n1106), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1112), .B(new_n1116), .C1(new_n1118), .C2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1040), .B1(new_n1103), .B2(new_n1122), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT111), .B1(new_n1067), .B2(new_n1041), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1052), .B2(new_n1042), .ZN(new_n1127));
  AND4_X1   g702(.A1(new_n1083), .A2(new_n1125), .A3(new_n1102), .A4(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1124), .A2(KEYINPUT125), .A3(new_n1128), .A4(new_n1092), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1039), .A2(new_n1123), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1120), .A2(KEYINPUT62), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1089), .A2(G171), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1115), .A2(new_n1106), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT122), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1115), .A2(new_n1106), .A3(new_n1117), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n1112), .A4(new_n1116), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1131), .A2(new_n1132), .A3(new_n1138), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1107), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1128), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT113), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1054), .B2(new_n1070), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1125), .A2(new_n1127), .A3(KEYINPUT113), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1102), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n602), .A2(new_n1043), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT114), .Z(new_n1148));
  AND2_X1   g723(.A1(new_n1066), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1056), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1050), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1146), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1096), .A2(G8), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT115), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT115), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1096), .A2(new_n1155), .A3(G8), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1154), .A2(new_n1076), .A3(new_n1156), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1107), .A2(G286), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1157), .A2(new_n1143), .A3(new_n1158), .A4(new_n1144), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1152), .B1(KEYINPUT63), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1130), .A2(new_n1141), .A3(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n838), .B(G2067), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n995), .A2(new_n977), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT105), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n1018), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(KEYINPUT104), .ZN(new_n1168));
  INV_X1    g743(.A(new_n792), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1163), .A2(G1996), .A3(new_n792), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1166), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT106), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n1172), .A2(KEYINPUT106), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n715), .A2(new_n724), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n715), .A2(new_n724), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1163), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(G290), .A2(G1986), .ZN(new_n1178));
  NOR2_X1   g753(.A1(G290), .A2(G1986), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1163), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  AND4_X1   g755(.A1(new_n1173), .A2(new_n1174), .A3(new_n1177), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1161), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1163), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1175), .B(KEYINPUT126), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1174), .A2(new_n1173), .A3(new_n1184), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n838), .A2(G2067), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1183), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1179), .A2(new_n1163), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT48), .ZN(new_n1189));
  AND4_X1   g764(.A1(new_n1173), .A2(new_n1174), .A3(new_n1177), .A4(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1163), .A2(new_n792), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1168), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1192), .A2(KEYINPUT46), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1192), .A2(KEYINPUT46), .ZN(new_n1194));
  OAI211_X1 g769(.A(new_n1191), .B(new_n1164), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT47), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1195), .B(new_n1196), .ZN(new_n1197));
  NOR3_X1   g772(.A1(new_n1187), .A2(new_n1190), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1182), .A2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g774(.A(G227), .ZN(new_n1201));
  NAND2_X1  g775(.A1(new_n1201), .A2(G319), .ZN(new_n1202));
  XNOR2_X1  g776(.A(new_n1202), .B(KEYINPUT127), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n1203), .B1(new_n965), .B2(new_n967), .ZN(new_n1204));
  NAND4_X1  g778(.A1(new_n1204), .A2(new_n669), .A3(new_n703), .A4(new_n916), .ZN(G225));
  INV_X1    g779(.A(G225), .ZN(G308));
endmodule


