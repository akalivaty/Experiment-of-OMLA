//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n634, new_n637, new_n639, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND3_X1  g030(.A1(new_n451), .A2(KEYINPUT67), .A3(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g033(.A(KEYINPUT67), .B1(new_n451), .B2(G2106), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT69), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT69), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  AND3_X1   g049(.A1(new_n472), .A2(new_n474), .A3(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n467), .B1(new_n470), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT71), .B1(new_n473), .B2(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT71), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(new_n471), .A3(G2104), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n477), .A2(new_n479), .A3(new_n474), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n480), .A2(G137), .A3(new_n466), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n462), .A2(G2104), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT72), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G101), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n476), .A2(new_n481), .A3(new_n484), .ZN(G160));
  NAND3_X1  g060(.A1(new_n477), .A2(new_n479), .A3(new_n474), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(new_n466), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n486), .A2(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  OAI221_X1 g065(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n466), .C2(G112), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT73), .Z(G162));
  AND2_X1   g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n477), .A2(new_n479), .A3(new_n474), .A4(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT74), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n462), .A2(G114), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n502), .A2(new_n497), .A3(KEYINPUT74), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n495), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n463), .A2(new_n465), .A3(G138), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n486), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT3), .B(G2104), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n466), .A2(new_n507), .A3(new_n508), .A4(G138), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n504), .B1(new_n506), .B2(new_n509), .ZN(G164));
  XNOR2_X1  g085(.A(KEYINPUT5), .B(G543), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT75), .B(G651), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT75), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT75), .A2(G651), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT6), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g096(.A(new_n516), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G50), .ZN(new_n523));
  AND2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n526), .B1(new_n519), .B2(new_n521), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G88), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n515), .A2(new_n523), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n526), .A2(KEYINPUT76), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n511), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n531), .A2(new_n533), .A3(G63), .A4(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT77), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XOR2_X1   g111(.A(new_n536), .B(KEYINPUT7), .Z(new_n537));
  AOI21_X1  g112(.A(new_n537), .B1(new_n522), .B2(G51), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n527), .A2(G89), .ZN(new_n539));
  AND2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g115(.A1(new_n535), .A2(new_n540), .ZN(G168));
  AOI22_X1  g116(.A1(G52), .A2(new_n522), .B1(new_n527), .B2(G90), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n531), .A2(new_n533), .A3(G64), .ZN(new_n544));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n514), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n543), .A2(new_n546), .ZN(G171));
  AOI22_X1  g122(.A1(G43), .A2(new_n522), .B1(new_n527), .B2(G81), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n531), .A2(new_n533), .A3(G56), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  AND2_X1   g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n548), .B1(new_n551), .B2(new_n514), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(KEYINPUT78), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n522), .A2(G43), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n519), .A2(new_n521), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(new_n511), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n554), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n514), .B1(new_n549), .B2(new_n550), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT78), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n553), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  AND2_X1   g143(.A1(KEYINPUT79), .A2(G53), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT6), .ZN(new_n570));
  OR2_X1    g145(.A1(KEYINPUT75), .A2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(KEYINPUT75), .A2(G651), .ZN(new_n572));
  AOI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g148(.A(G543), .B(new_n569), .C1(new_n573), .C2(new_n520), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n527), .A2(G91), .ZN(new_n577));
  OAI21_X1  g152(.A(G65), .B1(new_n524), .B2(new_n525), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT80), .B1(new_n580), .B2(G651), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  INV_X1    g157(.A(G651), .ZN(new_n583));
  AOI211_X1 g158(.A(new_n582), .B(new_n583), .C1(new_n578), .C2(new_n579), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n577), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  OR2_X1    g160(.A1(new_n576), .A2(new_n585), .ZN(G299));
  NAND2_X1  g161(.A1(new_n544), .A2(new_n545), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(new_n513), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(new_n542), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n589), .A2(KEYINPUT81), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n588), .B2(new_n542), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n590), .A2(new_n592), .ZN(G301));
  NAND2_X1  g168(.A1(new_n535), .A2(new_n540), .ZN(G286));
  AND2_X1   g169(.A1(new_n531), .A2(new_n533), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n595), .B2(G74), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n527), .A2(G87), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n522), .A2(G49), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G288));
  INV_X1    g174(.A(KEYINPUT83), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n520), .B1(new_n513), .B2(KEYINPUT6), .ZN(new_n601));
  NAND2_X1  g176(.A1(G48), .A2(G543), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n556), .A2(KEYINPUT83), .A3(G48), .A4(G543), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G73), .ZN(new_n606));
  OAI21_X1  g181(.A(KEYINPUT82), .B1(new_n606), .B2(new_n516), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n608), .A2(G73), .A3(G543), .ZN(new_n609));
  INV_X1    g184(.A(G61), .ZN(new_n610));
  OAI211_X1 g185(.A(new_n607), .B(new_n609), .C1(new_n526), .C2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(G86), .A2(new_n527), .B1(new_n611), .B2(new_n513), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT84), .ZN(G305));
  AOI22_X1  g189(.A1(new_n595), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n615), .A2(new_n514), .ZN(new_n616));
  AOI22_X1  g191(.A1(G47), .A2(new_n522), .B1(new_n527), .B2(G85), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(G290));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NOR2_X1   g194(.A1(G301), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n527), .A2(G92), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(G79), .ZN(new_n624));
  OR3_X1    g199(.A1(new_n624), .A2(new_n516), .A3(KEYINPUT85), .ZN(new_n625));
  OAI21_X1  g200(.A(KEYINPUT85), .B1(new_n624), .B2(new_n516), .ZN(new_n626));
  INV_X1    g201(.A(G66), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n526), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n628), .A2(G651), .B1(new_n522), .B2(G54), .ZN(new_n629));
  AND2_X1   g204(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT86), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n620), .B1(new_n631), .B2(new_n619), .ZN(G284));
  AOI21_X1  g207(.A(new_n620), .B1(new_n631), .B2(new_n619), .ZN(G321));
  NAND2_X1  g208(.A1(G299), .A2(new_n619), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n619), .B2(G168), .ZN(G297));
  OAI21_X1  g210(.A(new_n634), .B1(new_n619), .B2(G168), .ZN(G280));
  INV_X1    g211(.A(G559), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n631), .B1(new_n637), .B2(G860), .ZN(G148));
  NAND2_X1  g213(.A1(new_n631), .A2(new_n637), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT87), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G868), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(G868), .B2(new_n563), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g218(.A1(new_n483), .A2(new_n507), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT88), .B(KEYINPUT12), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT13), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT89), .B(G2100), .Z(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT90), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n487), .A2(G123), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n489), .A2(G135), .ZN(new_n652));
  OAI221_X1 g227(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n466), .C2(G111), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OAI22_X1  g229(.A1(new_n647), .A2(new_n648), .B1(G2096), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(G2096), .B2(new_n654), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n650), .A2(new_n656), .ZN(G156));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n661), .A2(KEYINPUT14), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT91), .B(KEYINPUT16), .Z(new_n669));
  XNOR2_X1  g244(.A(G2451), .B(G2454), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(G14), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n672), .B2(new_n668), .ZN(G401));
  XNOR2_X1  g249(.A(G2072), .B(G2078), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT17), .ZN(new_n676));
  XNOR2_X1  g251(.A(G2067), .B(G2678), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT93), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n682), .B(new_n679), .C1(new_n675), .C2(new_n677), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n678), .A2(new_n675), .A3(new_n677), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n681), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G2096), .B(G2100), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XOR2_X1   g264(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n690));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1956), .B(G2474), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1961), .B(G1966), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n693), .A2(new_n694), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n692), .A2(new_n695), .A3(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n692), .A2(new_n700), .ZN(new_n702));
  NOR4_X1   g277(.A1(new_n698), .A2(new_n699), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT96), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1981), .B(G1986), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(G229));
  MUX2_X1   g287(.A(G6), .B(G305), .S(G16), .Z(new_n713));
  XOR2_X1   g288(.A(KEYINPUT32), .B(G1981), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT99), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT98), .B(G16), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(G22), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G166), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G1971), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G23), .B(G288), .S(G16), .Z(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT33), .B(G1976), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n716), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT34), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n487), .A2(G119), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n489), .A2(G131), .ZN(new_n730));
  OAI221_X1 g305(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n466), .C2(G107), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT97), .B(G29), .Z(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G25), .B2(new_n735), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT35), .B(G1991), .Z(new_n738));
  AND2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n717), .A2(G24), .ZN(new_n740));
  INV_X1    g315(.A(G290), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(new_n717), .ZN(new_n742));
  OAI22_X1  g317(.A1(new_n742), .A2(G1986), .B1(new_n738), .B2(new_n737), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n739), .B(new_n743), .C1(G1986), .C2(new_n742), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n728), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT36), .ZN(new_n746));
  INV_X1    g321(.A(G16), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G4), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n631), .B2(new_n747), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(G1348), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n734), .A2(G26), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT28), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n487), .A2(G128), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n489), .A2(G140), .ZN(new_n754));
  OAI221_X1 g329(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n466), .C2(G116), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n752), .B1(new_n756), .B2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G2067), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n718), .A2(G19), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n563), .B2(new_n718), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G1341), .Z(new_n761));
  NAND3_X1  g336(.A1(new_n750), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT100), .ZN(new_n763));
  INV_X1    g338(.A(G21), .ZN(new_n764));
  AOI21_X1  g339(.A(KEYINPUT102), .B1(new_n747), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(G168), .A2(G16), .ZN(new_n766));
  MUX2_X1   g341(.A(KEYINPUT102), .B(new_n765), .S(new_n766), .Z(new_n767));
  NOR2_X1   g342(.A1(new_n767), .A2(G1966), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT103), .ZN(new_n769));
  NAND2_X1  g344(.A1(G162), .A2(new_n735), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G35), .B2(new_n735), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT29), .B(G2090), .Z(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n717), .A2(G20), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT23), .Z(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G299), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1956), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n773), .A2(new_n774), .A3(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n747), .A2(G5), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G171), .B2(new_n747), .ZN(new_n782));
  INV_X1    g357(.A(G1961), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(G160), .A2(G29), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT24), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(G34), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(G34), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n734), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G2084), .ZN(new_n792));
  INV_X1    g367(.A(G33), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n793), .A2(G29), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT25), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n489), .A2(G139), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n507), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n797), .B(new_n798), .C1(new_n466), .C2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n794), .B1(new_n800), .B2(G29), .ZN(new_n801));
  INV_X1    g376(.A(G2072), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(new_n654), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(new_n735), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT31), .B(G11), .Z(new_n806));
  INV_X1    g381(.A(G28), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(KEYINPUT30), .ZN(new_n808));
  AOI21_X1  g383(.A(G29), .B1(new_n807), .B2(KEYINPUT30), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n792), .A2(new_n803), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n735), .A2(G27), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G164), .B2(new_n735), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G2078), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n785), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT26), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n483), .A2(G105), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n487), .A2(G129), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n489), .A2(G141), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  MUX2_X1   g398(.A(G32), .B(new_n823), .S(G29), .Z(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT27), .B(G1996), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n824), .B(new_n825), .Z(new_n826));
  NOR2_X1   g401(.A1(new_n801), .A2(new_n802), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT101), .ZN(new_n828));
  AOI211_X1 g403(.A(new_n826), .B(new_n828), .C1(G1966), .C2(new_n767), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n769), .A2(new_n780), .A3(new_n815), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n763), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n746), .A2(new_n831), .ZN(G311));
  NAND2_X1  g407(.A1(new_n746), .A2(new_n831), .ZN(G150));
  INV_X1    g408(.A(G860), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n595), .A2(G67), .ZN(new_n835));
  NAND2_X1  g410(.A1(G80), .A2(G543), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n514), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n522), .A2(G55), .ZN(new_n838));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(new_n557), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n552), .A2(KEYINPUT78), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n560), .A2(new_n561), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n552), .A2(new_n837), .A3(new_n840), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n631), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n847), .B(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n834), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(KEYINPUT39), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n849), .A2(KEYINPUT104), .A3(KEYINPUT39), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n856));
  INV_X1    g431(.A(new_n841), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(G860), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT37), .ZN(new_n859));
  OR3_X1    g434(.A1(new_n855), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n856), .B1(new_n855), .B2(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(G145));
  XNOR2_X1  g437(.A(G162), .B(new_n804), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT106), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(G160), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n732), .B(KEYINPUT107), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n487), .A2(G130), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n489), .A2(G142), .ZN(new_n868));
  OAI221_X1 g443(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n466), .C2(G118), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n866), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n800), .B(new_n823), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n506), .A2(new_n509), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n498), .A2(new_n496), .A3(new_n500), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT74), .B1(new_n502), .B2(new_n497), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n480), .A2(new_n494), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n756), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n646), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n873), .B(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(G37), .B1(new_n865), .B2(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n865), .B2(new_n881), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g459(.A(G305), .B(G290), .ZN(new_n885));
  XNOR2_X1  g460(.A(G288), .B(G303), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT42), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT108), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n887), .A2(KEYINPUT42), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT109), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n890), .A2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n623), .A2(new_n629), .ZN(new_n895));
  XNOR2_X1  g470(.A(G299), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n639), .B(KEYINPUT87), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n846), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n897), .A2(new_n846), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n846), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n640), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n630), .B(G299), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(KEYINPUT41), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n896), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n903), .B(new_n898), .C1(new_n905), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n894), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n890), .B(new_n891), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n911), .A2(new_n889), .B1(new_n908), .B2(new_n901), .ZN(new_n912));
  OAI21_X1  g487(.A(G868), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n857), .A2(new_n619), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(G295));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n914), .ZN(G331));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n917));
  XOR2_X1   g492(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n857), .B1(new_n562), .B2(new_n553), .ZN(new_n920));
  INV_X1    g495(.A(new_n845), .ZN(new_n921));
  NAND2_X1  g496(.A1(G171), .A2(new_n591), .ZN(new_n922));
  INV_X1    g497(.A(new_n592), .ZN(new_n923));
  AOI21_X1  g498(.A(G286), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(G286), .A2(new_n589), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n920), .B(new_n921), .C1(new_n924), .C2(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(G168), .B1(new_n590), .B2(new_n592), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n928), .B(new_n925), .C1(new_n844), .C2(new_n845), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n931), .A3(new_n904), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n904), .A2(KEYINPUT41), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n896), .A2(new_n906), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n933), .A2(new_n934), .A3(new_n927), .A4(new_n929), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n896), .B1(new_n927), .B2(new_n929), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n937), .A2(new_n931), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n919), .B1(new_n939), .B2(new_n887), .ZN(new_n940));
  INV_X1    g515(.A(new_n887), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n936), .B2(new_n938), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n943));
  INV_X1    g518(.A(G37), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n942), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n940), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n935), .ZN(new_n948));
  OR2_X1    g523(.A1(new_n948), .A2(new_n937), .ZN(new_n949));
  AOI21_X1  g524(.A(G37), .B1(new_n949), .B2(new_n941), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n939), .A2(new_n887), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n917), .B1(new_n947), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n951), .B1(new_n945), .B2(new_n946), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n955), .A2(new_n919), .B1(new_n950), .B2(new_n940), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n956), .B2(new_n917), .ZN(G397));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(G164), .B2(G1384), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n476), .A2(new_n481), .A3(new_n484), .A4(G40), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n959), .A2(G1996), .A3(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT46), .Z(new_n962));
  NOR2_X1   g537(.A1(new_n959), .A2(new_n960), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n756), .B(G2067), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n823), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT47), .Z(new_n967));
  XNOR2_X1  g542(.A(new_n823), .B(G1996), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(new_n964), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n732), .B(new_n738), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n963), .ZN(new_n972));
  INV_X1    g547(.A(G1986), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n741), .A2(new_n973), .A3(new_n963), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n974), .B(KEYINPUT127), .Z(new_n975));
  OAI21_X1  g550(.A(new_n972), .B1(new_n975), .B2(KEYINPUT48), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(KEYINPUT48), .B2(new_n975), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n969), .A2(new_n738), .A3(new_n733), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(G2067), .B2(new_n756), .ZN(new_n979));
  AOI211_X1 g554(.A(new_n967), .B(new_n977), .C1(new_n963), .C2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n981));
  INV_X1    g556(.A(G8), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n983));
  NOR3_X1   g558(.A1(G166), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n985));
  AOI22_X1  g560(.A1(G303), .A2(G8), .B1(new_n985), .B2(KEYINPUT55), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  AND4_X1   g562(.A1(G40), .A2(new_n476), .A3(new_n481), .A4(new_n484), .ZN(new_n988));
  AOI21_X1  g563(.A(G1384), .B1(new_n874), .B2(new_n877), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NOR3_X1   g566(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G2090), .ZN(new_n994));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n878), .A2(KEYINPUT45), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n959), .A2(new_n988), .A3(new_n996), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n993), .A2(new_n994), .B1(new_n997), .B2(new_n721), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n981), .B(new_n987), .C1(new_n998), .C2(new_n982), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n988), .B1(new_n989), .B2(KEYINPUT45), .ZN(new_n1000));
  AOI211_X1 g575(.A(new_n958), .B(G1384), .C1(new_n874), .C2(new_n877), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n721), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n989), .A2(new_n990), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n994), .A4(new_n988), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n982), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n987), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT114), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n1010));
  INV_X1    g585(.A(G1981), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n605), .A2(new_n612), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1011), .B1(new_n605), .B2(new_n612), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n613), .A2(G1981), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1016), .A2(KEYINPUT49), .A3(new_n1012), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n982), .B1(new_n988), .B2(new_n989), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1021), .B(new_n1018), .C1(new_n1020), .C2(G288), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n988), .A2(new_n989), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(G8), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G288), .A2(new_n1020), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT52), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1019), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n999), .A2(new_n1008), .A3(new_n1009), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT125), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1019), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1032), .A2(KEYINPUT125), .A3(new_n1008), .A4(new_n999), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g609(.A1(G286), .A2(G8), .B1(KEYINPUT122), .B2(KEYINPUT51), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n878), .A2(new_n995), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n960), .B1(new_n1037), .B2(KEYINPUT50), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n1004), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1036), .B1(new_n1039), .B2(G2084), .ZN(new_n1040));
  INV_X1    g615(.A(G2084), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n993), .A2(KEYINPUT116), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT115), .B1(new_n1043), .B2(G1966), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n1045));
  INV_X1    g620(.A(G1966), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n997), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1040), .A2(new_n1042), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1035), .B1(new_n1048), .B2(new_n982), .ZN(new_n1049));
  NOR2_X1   g624(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  OAI221_X1 g626(.A(new_n1035), .B1(KEYINPUT122), .B2(KEYINPUT51), .C1(new_n1048), .C2(new_n982), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G286), .A2(G8), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT117), .B1(new_n576), .B2(new_n585), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(KEYINPUT117), .B(new_n1058), .C1(new_n576), .C2(new_n585), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(G1956), .B1(new_n1038), .B2(new_n1004), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT56), .B(G2072), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1000), .A2(new_n1001), .A3(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1062), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1348), .B1(new_n1038), .B2(new_n1004), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1023), .A2(G2067), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1067), .B1(new_n1070), .B2(new_n895), .ZN(new_n1071));
  INV_X1    g646(.A(G1956), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n991), .B2(new_n992), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n959), .A2(new_n988), .A3(new_n996), .A4(new_n1064), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1073), .A2(new_n1061), .A3(new_n1060), .A4(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1071), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1067), .A2(KEYINPUT121), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1062), .B(new_n1078), .C1(new_n1063), .C2(new_n1066), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT61), .B1(new_n1080), .B2(new_n1075), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT119), .B(G1996), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n959), .A2(new_n988), .A3(new_n996), .A4(new_n1083), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT58), .B(G1341), .Z(new_n1085));
  NAND2_X1  g660(.A1(new_n1023), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n563), .ZN(new_n1088));
  NAND2_X1  g663(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n563), .A3(new_n1089), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT60), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1023), .A2(G2067), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1096), .B(KEYINPUT60), .C1(new_n993), .C2(G1348), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n630), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n895), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1067), .A2(KEYINPUT61), .A3(new_n1075), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1093), .A2(new_n1098), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1076), .B1(new_n1081), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n997), .B2(G2078), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(G2078), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n959), .A2(new_n988), .A3(new_n996), .A4(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n783), .B1(new_n991), .B2(new_n992), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1104), .A2(G301), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT124), .ZN(new_n1109));
  AOI21_X1  g684(.A(G1961), .B1(new_n1038), .B2(new_n1004), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1105), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1000), .A2(new_n1001), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1113), .A2(new_n1114), .A3(G301), .A4(new_n1104), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1104), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1107), .A2(KEYINPUT123), .A3(new_n1106), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1116), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1109), .B(new_n1115), .C1(new_n1120), .C2(G301), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(G301), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1113), .A2(new_n1104), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1122), .B1(new_n1124), .B2(G171), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1121), .A2(new_n1122), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1034), .A2(new_n1056), .A3(new_n1102), .A4(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(G288), .A2(G1976), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1013), .B1(new_n1019), .B2(new_n1128), .ZN(new_n1129));
  OAI22_X1  g704(.A1(new_n1009), .A2(new_n1031), .B1(new_n1129), .B2(new_n1024), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1048), .A2(new_n982), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(G168), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1133), .B2(new_n1028), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(new_n1131), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1132), .A2(new_n1032), .A3(new_n1136), .A4(G168), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1130), .B1(new_n1134), .B2(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1127), .A2(KEYINPUT126), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT126), .B1(new_n1127), .B2(new_n1138), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1056), .A2(KEYINPUT62), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1054), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(new_n1052), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1120), .A2(G301), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1030), .A2(new_n1033), .A3(new_n1145), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1141), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1139), .A2(new_n1140), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n971), .ZN(new_n1149));
  XNOR2_X1  g724(.A(G290), .B(new_n973), .ZN(new_n1150));
  AOI211_X1 g725(.A(new_n959), .B(new_n960), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n980), .B1(new_n1148), .B2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g727(.A(new_n460), .ZN(new_n1154));
  NOR4_X1   g728(.A1(G229), .A2(new_n1154), .A3(G401), .A4(G227), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n883), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g730(.A1(new_n956), .A2(new_n1156), .ZN(G308));
  OR2_X1    g731(.A1(new_n956), .A2(new_n1156), .ZN(G225));
endmodule


